module normal_multiplier (A,
    B,
    P);
 input [31:0] A;
 input [31:0] B;
 output [63:0] P;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;

 sky130_fd_sc_hd__inv_2 _11277_ (.A(net33),
    .Y(_01737_));
 sky130_fd_sc_hd__inv_12 _11278_ (.A(net28),
    .Y(_01748_));
 sky130_fd_sc_hd__clkinv_4 _11279_ (.A(net44),
    .Y(_01759_));
 sky130_fd_sc_hd__clkinv_16 _11280_ (.A(net27),
    .Y(_01769_));
 sky130_fd_sc_hd__clkinv_16 _11281_ (.A(net55),
    .Y(_01780_));
 sky130_fd_sc_hd__inv_12 _11282_ (.A(net26),
    .Y(_01791_));
 sky130_fd_sc_hd__inv_12 _11283_ (.A(net23),
    .Y(_01802_));
 sky130_fd_sc_hd__clkinv_4 _11284_ (.A(net59),
    .Y(_01813_));
 sky130_fd_sc_hd__inv_12 _11285_ (.A(net12),
    .Y(_01824_));
 sky130_fd_sc_hd__clkinv_16 _11286_ (.A(net60),
    .Y(_01835_));
 sky130_fd_sc_hd__inv_12 _11287_ (.A(net1),
    .Y(_01846_));
 sky130_fd_sc_hd__inv_12 _11288_ (.A(net29),
    .Y(_01857_));
 sky130_fd_sc_hd__clkinv_16 _11289_ (.A(net30),
    .Y(_01868_));
 sky130_fd_sc_hd__clkinv_16 _11290_ (.A(net31),
    .Y(_01879_));
 sky130_fd_sc_hd__clkinv_16 _11291_ (.A(net63),
    .Y(_01890_));
 sky130_fd_sc_hd__inv_12 _11292_ (.A(net2),
    .Y(_01901_));
 sky130_fd_sc_hd__inv_12 _11293_ (.A(net32),
    .Y(_01912_));
 sky130_fd_sc_hd__inv_12 _11294_ (.A(net3),
    .Y(_01923_));
 sky130_fd_sc_hd__clkinv_16 _11295_ (.A(net35),
    .Y(_01934_));
 sky130_fd_sc_hd__inv_16 _11296_ (.A(net4),
    .Y(_01945_));
 sky130_fd_sc_hd__inv_8 _11297_ (.A(net5),
    .Y(_01956_));
 sky130_fd_sc_hd__inv_12 _11298_ (.A(net6),
    .Y(_01966_));
 sky130_fd_sc_hd__inv_16 _11299_ (.A(net7),
    .Y(_01977_));
 sky130_fd_sc_hd__inv_12 _11300_ (.A(net8),
    .Y(_01988_));
 sky130_fd_sc_hd__inv_12 _11301_ (.A(net9),
    .Y(_01999_));
 sky130_fd_sc_hd__clkinv_16 _11302_ (.A(net41),
    .Y(_02010_));
 sky130_fd_sc_hd__inv_12 _11303_ (.A(net10),
    .Y(_02021_));
 sky130_fd_sc_hd__inv_12 _11304_ (.A(net11),
    .Y(_02032_));
 sky130_fd_sc_hd__inv_8 _11305_ (.A(net13),
    .Y(_02043_));
 sky130_fd_sc_hd__clkinv_16 _11306_ (.A(net45),
    .Y(_02054_));
 sky130_fd_sc_hd__clkinv_16 _11307_ (.A(net14),
    .Y(_02065_));
 sky130_fd_sc_hd__inv_12 _11308_ (.A(net15),
    .Y(_02076_));
 sky130_fd_sc_hd__clkinv_8 _11309_ (.A(net47),
    .Y(_02087_));
 sky130_fd_sc_hd__inv_8 _11310_ (.A(net16),
    .Y(_02098_));
 sky130_fd_sc_hd__inv_16 _11311_ (.A(net48),
    .Y(_02109_));
 sky130_fd_sc_hd__inv_12 _11312_ (.A(net49),
    .Y(_02120_));
 sky130_fd_sc_hd__clkinv_16 _11313_ (.A(net18),
    .Y(_02131_));
 sky130_fd_sc_hd__inv_12 _11314_ (.A(net19),
    .Y(_02142_));
 sky130_fd_sc_hd__clkinv_16 _11315_ (.A(net51),
    .Y(_02152_));
 sky130_fd_sc_hd__clkinv_16 _11316_ (.A(net20),
    .Y(_02163_));
 sky130_fd_sc_hd__inv_4 _11317_ (.A(net52),
    .Y(_02174_));
 sky130_fd_sc_hd__clkinv_16 _11318_ (.A(net21),
    .Y(_02185_));
 sky130_fd_sc_hd__inv_8 _11319_ (.A(net22),
    .Y(_02196_));
 sky130_fd_sc_hd__inv_16 _11320_ (.A(net54),
    .Y(_02207_));
 sky130_fd_sc_hd__inv_16 _11321_ (.A(net24),
    .Y(_02218_));
 sky130_fd_sc_hd__inv_16 _11322_ (.A(net56),
    .Y(_02229_));
 sky130_fd_sc_hd__inv_16 _11323_ (.A(net57),
    .Y(_02240_));
 sky130_fd_sc_hd__inv_12 _11324_ (.A(net25),
    .Y(_02251_));
 sky130_fd_sc_hd__nor2_1 _11325_ (.A(_01737_),
    .B(_01846_),
    .Y(net65));
 sky130_fd_sc_hd__or4_4 _11326_ (.A(_01737_),
    .B(_01759_),
    .C(_01824_),
    .D(_01846_),
    .X(_02272_));
 sky130_fd_sc_hd__nand4_2 _11327_ (.A(net33),
    .B(net44),
    .C(net23),
    .D(net12),
    .Y(_02283_));
 sky130_fd_sc_hd__a22o_1 _11328_ (.A1(net33),
    .A2(net23),
    .B1(net12),
    .B2(net44),
    .X(_02294_));
 sky130_fd_sc_hd__nand4_1 _11329_ (.A(_02294_),
    .B(net1),
    .C(net55),
    .D(_02283_),
    .Y(_02305_));
 sky130_fd_sc_hd__a22o_1 _11330_ (.A1(net55),
    .A2(net1),
    .B1(_02283_),
    .B2(_02294_),
    .X(_02316_));
 sky130_fd_sc_hd__nand2_1 _11331_ (.A(_02305_),
    .B(_02316_),
    .Y(_02327_));
 sky130_fd_sc_hd__nand2_1 _11332_ (.A(net58),
    .B(net1),
    .Y(_02338_));
 sky130_fd_sc_hd__nand2_1 _11333_ (.A(net44),
    .B(net26),
    .Y(_02349_));
 sky130_fd_sc_hd__and4_1 _11334_ (.A(net33),
    .B(net44),
    .C(net26),
    .D(net23),
    .X(_02360_));
 sky130_fd_sc_hd__nand4_1 _11335_ (.A(net33),
    .B(net44),
    .C(net26),
    .D(net23),
    .Y(_02370_));
 sky130_fd_sc_hd__a22o_1 _11336_ (.A1(net33),
    .A2(net26),
    .B1(net23),
    .B2(net44),
    .X(_02381_));
 sky130_fd_sc_hd__o2bb2a_1 _11337_ (.A1_N(_02370_),
    .A2_N(_02381_),
    .B1(_01780_),
    .B2(_01824_),
    .X(_02392_));
 sky130_fd_sc_hd__and4_1 _11338_ (.A(_02381_),
    .B(net12),
    .C(net55),
    .D(_02370_),
    .X(_02403_));
 sky130_fd_sc_hd__a211oi_1 _11339_ (.A1(_02283_),
    .A2(_02305_),
    .B1(_02392_),
    .C1(_02403_),
    .Y(_02414_));
 sky130_fd_sc_hd__o211a_1 _11340_ (.A1(_02392_),
    .A2(_02403_),
    .B1(_02283_),
    .C1(_02305_),
    .X(_02425_));
 sky130_fd_sc_hd__or3_1 _11341_ (.A(_02338_),
    .B(_02414_),
    .C(_02425_),
    .X(_02436_));
 sky130_fd_sc_hd__a2bb2o_1 _11342_ (.A1_N(_02414_),
    .A2_N(_02425_),
    .B1(net58),
    .B2(net1),
    .X(_02447_));
 sky130_fd_sc_hd__or4bb_2 _11343_ (.A(_02272_),
    .B(_02327_),
    .C_N(_02436_),
    .D_N(_02447_),
    .X(_02458_));
 sky130_fd_sc_hd__o21ba_1 _11344_ (.A1(_02338_),
    .A2(_02425_),
    .B1_N(_02414_),
    .X(_02469_));
 sky130_fd_sc_hd__a31o_1 _11345_ (.A1(_02381_),
    .A2(net12),
    .A3(net55),
    .B1(_02360_),
    .X(_02480_));
 sky130_fd_sc_hd__nand2_1 _11346_ (.A(net55),
    .B(net23),
    .Y(_02491_));
 sky130_fd_sc_hd__nand2_2 _11347_ (.A(net33),
    .B(net27),
    .Y(_02502_));
 sky130_fd_sc_hd__a22o_1 _11348_ (.A1(net33),
    .A2(net27),
    .B1(net26),
    .B2(net44),
    .X(_02513_));
 sky130_fd_sc_hd__and4_1 _11349_ (.A(net33),
    .B(net44),
    .C(net27),
    .D(net26),
    .X(_02524_));
 sky130_fd_sc_hd__nand4_1 _11350_ (.A(net33),
    .B(net44),
    .C(net27),
    .D(net26),
    .Y(_02535_));
 sky130_fd_sc_hd__a22o_1 _11351_ (.A1(net55),
    .A2(net23),
    .B1(_02513_),
    .B2(_02535_),
    .X(_02546_));
 sky130_fd_sc_hd__nand4_1 _11352_ (.A(_02513_),
    .B(_02535_),
    .C(net55),
    .D(net23),
    .Y(_02557_));
 sky130_fd_sc_hd__a21o_1 _11353_ (.A1(_02546_),
    .A2(_02557_),
    .B1(_02480_),
    .X(_02568_));
 sky130_fd_sc_hd__o211ai_2 _11354_ (.A1(_02360_),
    .A2(_02403_),
    .B1(_02546_),
    .C1(_02557_),
    .Y(_02578_));
 sky130_fd_sc_hd__nor2_1 _11355_ (.A(_01813_),
    .B(_01824_),
    .Y(_02589_));
 sky130_fd_sc_hd__and3_1 _11356_ (.A(net58),
    .B(net1),
    .C(_02589_),
    .X(_02600_));
 sky130_fd_sc_hd__o2bb2a_1 _11357_ (.A1_N(net58),
    .A2_N(net12),
    .B1(_01846_),
    .B2(_01813_),
    .X(_02611_));
 sky130_fd_sc_hd__a31o_1 _11358_ (.A1(net58),
    .A2(net1),
    .A3(_02589_),
    .B1(_02611_),
    .X(_02622_));
 sky130_fd_sc_hd__a21bo_1 _11359_ (.A1(_02568_),
    .A2(_02578_),
    .B1_N(_02622_),
    .X(_02633_));
 sky130_fd_sc_hd__nand3b_1 _11360_ (.A_N(_02622_),
    .B(_02578_),
    .C(_02568_),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2_1 _11361_ (.A(_02633_),
    .B(_02644_),
    .Y(_02655_));
 sky130_fd_sc_hd__nor2_1 _11362_ (.A(_02469_),
    .B(_02655_),
    .Y(_02666_));
 sky130_fd_sc_hd__and2_1 _11363_ (.A(_02655_),
    .B(_02469_),
    .X(_02677_));
 sky130_fd_sc_hd__or2_1 _11364_ (.A(_02666_),
    .B(_02677_),
    .X(_02688_));
 sky130_fd_sc_hd__nor2_1 _11365_ (.A(_02458_),
    .B(_02688_),
    .Y(_02699_));
 sky130_fd_sc_hd__a21boi_1 _11366_ (.A1(_02578_),
    .A2(_02622_),
    .B1_N(_02568_),
    .Y(_02710_));
 sky130_fd_sc_hd__and4_1 _11367_ (.A(net23),
    .B(net58),
    .C(net59),
    .D(net12),
    .X(_02721_));
 sky130_fd_sc_hd__nand4_1 _11368_ (.A(net23),
    .B(net58),
    .C(net59),
    .D(net12),
    .Y(_02732_));
 sky130_fd_sc_hd__a22o_1 _11369_ (.A1(net23),
    .A2(net58),
    .B1(net59),
    .B2(net12),
    .X(_02743_));
 sky130_fd_sc_hd__a22oi_1 _11370_ (.A1(net60),
    .A2(net1),
    .B1(_02732_),
    .B2(_02743_),
    .Y(_02754_));
 sky130_fd_sc_hd__and4_1 _11371_ (.A(_02743_),
    .B(net1),
    .C(net60),
    .D(_02732_),
    .X(_02765_));
 sky130_fd_sc_hd__nor2_1 _11372_ (.A(_02754_),
    .B(_02765_),
    .Y(_02776_));
 sky130_fd_sc_hd__o21ai_1 _11373_ (.A1(_02349_),
    .A2(_02502_),
    .B1(_02491_),
    .Y(_02787_));
 sky130_fd_sc_hd__a21oi_1 _11374_ (.A1(_02349_),
    .A2(_02502_),
    .B1(_02491_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_1 _11375_ (.A(net55),
    .B(net26),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _11376_ (.A(net28),
    .B(net44),
    .Y(_02819_));
 sky130_fd_sc_hd__nand4_2 _11377_ (.A(net33),
    .B(net28),
    .C(net44),
    .D(net27),
    .Y(_02830_));
 sky130_fd_sc_hd__a22oi_1 _11378_ (.A1(net33),
    .A2(net28),
    .B1(net44),
    .B2(net27),
    .Y(_02841_));
 sky130_fd_sc_hd__a22o_2 _11379_ (.A1(net33),
    .A2(net28),
    .B1(net44),
    .B2(net27),
    .X(_02852_));
 sky130_fd_sc_hd__a22oi_1 _11380_ (.A1(net55),
    .A2(net26),
    .B1(_02830_),
    .B2(_02852_),
    .Y(_02863_));
 sky130_fd_sc_hd__a22o_1 _11381_ (.A1(net55),
    .A2(net26),
    .B1(_02830_),
    .B2(_02852_),
    .X(_02874_));
 sky130_fd_sc_hd__and4_1 _11382_ (.A(_02852_),
    .B(net26),
    .C(net55),
    .D(_02830_),
    .X(_02885_));
 sky130_fd_sc_hd__o2111ai_2 _11383_ (.A1(_02502_),
    .A2(_02819_),
    .B1(net55),
    .C1(net26),
    .D1(_02852_),
    .Y(_02896_));
 sky130_fd_sc_hd__o211a_1 _11384_ (.A1(_02524_),
    .A2(_02798_),
    .B1(_02874_),
    .C1(_02896_),
    .X(_02907_));
 sky130_fd_sc_hd__o211ai_2 _11385_ (.A1(_02524_),
    .A2(_02798_),
    .B1(_02874_),
    .C1(_02896_),
    .Y(_02918_));
 sky130_fd_sc_hd__o2bb2ai_2 _11386_ (.A1_N(_02513_),
    .A2_N(_02787_),
    .B1(_02863_),
    .B2(_02885_),
    .Y(_02929_));
 sky130_fd_sc_hd__nand2_1 _11387_ (.A(_02929_),
    .B(_02776_),
    .Y(_02940_));
 sky130_fd_sc_hd__nand3_1 _11388_ (.A(_02929_),
    .B(_02776_),
    .C(_02918_),
    .Y(_02951_));
 sky130_fd_sc_hd__a2bb2o_1 _11389_ (.A1_N(_02754_),
    .A2_N(_02765_),
    .B1(_02918_),
    .B2(_02929_),
    .X(_02962_));
 sky130_fd_sc_hd__a21o_1 _11390_ (.A1(_02951_),
    .A2(_02962_),
    .B1(_02710_),
    .X(_02973_));
 sky130_fd_sc_hd__o211ai_2 _11391_ (.A1(_02907_),
    .A2(_02940_),
    .B1(_02962_),
    .C1(_02710_),
    .Y(_02984_));
 sky130_fd_sc_hd__a32o_1 _11392_ (.A1(net58),
    .A2(net1),
    .A3(_02589_),
    .B1(_02973_),
    .B2(_02984_),
    .X(_02995_));
 sky130_fd_sc_hd__nand3_2 _11393_ (.A(_02973_),
    .B(_02984_),
    .C(_02600_),
    .Y(_03006_));
 sky130_fd_sc_hd__o2bb2a_1 _11394_ (.A1_N(_02995_),
    .A2_N(_03006_),
    .B1(_02469_),
    .B2(_02655_),
    .X(_03017_));
 sky130_fd_sc_hd__a2bb2o_1 _11395_ (.A1_N(_02655_),
    .A2_N(_02469_),
    .B1(_03006_),
    .B2(_02995_),
    .X(_03028_));
 sky130_fd_sc_hd__nand3_1 _11396_ (.A(_02995_),
    .B(_03006_),
    .C(_02666_),
    .Y(_03039_));
 sky130_fd_sc_hd__a2bb2o_1 _11397_ (.A1_N(_02458_),
    .A2_N(_02688_),
    .B1(_03028_),
    .B2(_03039_),
    .X(_03050_));
 sky130_fd_sc_hd__nand2_1 _11398_ (.A(_02699_),
    .B(_03028_),
    .Y(_03060_));
 sky130_fd_sc_hd__o31a_1 _11399_ (.A1(_02458_),
    .A2(_02688_),
    .A3(_03017_),
    .B1(_03050_),
    .X(net120));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(_02984_),
    .B(_03006_),
    .Y(_03081_));
 sky130_fd_sc_hd__nand2_2 _11401_ (.A(net1),
    .B(net61),
    .Y(_03092_));
 sky130_fd_sc_hd__a31oi_4 _11402_ (.A1(_02743_),
    .A2(net1),
    .A3(net60),
    .B1(_02721_),
    .Y(_03103_));
 sky130_fd_sc_hd__or3b_2 _11403_ (.A(_01846_),
    .B(_03103_),
    .C_N(net61),
    .X(_03114_));
 sky130_fd_sc_hd__a211o_1 _11404_ (.A1(net1),
    .A2(net61),
    .B1(_02721_),
    .C1(_02765_),
    .X(_03125_));
 sky130_fd_sc_hd__xor2_1 _11405_ (.A(_03092_),
    .B(_03103_),
    .X(_03136_));
 sky130_fd_sc_hd__nand2_1 _11406_ (.A(_03114_),
    .B(_03125_),
    .Y(_03147_));
 sky130_fd_sc_hd__a21oi_2 _11407_ (.A1(_02929_),
    .A2(_02776_),
    .B1(_02907_),
    .Y(_03158_));
 sky130_fd_sc_hd__nand2_1 _11408_ (.A(net12),
    .B(net60),
    .Y(_03169_));
 sky130_fd_sc_hd__a22oi_1 _11409_ (.A1(net26),
    .A2(net58),
    .B1(net59),
    .B2(net23),
    .Y(_03180_));
 sky130_fd_sc_hd__a22o_1 _11410_ (.A1(net26),
    .A2(net58),
    .B1(net59),
    .B2(net23),
    .X(_03191_));
 sky130_fd_sc_hd__nand4_4 _11411_ (.A(net26),
    .B(net23),
    .C(net58),
    .D(net59),
    .Y(_03202_));
 sky130_fd_sc_hd__and3_2 _11412_ (.A(_03169_),
    .B(_03191_),
    .C(_03202_),
    .X(_03213_));
 sky130_fd_sc_hd__a21oi_2 _11413_ (.A1(_03191_),
    .A2(_03202_),
    .B1(_03169_),
    .Y(_03224_));
 sky130_fd_sc_hd__o2bb2ai_1 _11414_ (.A1_N(_03191_),
    .A2_N(_03202_),
    .B1(_01824_),
    .B2(_01835_),
    .Y(_03235_));
 sky130_fd_sc_hd__nand4_1 _11415_ (.A(_03191_),
    .B(_03202_),
    .C(net12),
    .D(net60),
    .Y(_03246_));
 sky130_fd_sc_hd__nand2_1 _11416_ (.A(_03235_),
    .B(_03246_),
    .Y(_03257_));
 sky130_fd_sc_hd__o21ai_2 _11417_ (.A1(_02502_),
    .A2(_02819_),
    .B1(_02808_),
    .Y(_03268_));
 sky130_fd_sc_hd__o21ai_2 _11418_ (.A1(_02808_),
    .A2(_02841_),
    .B1(_02830_),
    .Y(_03279_));
 sky130_fd_sc_hd__nand2_2 _11419_ (.A(net33),
    .B(net29),
    .Y(_03290_));
 sky130_fd_sc_hd__a22oi_4 _11420_ (.A1(net28),
    .A2(net44),
    .B1(net29),
    .B2(net33),
    .Y(_03301_));
 sky130_fd_sc_hd__a22o_1 _11421_ (.A1(net28),
    .A2(net44),
    .B1(net29),
    .B2(net33),
    .X(_03312_));
 sky130_fd_sc_hd__and4_2 _11422_ (.A(net33),
    .B(net28),
    .C(net44),
    .D(net29),
    .X(_03322_));
 sky130_fd_sc_hd__nand4_4 _11423_ (.A(net33),
    .B(net28),
    .C(net44),
    .D(net29),
    .Y(_03333_));
 sky130_fd_sc_hd__nand2_1 _11424_ (.A(net27),
    .B(net55),
    .Y(_03344_));
 sky130_fd_sc_hd__o22ai_4 _11425_ (.A1(_01769_),
    .A2(_01780_),
    .B1(_03301_),
    .B2(_03322_),
    .Y(_03355_));
 sky130_fd_sc_hd__nand4_4 _11426_ (.A(_03312_),
    .B(_03333_),
    .C(net27),
    .D(net55),
    .Y(_03366_));
 sky130_fd_sc_hd__and3_1 _11427_ (.A(_03355_),
    .B(_03366_),
    .C(_03279_),
    .X(_03377_));
 sky130_fd_sc_hd__nand4_1 _11428_ (.A(_02852_),
    .B(_03268_),
    .C(_03355_),
    .D(_03366_),
    .Y(_03388_));
 sky130_fd_sc_hd__a22oi_4 _11429_ (.A1(_02852_),
    .A2(_03268_),
    .B1(_03355_),
    .B2(_03366_),
    .Y(_03399_));
 sky130_fd_sc_hd__o22ai_4 _11430_ (.A1(_03213_),
    .A2(_03224_),
    .B1(_03377_),
    .B2(_03399_),
    .Y(_03410_));
 sky130_fd_sc_hd__nand3b_2 _11431_ (.A_N(_03399_),
    .B(_03257_),
    .C(_03388_),
    .Y(_03421_));
 sky130_fd_sc_hd__nor2_1 _11432_ (.A(_03257_),
    .B(_03399_),
    .Y(_03432_));
 sky130_fd_sc_hd__a21oi_2 _11433_ (.A1(_03410_),
    .A2(_03421_),
    .B1(_03158_),
    .Y(_03443_));
 sky130_fd_sc_hd__a22o_1 _11434_ (.A1(_02918_),
    .A2(_02940_),
    .B1(_03410_),
    .B2(_03421_),
    .X(_03454_));
 sky130_fd_sc_hd__nand4_1 _11435_ (.A(_02918_),
    .B(_02940_),
    .C(_03410_),
    .D(_03421_),
    .Y(_03465_));
 sky130_fd_sc_hd__a31oi_4 _11436_ (.A1(_03158_),
    .A2(_03410_),
    .A3(_03421_),
    .B1(_03147_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _11437_ (.A(_03476_),
    .B(_03454_),
    .Y(_03487_));
 sky130_fd_sc_hd__a21o_1 _11438_ (.A1(_03454_),
    .A2(_03465_),
    .B1(_03136_),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_1 _11439_ (.A1(_03487_),
    .A2(_03498_),
    .B1(_03081_),
    .X(_03509_));
 sky130_fd_sc_hd__nand3_2 _11440_ (.A(_03081_),
    .B(_03487_),
    .C(_03498_),
    .Y(_03520_));
 sky130_fd_sc_hd__inv_2 _11441_ (.A(_03520_),
    .Y(_03531_));
 sky130_fd_sc_hd__nand2_1 _11442_ (.A(_03509_),
    .B(_03520_),
    .Y(_03542_));
 sky130_fd_sc_hd__o31a_1 _11443_ (.A1(_02458_),
    .A2(_02688_),
    .A3(_03017_),
    .B1(_03039_),
    .X(_03553_));
 sky130_fd_sc_hd__a32o_1 _11444_ (.A1(_02666_),
    .A2(_02995_),
    .A3(_03006_),
    .B1(_02699_),
    .B2(_03028_),
    .X(_03564_));
 sky130_fd_sc_hd__a21o_1 _11445_ (.A1(_03509_),
    .A2(_03520_),
    .B1(_03564_),
    .X(_03575_));
 sky130_fd_sc_hd__nand4_2 _11446_ (.A(_02995_),
    .B(_03006_),
    .C(_03509_),
    .D(_02666_),
    .Y(_03586_));
 sky130_fd_sc_hd__o211a_1 _11447_ (.A1(_03060_),
    .A2(_03542_),
    .B1(_03575_),
    .C1(_03586_),
    .X(net125));
 sky130_fd_sc_hd__a21o_1 _11448_ (.A1(_03465_),
    .A2(_03136_),
    .B1(_03443_),
    .X(_03606_));
 sky130_fd_sc_hd__a311oi_4 _11449_ (.A1(_03355_),
    .A2(_03366_),
    .A3(_03279_),
    .B1(_03224_),
    .C1(_03213_),
    .Y(_03617_));
 sky130_fd_sc_hd__o21ai_1 _11450_ (.A1(_03257_),
    .A2(_03399_),
    .B1(_03388_),
    .Y(_03628_));
 sky130_fd_sc_hd__nand2_1 _11451_ (.A(net23),
    .B(net60),
    .Y(_03639_));
 sky130_fd_sc_hd__a22oi_4 _11452_ (.A1(net27),
    .A2(net58),
    .B1(net59),
    .B2(net26),
    .Y(_03650_));
 sky130_fd_sc_hd__a22o_1 _11453_ (.A1(net27),
    .A2(net58),
    .B1(net59),
    .B2(net26),
    .X(_03661_));
 sky130_fd_sc_hd__and4_1 _11454_ (.A(net27),
    .B(net26),
    .C(net58),
    .D(net59),
    .X(_03672_));
 sky130_fd_sc_hd__nand4_4 _11455_ (.A(net27),
    .B(net26),
    .C(net58),
    .D(net59),
    .Y(_03683_));
 sky130_fd_sc_hd__and4_1 _11456_ (.A(_03661_),
    .B(_03683_),
    .C(net23),
    .D(net60),
    .X(_03694_));
 sky130_fd_sc_hd__nand4_2 _11457_ (.A(_03661_),
    .B(_03683_),
    .C(net23),
    .D(net60),
    .Y(_03705_));
 sky130_fd_sc_hd__o22a_1 _11458_ (.A1(_01802_),
    .A2(_01835_),
    .B1(_03650_),
    .B2(_03672_),
    .X(_03716_));
 sky130_fd_sc_hd__o22ai_4 _11459_ (.A1(_01802_),
    .A2(_01835_),
    .B1(_03650_),
    .B2(_03672_),
    .Y(_03727_));
 sky130_fd_sc_hd__nand2_1 _11460_ (.A(_03705_),
    .B(_03727_),
    .Y(_03738_));
 sky130_fd_sc_hd__a21oi_2 _11461_ (.A1(_02819_),
    .A2(_03290_),
    .B1(_03344_),
    .Y(_03749_));
 sky130_fd_sc_hd__o21ai_2 _11462_ (.A1(_03344_),
    .A2(_03301_),
    .B1(_03333_),
    .Y(_03760_));
 sky130_fd_sc_hd__o31a_1 _11463_ (.A1(_01769_),
    .A2(_01780_),
    .A3(_03301_),
    .B1(_03333_),
    .X(_03771_));
 sky130_fd_sc_hd__nand2_1 _11464_ (.A(net28),
    .B(net55),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_2 _11465_ (.A(net44),
    .B(net30),
    .Y(_03793_));
 sky130_fd_sc_hd__nand4_4 _11466_ (.A(net33),
    .B(net44),
    .C(net29),
    .D(net30),
    .Y(_03804_));
 sky130_fd_sc_hd__a22oi_2 _11467_ (.A1(net44),
    .A2(net29),
    .B1(net30),
    .B2(net33),
    .Y(_03815_));
 sky130_fd_sc_hd__a22o_2 _11468_ (.A1(net44),
    .A2(net29),
    .B1(net30),
    .B2(net33),
    .X(_03826_));
 sky130_fd_sc_hd__o221ai_4 _11469_ (.A1(_01748_),
    .A2(_01780_),
    .B1(_03290_),
    .B2(_03793_),
    .C1(_03826_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21o_1 _11470_ (.A1(_03804_),
    .A2(_03826_),
    .B1(_03782_),
    .X(_03848_));
 sky130_fd_sc_hd__o2bb2ai_4 _11471_ (.A1_N(_03804_),
    .A2_N(_03826_),
    .B1(_01748_),
    .B2(_01780_),
    .Y(_03859_));
 sky130_fd_sc_hd__o2111ai_4 _11472_ (.A1(_03290_),
    .A2(_03793_),
    .B1(net28),
    .C1(net55),
    .D1(_03826_),
    .Y(_03870_));
 sky130_fd_sc_hd__a21oi_2 _11473_ (.A1(_03859_),
    .A2(_03870_),
    .B1(_03760_),
    .Y(_03880_));
 sky130_fd_sc_hd__nand3_1 _11474_ (.A(_03771_),
    .B(_03837_),
    .C(_03848_),
    .Y(_03891_));
 sky130_fd_sc_hd__o211a_1 _11475_ (.A1(_03322_),
    .A2(_03749_),
    .B1(_03859_),
    .C1(_03870_),
    .X(_03902_));
 sky130_fd_sc_hd__o211ai_4 _11476_ (.A1(_03322_),
    .A2(_03749_),
    .B1(_03859_),
    .C1(_03870_),
    .Y(_03913_));
 sky130_fd_sc_hd__and4_1 _11477_ (.A(_03705_),
    .B(_03727_),
    .C(_03891_),
    .D(_03913_),
    .X(_03924_));
 sky130_fd_sc_hd__nand3b_2 _11478_ (.A_N(_03738_),
    .B(_03891_),
    .C(_03913_),
    .Y(_03935_));
 sky130_fd_sc_hd__o22ai_4 _11479_ (.A1(_03694_),
    .A2(_03716_),
    .B1(_03880_),
    .B2(_03902_),
    .Y(_03946_));
 sky130_fd_sc_hd__a2bb2oi_4 _11480_ (.A1_N(_03399_),
    .A2_N(_03617_),
    .B1(_03935_),
    .B2(_03946_),
    .Y(_03957_));
 sky130_fd_sc_hd__a2bb2o_1 _11481_ (.A1_N(_03399_),
    .A2_N(_03617_),
    .B1(_03935_),
    .B2(_03946_),
    .X(_03968_));
 sky130_fd_sc_hd__o21ai_2 _11482_ (.A1(_03377_),
    .A2(_03432_),
    .B1(_03946_),
    .Y(_03979_));
 sky130_fd_sc_hd__o211a_1 _11483_ (.A1(_03377_),
    .A2(_03432_),
    .B1(_03935_),
    .C1(_03946_),
    .X(_03990_));
 sky130_fd_sc_hd__and2_1 _11484_ (.A(net12),
    .B(net62),
    .X(_04001_));
 sky130_fd_sc_hd__nand2_1 _11485_ (.A(net12),
    .B(net62),
    .Y(_04012_));
 sky130_fd_sc_hd__nand2_2 _11486_ (.A(net12),
    .B(net61),
    .Y(_04023_));
 sky130_fd_sc_hd__and3_1 _11487_ (.A(net1),
    .B(net61),
    .C(_04001_),
    .X(_04034_));
 sky130_fd_sc_hd__a22oi_1 _11488_ (.A1(net12),
    .A2(net61),
    .B1(net62),
    .B2(net1),
    .Y(_04045_));
 sky130_fd_sc_hd__a31o_1 _11489_ (.A1(net1),
    .A2(net61),
    .A3(_04001_),
    .B1(_04045_),
    .X(_04056_));
 sky130_fd_sc_hd__o31a_1 _11490_ (.A1(_01824_),
    .A2(_01835_),
    .A3(_03180_),
    .B1(_03202_),
    .X(_04067_));
 sky130_fd_sc_hd__a21oi_2 _11491_ (.A1(_03202_),
    .A2(_03246_),
    .B1(_04056_),
    .Y(_04078_));
 sky130_fd_sc_hd__o311a_1 _11492_ (.A1(_01824_),
    .A2(_01835_),
    .A3(_03180_),
    .B1(_03202_),
    .C1(_04056_),
    .X(_04089_));
 sky130_fd_sc_hd__nor2_1 _11493_ (.A(_04078_),
    .B(_04089_),
    .Y(_04100_));
 sky130_fd_sc_hd__or2_1 _11494_ (.A(_04078_),
    .B(_04089_),
    .X(_04111_));
 sky130_fd_sc_hd__o21ai_4 _11495_ (.A1(_03957_),
    .A2(_03990_),
    .B1(_04111_),
    .Y(_04122_));
 sky130_fd_sc_hd__o211ai_4 _11496_ (.A1(_03924_),
    .A2(_03979_),
    .B1(_04100_),
    .C1(_03968_),
    .Y(_04133_));
 sky130_fd_sc_hd__a21oi_2 _11497_ (.A1(_04122_),
    .A2(_04133_),
    .B1(_03606_),
    .Y(_04144_));
 sky130_fd_sc_hd__a21o_2 _11498_ (.A1(_04122_),
    .A2(_04133_),
    .B1(_03606_),
    .X(_04155_));
 sky130_fd_sc_hd__o211a_1 _11499_ (.A1(_03443_),
    .A2(_03476_),
    .B1(_04122_),
    .C1(_04133_),
    .X(_04166_));
 sky130_fd_sc_hd__o211ai_4 _11500_ (.A1(_03443_),
    .A2(_03476_),
    .B1(_04122_),
    .C1(_04133_),
    .Y(_04176_));
 sky130_fd_sc_hd__o22ai_4 _11501_ (.A1(_03092_),
    .A2(_03103_),
    .B1(_04144_),
    .B2(_04166_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand3b_4 _11502_ (.A_N(_03114_),
    .B(_04155_),
    .C(_04176_),
    .Y(_04198_));
 sky130_fd_sc_hd__nand2_1 _11503_ (.A(_04187_),
    .B(_04198_),
    .Y(_04209_));
 sky130_fd_sc_hd__a32o_1 _11504_ (.A1(_03081_),
    .A2(_03487_),
    .A3(_03498_),
    .B1(_04187_),
    .B2(_04198_),
    .X(_04220_));
 sky130_fd_sc_hd__nand3b_1 _11505_ (.A_N(_03520_),
    .B(_04187_),
    .C(_04198_),
    .Y(_04231_));
 sky130_fd_sc_hd__o211a_1 _11506_ (.A1(_03542_),
    .A2(_03553_),
    .B1(_04220_),
    .C1(_04231_),
    .X(_04242_));
 sky130_fd_sc_hd__a41o_1 _11507_ (.A1(_03509_),
    .A2(_03520_),
    .A3(_03564_),
    .A4(_04209_),
    .B1(_04242_),
    .X(net126));
 sky130_fd_sc_hd__nor3_1 _11508_ (.A(_03060_),
    .B(_03542_),
    .C(_04209_),
    .Y(_04263_));
 sky130_fd_sc_hd__o21ai_4 _11509_ (.A1(_03639_),
    .A2(_03650_),
    .B1(_03683_),
    .Y(_04274_));
 sky130_fd_sc_hd__nand2_2 _11510_ (.A(net23),
    .B(net62),
    .Y(_04285_));
 sky130_fd_sc_hd__and4_1 _11511_ (.A(net23),
    .B(net12),
    .C(net61),
    .D(net62),
    .X(_04296_));
 sky130_fd_sc_hd__nand2_1 _11512_ (.A(net23),
    .B(net61),
    .Y(_04307_));
 sky130_fd_sc_hd__a22o_1 _11513_ (.A1(net23),
    .A2(net61),
    .B1(net62),
    .B2(net12),
    .X(_04318_));
 sky130_fd_sc_hd__o2bb2ai_1 _11514_ (.A1_N(_04012_),
    .A2_N(_04307_),
    .B1(_04285_),
    .B2(_04023_),
    .Y(_04329_));
 sky130_fd_sc_hd__o221ai_2 _11515_ (.A1(_01846_),
    .A2(_01890_),
    .B1(_04023_),
    .B2(_04285_),
    .C1(_04318_),
    .Y(_04340_));
 sky130_fd_sc_hd__nand3_1 _11516_ (.A(_04329_),
    .B(net63),
    .C(net1),
    .Y(_04351_));
 sky130_fd_sc_hd__o21ai_2 _11517_ (.A1(_01846_),
    .A2(_01890_),
    .B1(_04329_),
    .Y(_04362_));
 sky130_fd_sc_hd__o2111ai_4 _11518_ (.A1(_04023_),
    .A2(_04285_),
    .B1(net1),
    .C1(net63),
    .D1(_04318_),
    .Y(_04373_));
 sky130_fd_sc_hd__nand3b_2 _11519_ (.A_N(_04274_),
    .B(_04340_),
    .C(_04351_),
    .Y(_04384_));
 sky130_fd_sc_hd__nand3_2 _11520_ (.A(_04274_),
    .B(_04362_),
    .C(_04373_),
    .Y(_04395_));
 sky130_fd_sc_hd__a21oi_1 _11521_ (.A1(_04384_),
    .A2(_04395_),
    .B1(_04034_),
    .Y(_04406_));
 sky130_fd_sc_hd__a32o_1 _11522_ (.A1(net1),
    .A2(net61),
    .A3(_04001_),
    .B1(_04384_),
    .B2(_04395_),
    .X(_04417_));
 sky130_fd_sc_hd__and3_2 _11523_ (.A(_04384_),
    .B(_04395_),
    .C(_04034_),
    .X(_04428_));
 sky130_fd_sc_hd__nand3_2 _11524_ (.A(_04384_),
    .B(_04395_),
    .C(_04034_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_1 _11525_ (.A(_04417_),
    .B(_04439_),
    .Y(_04450_));
 sky130_fd_sc_hd__o21ai_2 _11526_ (.A1(_03782_),
    .A2(_03815_),
    .B1(_03804_),
    .Y(_04461_));
 sky130_fd_sc_hd__o22a_1 _11527_ (.A1(_03290_),
    .A2(_03793_),
    .B1(_03782_),
    .B2(_03815_),
    .X(_04472_));
 sky130_fd_sc_hd__nand2_1 _11528_ (.A(net55),
    .B(net29),
    .Y(_04483_));
 sky130_fd_sc_hd__a22oi_4 _11529_ (.A1(net44),
    .A2(net30),
    .B1(net31),
    .B2(net33),
    .Y(_04494_));
 sky130_fd_sc_hd__a22o_1 _11530_ (.A1(net44),
    .A2(net30),
    .B1(net31),
    .B2(net33),
    .X(_04505_));
 sky130_fd_sc_hd__and4_1 _11531_ (.A(net33),
    .B(net44),
    .C(net30),
    .D(net31),
    .X(_04515_));
 sky130_fd_sc_hd__nand4_2 _11532_ (.A(net33),
    .B(net44),
    .C(net30),
    .D(net31),
    .Y(_04526_));
 sky130_fd_sc_hd__o211ai_2 _11533_ (.A1(_01780_),
    .A2(_01857_),
    .B1(_04505_),
    .C1(_04526_),
    .Y(_04537_));
 sky130_fd_sc_hd__o21bai_1 _11534_ (.A1(_04494_),
    .A2(_04515_),
    .B1_N(_04483_),
    .Y(_04548_));
 sky130_fd_sc_hd__o22a_2 _11535_ (.A1(_01780_),
    .A2(_01857_),
    .B1(_04494_),
    .B2(_04515_),
    .X(_04559_));
 sky130_fd_sc_hd__a22o_1 _11536_ (.A1(net55),
    .A2(net29),
    .B1(_04505_),
    .B2(_04526_),
    .X(_04570_));
 sky130_fd_sc_hd__a41o_1 _11537_ (.A1(net33),
    .A2(net44),
    .A3(net30),
    .A4(net31),
    .B1(_04483_),
    .X(_04581_));
 sky130_fd_sc_hd__nand3_4 _11538_ (.A(_04472_),
    .B(_04537_),
    .C(_04548_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_4 _11539_ (.A1(_04494_),
    .A2(_04581_),
    .B1(_04461_),
    .Y(_04603_));
 sky130_fd_sc_hd__o211ai_2 _11540_ (.A1(_04494_),
    .A2(_04581_),
    .B1(_04461_),
    .C1(_04570_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2_1 _11541_ (.A(net26),
    .B(net60),
    .Y(_04625_));
 sky130_fd_sc_hd__and4_1 _11542_ (.A(net28),
    .B(net27),
    .C(net58),
    .D(net59),
    .X(_04636_));
 sky130_fd_sc_hd__nand4_2 _11543_ (.A(net28),
    .B(net27),
    .C(net58),
    .D(net59),
    .Y(_04647_));
 sky130_fd_sc_hd__a22oi_2 _11544_ (.A1(net28),
    .A2(net58),
    .B1(net59),
    .B2(net27),
    .Y(_04658_));
 sky130_fd_sc_hd__a22o_1 _11545_ (.A1(net28),
    .A2(net58),
    .B1(net59),
    .B2(net27),
    .X(_04669_));
 sky130_fd_sc_hd__and3_1 _11546_ (.A(_04625_),
    .B(_04647_),
    .C(_04669_),
    .X(_04680_));
 sky130_fd_sc_hd__o211ai_1 _11547_ (.A1(_01791_),
    .A2(_01835_),
    .B1(_04647_),
    .C1(_04669_),
    .Y(_04691_));
 sky130_fd_sc_hd__o211a_1 _11548_ (.A1(_04636_),
    .A2(_04658_),
    .B1(net26),
    .C1(net60),
    .X(_04702_));
 sky130_fd_sc_hd__a21o_1 _11549_ (.A1(_04647_),
    .A2(_04669_),
    .B1(_04625_),
    .X(_04713_));
 sky130_fd_sc_hd__o22a_1 _11550_ (.A1(_01791_),
    .A2(_01835_),
    .B1(_04636_),
    .B2(_04658_),
    .X(_04724_));
 sky130_fd_sc_hd__and4_1 _11551_ (.A(_04669_),
    .B(net60),
    .C(net26),
    .D(_04647_),
    .X(_04735_));
 sky130_fd_sc_hd__nand2_1 _11552_ (.A(_04691_),
    .B(_04713_),
    .Y(_04746_));
 sky130_fd_sc_hd__o2bb2ai_2 _11553_ (.A1_N(_04592_),
    .A2_N(_04614_),
    .B1(_04680_),
    .B2(_04702_),
    .Y(_04757_));
 sky130_fd_sc_hd__o221ai_4 _11554_ (.A1(_04559_),
    .A2(_04603_),
    .B1(_04724_),
    .B2(_04735_),
    .C1(_04592_),
    .Y(_04768_));
 sky130_fd_sc_hd__o2bb2ai_1 _11555_ (.A1_N(_04592_),
    .A2_N(_04614_),
    .B1(_04724_),
    .B2(_04735_),
    .Y(_04779_));
 sky130_fd_sc_hd__o211ai_2 _11556_ (.A1(_04603_),
    .A2(_04559_),
    .B1(_04592_),
    .C1(_04746_),
    .Y(_04790_));
 sky130_fd_sc_hd__nand2_1 _11557_ (.A(_04757_),
    .B(_04768_),
    .Y(_04801_));
 sky130_fd_sc_hd__a32oi_4 _11558_ (.A1(_03859_),
    .A2(_03870_),
    .A3(_03760_),
    .B1(_03727_),
    .B2(_03705_),
    .Y(_04812_));
 sky130_fd_sc_hd__a32oi_4 _11559_ (.A1(_03771_),
    .A2(_03837_),
    .A3(_03848_),
    .B1(_03913_),
    .B2(_03738_),
    .Y(_04822_));
 sky130_fd_sc_hd__o211ai_4 _11560_ (.A1(_03880_),
    .A2(_04812_),
    .B1(_04768_),
    .C1(_04757_),
    .Y(_04833_));
 sky130_fd_sc_hd__and3_1 _11561_ (.A(_04779_),
    .B(_04822_),
    .C(_04790_),
    .X(_04844_));
 sky130_fd_sc_hd__nand3_2 _11562_ (.A(_04779_),
    .B(_04822_),
    .C(_04790_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand3_1 _11563_ (.A(_04417_),
    .B(_04439_),
    .C(_04833_),
    .Y(_04866_));
 sky130_fd_sc_hd__a22o_1 _11564_ (.A1(_04417_),
    .A2(_04439_),
    .B1(_04833_),
    .B2(_04855_),
    .X(_04877_));
 sky130_fd_sc_hd__a21o_1 _11565_ (.A1(_04833_),
    .A2(_04855_),
    .B1(_04450_),
    .X(_04888_));
 sky130_fd_sc_hd__o211ai_2 _11566_ (.A1(_04406_),
    .A2(_04428_),
    .B1(_04833_),
    .C1(_04855_),
    .Y(_04899_));
 sky130_fd_sc_hd__a31oi_2 _11567_ (.A1(_03946_),
    .A2(_03628_),
    .A3(_03935_),
    .B1(_04100_),
    .Y(_04910_));
 sky130_fd_sc_hd__o22ai_2 _11568_ (.A1(_03924_),
    .A2(_03979_),
    .B1(_04111_),
    .B2(_03957_),
    .Y(_04921_));
 sky130_fd_sc_hd__o211ai_4 _11569_ (.A1(_03957_),
    .A2(_04910_),
    .B1(_04899_),
    .C1(_04888_),
    .Y(_04932_));
 sky130_fd_sc_hd__o211a_1 _11570_ (.A1(_04844_),
    .A2(_04866_),
    .B1(_04921_),
    .C1(_04877_),
    .X(_04943_));
 sky130_fd_sc_hd__o211ai_2 _11571_ (.A1(_04844_),
    .A2(_04866_),
    .B1(_04921_),
    .C1(_04877_),
    .Y(_04954_));
 sky130_fd_sc_hd__o2bb2ai_4 _11572_ (.A1_N(_04932_),
    .A2_N(_04954_),
    .B1(_04056_),
    .B2(_04067_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_1 _11573_ (.A(_04932_),
    .B(_04078_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand3_1 _11574_ (.A(_04932_),
    .B(_04954_),
    .C(_04078_),
    .Y(_04987_));
 sky130_fd_sc_hd__o21a_1 _11575_ (.A1(_04943_),
    .A2(_04976_),
    .B1(_04965_),
    .X(_04998_));
 sky130_fd_sc_hd__o21a_1 _11576_ (.A1(_03092_),
    .A2(_03103_),
    .B1(_04176_),
    .X(_05009_));
 sky130_fd_sc_hd__o21ai_2 _11577_ (.A1(_03092_),
    .A2(_03103_),
    .B1(_04176_),
    .Y(_05020_));
 sky130_fd_sc_hd__o21ai_2 _11578_ (.A1(_03114_),
    .A2(_04144_),
    .B1(_04176_),
    .Y(_05031_));
 sky130_fd_sc_hd__a22oi_2 _11579_ (.A1(_04965_),
    .A2(_04987_),
    .B1(_05020_),
    .B2(_04155_),
    .Y(_05042_));
 sky130_fd_sc_hd__o2bb2ai_2 _11580_ (.A1_N(_04965_),
    .A2_N(_04987_),
    .B1(_05009_),
    .B2(_04144_),
    .Y(_05053_));
 sky130_fd_sc_hd__o2111ai_4 _11581_ (.A1(_04943_),
    .A2(_04976_),
    .B1(_05020_),
    .C1(_04965_),
    .D1(_04155_),
    .Y(_05064_));
 sky130_fd_sc_hd__a32oi_4 _11582_ (.A1(_03531_),
    .A2(_04187_),
    .A3(_04198_),
    .B1(_05053_),
    .B2(_05064_),
    .Y(_05075_));
 sky130_fd_sc_hd__a32o_1 _11583_ (.A1(_03531_),
    .A2(_04187_),
    .A3(_04198_),
    .B1(_05053_),
    .B2(_05064_),
    .X(_05086_));
 sky130_fd_sc_hd__nor2_1 _11584_ (.A(_05042_),
    .B(_04231_),
    .Y(_05097_));
 sky130_fd_sc_hd__nand4_2 _11585_ (.A(_04187_),
    .B(_04198_),
    .C(_05053_),
    .D(_03531_),
    .Y(_05108_));
 sky130_fd_sc_hd__and4b_1 _11586_ (.A_N(_03039_),
    .B(_03509_),
    .C(_04187_),
    .D(_04198_),
    .X(_05119_));
 sky130_fd_sc_hd__o22ai_2 _11587_ (.A1(_03586_),
    .A2(_04209_),
    .B1(_05075_),
    .B2(_05097_),
    .Y(_05130_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(_05086_),
    .B(_05119_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _11589_ (.A(_05130_),
    .B(_04263_),
    .Y(_05152_));
 sky130_fd_sc_hd__a21oi_1 _11590_ (.A1(_05130_),
    .A2(_05141_),
    .B1(_04263_),
    .Y(_05163_));
 sky130_fd_sc_hd__a21oi_1 _11591_ (.A1(_04263_),
    .A2(_05130_),
    .B1(_05163_),
    .Y(net127));
 sky130_fd_sc_hd__a21oi_1 _11592_ (.A1(_04078_),
    .A2(_04932_),
    .B1(_04943_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21o_1 _11593_ (.A1(_04078_),
    .A2(_04932_),
    .B1(_04943_),
    .X(_05194_));
 sky130_fd_sc_hd__nand2_2 _11594_ (.A(net1),
    .B(net64),
    .Y(_05205_));
 sky130_fd_sc_hd__a31oi_4 _11595_ (.A1(_04274_),
    .A2(_04362_),
    .A3(_04373_),
    .B1(_04428_),
    .Y(_05216_));
 sky130_fd_sc_hd__a21o_1 _11596_ (.A1(_04395_),
    .A2(_04439_),
    .B1(_05205_),
    .X(_05227_));
 sky130_fd_sc_hd__a22o_1 _11597_ (.A1(net1),
    .A2(net64),
    .B1(_04395_),
    .B2(_04439_),
    .X(_05238_));
 sky130_fd_sc_hd__a311o_1 _11598_ (.A1(_04274_),
    .A2(_04362_),
    .A3(_04373_),
    .B1(_05205_),
    .C1(_04428_),
    .X(_05249_));
 sky130_fd_sc_hd__nand2_2 _11599_ (.A(_05238_),
    .B(_05249_),
    .Y(_05260_));
 sky130_fd_sc_hd__o21ai_1 _11600_ (.A1(_04406_),
    .A2(_04428_),
    .B1(_04855_),
    .Y(_05271_));
 sky130_fd_sc_hd__o21ai_2 _11601_ (.A1(_04801_),
    .A2(_04822_),
    .B1(_05271_),
    .Y(_05282_));
 sky130_fd_sc_hd__a21boi_1 _11602_ (.A1(_04450_),
    .A2(_04855_),
    .B1_N(_04833_),
    .Y(_05293_));
 sky130_fd_sc_hd__o21ai_2 _11603_ (.A1(_04625_),
    .A2(_04658_),
    .B1(_04647_),
    .Y(_05304_));
 sky130_fd_sc_hd__nand2_1 _11604_ (.A(net26),
    .B(net61),
    .Y(_05315_));
 sky130_fd_sc_hd__a22o_2 _11605_ (.A1(net26),
    .A2(net61),
    .B1(net62),
    .B2(net23),
    .X(_05326_));
 sky130_fd_sc_hd__nand2_1 _11606_ (.A(net26),
    .B(net62),
    .Y(_05337_));
 sky130_fd_sc_hd__and4_1 _11607_ (.A(net26),
    .B(net23),
    .C(net61),
    .D(net62),
    .X(_05348_));
 sky130_fd_sc_hd__nand4_1 _11608_ (.A(net26),
    .B(net23),
    .C(net61),
    .D(net62),
    .Y(_05359_));
 sky130_fd_sc_hd__a22oi_1 _11609_ (.A1(net12),
    .A2(net63),
    .B1(_05326_),
    .B2(_05359_),
    .Y(_05370_));
 sky130_fd_sc_hd__a22o_1 _11610_ (.A1(net12),
    .A2(net63),
    .B1(_05326_),
    .B2(_05359_),
    .X(_05381_));
 sky130_fd_sc_hd__o2111a_1 _11611_ (.A1(_04307_),
    .A2(_05337_),
    .B1(net12),
    .C1(net63),
    .D1(_05326_),
    .X(_05392_));
 sky130_fd_sc_hd__o2111ai_4 _11612_ (.A1(_04307_),
    .A2(_05337_),
    .B1(net12),
    .C1(net63),
    .D1(_05326_),
    .Y(_05403_));
 sky130_fd_sc_hd__o21bai_2 _11613_ (.A1(_05370_),
    .A2(_05392_),
    .B1_N(_05304_),
    .Y(_05414_));
 sky130_fd_sc_hd__nand3_4 _11614_ (.A(_05381_),
    .B(_05403_),
    .C(_05304_),
    .Y(_05425_));
 sky130_fd_sc_hd__inv_2 _11615_ (.A(_05425_),
    .Y(_05436_));
 sky130_fd_sc_hd__a31o_1 _11616_ (.A1(_04318_),
    .A2(net63),
    .A3(net1),
    .B1(_04296_),
    .X(_05447_));
 sky130_fd_sc_hd__a21oi_2 _11617_ (.A1(_05414_),
    .A2(_05425_),
    .B1(_05447_),
    .Y(_05458_));
 sky130_fd_sc_hd__a21o_1 _11618_ (.A1(_05414_),
    .A2(_05425_),
    .B1(_05447_),
    .X(_05469_));
 sky130_fd_sc_hd__and3_2 _11619_ (.A(_05414_),
    .B(_05425_),
    .C(_05447_),
    .X(_05480_));
 sky130_fd_sc_hd__nand3_1 _11620_ (.A(_05414_),
    .B(_05425_),
    .C(_05447_),
    .Y(_05491_));
 sky130_fd_sc_hd__nand2_1 _11621_ (.A(_05469_),
    .B(_05491_),
    .Y(_05502_));
 sky130_fd_sc_hd__o21ai_2 _11622_ (.A1(_04483_),
    .A2(_04494_),
    .B1(_04526_),
    .Y(_05513_));
 sky130_fd_sc_hd__o21a_1 _11623_ (.A1(_04483_),
    .A2(_04494_),
    .B1(_04526_),
    .X(_05523_));
 sky130_fd_sc_hd__nand2_1 _11624_ (.A(net55),
    .B(net30),
    .Y(_05534_));
 sky130_fd_sc_hd__a22oi_4 _11625_ (.A1(net44),
    .A2(net31),
    .B1(net32),
    .B2(net33),
    .Y(_05545_));
 sky130_fd_sc_hd__a22o_1 _11626_ (.A1(net44),
    .A2(net31),
    .B1(net32),
    .B2(net33),
    .X(_05556_));
 sky130_fd_sc_hd__and4_1 _11627_ (.A(net33),
    .B(net44),
    .C(net31),
    .D(net32),
    .X(_05567_));
 sky130_fd_sc_hd__nand4_2 _11628_ (.A(net33),
    .B(net44),
    .C(net31),
    .D(net32),
    .Y(_05578_));
 sky130_fd_sc_hd__o211ai_4 _11629_ (.A1(_01780_),
    .A2(_01868_),
    .B1(_05556_),
    .C1(_05578_),
    .Y(_05589_));
 sky130_fd_sc_hd__o21bai_4 _11630_ (.A1(_05545_),
    .A2(_05567_),
    .B1_N(_05534_),
    .Y(_05600_));
 sky130_fd_sc_hd__o22a_2 _11631_ (.A1(_01780_),
    .A2(_01868_),
    .B1(_05545_),
    .B2(_05567_),
    .X(_05611_));
 sky130_fd_sc_hd__o21ai_1 _11632_ (.A1(_05545_),
    .A2(_05567_),
    .B1(_05534_),
    .Y(_05622_));
 sky130_fd_sc_hd__a41o_1 _11633_ (.A1(net33),
    .A2(net44),
    .A3(net31),
    .A4(net32),
    .B1(_05534_),
    .X(_05633_));
 sky130_fd_sc_hd__nand3_4 _11634_ (.A(_05523_),
    .B(_05589_),
    .C(_05600_),
    .Y(_05644_));
 sky130_fd_sc_hd__o21ai_4 _11635_ (.A1(_05545_),
    .A2(_05633_),
    .B1(_05513_),
    .Y(_05655_));
 sky130_fd_sc_hd__o211a_1 _11636_ (.A1(_05545_),
    .A2(_05633_),
    .B1(_05513_),
    .C1(_05622_),
    .X(_05666_));
 sky130_fd_sc_hd__o211ai_2 _11637_ (.A1(_05545_),
    .A2(_05633_),
    .B1(_05513_),
    .C1(_05622_),
    .Y(_05677_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(net27),
    .B(net60),
    .Y(_05688_));
 sky130_fd_sc_hd__nand4_4 _11639_ (.A(net28),
    .B(net58),
    .C(net59),
    .D(net29),
    .Y(_05699_));
 sky130_fd_sc_hd__a22oi_1 _11640_ (.A1(net28),
    .A2(net59),
    .B1(net29),
    .B2(net58),
    .Y(_05710_));
 sky130_fd_sc_hd__a22o_1 _11641_ (.A1(net28),
    .A2(net59),
    .B1(net29),
    .B2(net58),
    .X(_05721_));
 sky130_fd_sc_hd__and3_1 _11642_ (.A(_05688_),
    .B(_05699_),
    .C(_05721_),
    .X(_05732_));
 sky130_fd_sc_hd__o211ai_4 _11643_ (.A1(_01769_),
    .A2(_01835_),
    .B1(_05699_),
    .C1(_05721_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21oi_2 _11644_ (.A1(_05699_),
    .A2(_05721_),
    .B1(_05688_),
    .Y(_05754_));
 sky130_fd_sc_hd__a21o_2 _11645_ (.A1(_05699_),
    .A2(_05721_),
    .B1(_05688_),
    .X(_05765_));
 sky130_fd_sc_hd__nand2_1 _11646_ (.A(_05743_),
    .B(_05765_),
    .Y(_05776_));
 sky130_fd_sc_hd__o2bb2ai_2 _11647_ (.A1_N(_05644_),
    .A2_N(_05677_),
    .B1(_05732_),
    .B2(_05754_),
    .Y(_05787_));
 sky130_fd_sc_hd__o2111ai_4 _11648_ (.A1(_05611_),
    .A2(_05655_),
    .B1(_05743_),
    .C1(_05765_),
    .D1(_05644_),
    .Y(_05798_));
 sky130_fd_sc_hd__a21o_1 _11649_ (.A1(_05644_),
    .A2(_05677_),
    .B1(_05776_),
    .X(_05809_));
 sky130_fd_sc_hd__o221ai_4 _11650_ (.A1(_05611_),
    .A2(_05655_),
    .B1(_05732_),
    .B2(_05754_),
    .C1(_05644_),
    .Y(_05820_));
 sky130_fd_sc_hd__a2bb2oi_2 _11651_ (.A1_N(_04603_),
    .A2_N(_04559_),
    .B1(_04592_),
    .B2(_04746_),
    .Y(_05831_));
 sky130_fd_sc_hd__o2bb2ai_2 _11652_ (.A1_N(_04592_),
    .A2_N(_04746_),
    .B1(_04603_),
    .B2(_04559_),
    .Y(_05842_));
 sky130_fd_sc_hd__a21oi_2 _11653_ (.A1(_05787_),
    .A2(_05798_),
    .B1(_05831_),
    .Y(_05853_));
 sky130_fd_sc_hd__nand3_4 _11654_ (.A(_05809_),
    .B(_05820_),
    .C(_05842_),
    .Y(_05864_));
 sky130_fd_sc_hd__a21oi_2 _11655_ (.A1(_05809_),
    .A2(_05820_),
    .B1(_05842_),
    .Y(_05874_));
 sky130_fd_sc_hd__nand3_1 _11656_ (.A(_05831_),
    .B(_05798_),
    .C(_05787_),
    .Y(_05885_));
 sky130_fd_sc_hd__a21o_1 _11657_ (.A1(_05864_),
    .A2(_05885_),
    .B1(_05502_),
    .X(_05896_));
 sky130_fd_sc_hd__o211ai_2 _11658_ (.A1(_05458_),
    .A2(_05480_),
    .B1(_05864_),
    .C1(_05885_),
    .Y(_05907_));
 sky130_fd_sc_hd__a311oi_2 _11659_ (.A1(_05787_),
    .A2(_05831_),
    .A3(_05798_),
    .B1(_05458_),
    .C1(_05480_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand4_1 _11660_ (.A(_05469_),
    .B(_05491_),
    .C(_05864_),
    .D(_05885_),
    .Y(_05929_));
 sky130_fd_sc_hd__inv_2 _11661_ (.A(_05929_),
    .Y(_05940_));
 sky130_fd_sc_hd__o22ai_1 _11662_ (.A1(_05458_),
    .A2(_05480_),
    .B1(_05853_),
    .B2(_05874_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_05293_),
    .B(_05951_),
    .Y(_05962_));
 sky130_fd_sc_hd__nand3_1 _11664_ (.A(_05293_),
    .B(_05929_),
    .C(_05951_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand3_4 _11665_ (.A(_05896_),
    .B(_05907_),
    .C(_05282_),
    .Y(_05984_));
 sky130_fd_sc_hd__a22o_1 _11666_ (.A1(_05238_),
    .A2(_05249_),
    .B1(_05973_),
    .B2(_05984_),
    .X(_05995_));
 sky130_fd_sc_hd__nand4_1 _11667_ (.A(_05238_),
    .B(_05249_),
    .C(_05973_),
    .D(_05984_),
    .Y(_06006_));
 sky130_fd_sc_hd__and3_1 _11668_ (.A(_05973_),
    .B(_05984_),
    .C(_05260_),
    .X(_06017_));
 sky130_fd_sc_hd__o211ai_2 _11669_ (.A1(_05940_),
    .A2(_05962_),
    .B1(_05984_),
    .C1(_05260_),
    .Y(_06028_));
 sky130_fd_sc_hd__a21o_1 _11670_ (.A1(_05973_),
    .A2(_05984_),
    .B1(_05260_),
    .X(_06039_));
 sky130_fd_sc_hd__nand2_1 _11671_ (.A(_05194_),
    .B(_06039_),
    .Y(_06050_));
 sky130_fd_sc_hd__and3_1 _11672_ (.A(_05194_),
    .B(_06028_),
    .C(_06039_),
    .X(_06061_));
 sky130_fd_sc_hd__nand3_2 _11673_ (.A(_05194_),
    .B(_06028_),
    .C(_06039_),
    .Y(_06072_));
 sky130_fd_sc_hd__nand3_1 _11674_ (.A(_05995_),
    .B(_06006_),
    .C(_05183_),
    .Y(_06083_));
 sky130_fd_sc_hd__a22oi_4 _11675_ (.A1(_04998_),
    .A2(_05031_),
    .B1(_06072_),
    .B2(_06083_),
    .Y(_06094_));
 sky130_fd_sc_hd__a31oi_2 _11676_ (.A1(_05183_),
    .A2(_05995_),
    .A3(_06006_),
    .B1(_05064_),
    .Y(_06105_));
 sky130_fd_sc_hd__and4_1 _11677_ (.A(_06072_),
    .B(_06083_),
    .C(_04998_),
    .D(_05031_),
    .X(_06116_));
 sky130_fd_sc_hd__o21ai_2 _11678_ (.A1(_06017_),
    .A2(_06050_),
    .B1(_06105_),
    .Y(_06127_));
 sky130_fd_sc_hd__a21oi_1 _11679_ (.A1(_06105_),
    .A2(_06072_),
    .B1(_06094_),
    .Y(_06138_));
 sky130_fd_sc_hd__a21o_1 _11680_ (.A1(_06105_),
    .A2(_06072_),
    .B1(_06094_),
    .X(_06149_));
 sky130_fd_sc_hd__o22a_1 _11681_ (.A1(_05042_),
    .A2(_04231_),
    .B1(_04209_),
    .B2(_03586_),
    .X(_06160_));
 sky130_fd_sc_hd__o221ai_2 _11682_ (.A1(_05097_),
    .A2(_05119_),
    .B1(_06094_),
    .B2(_06116_),
    .C1(_05086_),
    .Y(_06171_));
 sky130_fd_sc_hd__o21ai_1 _11683_ (.A1(_05075_),
    .A2(_06160_),
    .B1(_06138_),
    .Y(_06182_));
 sky130_fd_sc_hd__nor2_1 _11684_ (.A(_06094_),
    .B(_05108_),
    .Y(_06193_));
 sky130_fd_sc_hd__and3_1 _11685_ (.A(_06138_),
    .B(_05086_),
    .C(_05119_),
    .X(_06204_));
 sky130_fd_sc_hd__o31a_1 _11686_ (.A1(_05075_),
    .A2(_06138_),
    .A3(_06160_),
    .B1(_06182_),
    .X(_06215_));
 sky130_fd_sc_hd__a21oi_1 _11687_ (.A1(_06171_),
    .A2(_06182_),
    .B1(_05152_),
    .Y(_06225_));
 sky130_fd_sc_hd__o2bb2ai_1 _11688_ (.A1_N(_05260_),
    .A2_N(_05984_),
    .B1(_05940_),
    .B2(_05962_),
    .Y(_06236_));
 sky130_fd_sc_hd__a21boi_2 _11689_ (.A1(_05260_),
    .A2(_05984_),
    .B1_N(_05973_),
    .Y(_06247_));
 sky130_fd_sc_hd__o31a_1 _11690_ (.A1(_05458_),
    .A2(_05480_),
    .A3(_05874_),
    .B1(_05864_),
    .X(_06258_));
 sky130_fd_sc_hd__o21ai_1 _11691_ (.A1(_05688_),
    .A2(_05710_),
    .B1(_05699_),
    .Y(_06269_));
 sky130_fd_sc_hd__o21a_1 _11692_ (.A1(_05688_),
    .A2(_05710_),
    .B1(_05699_),
    .X(_06280_));
 sky130_fd_sc_hd__nand2_1 _11693_ (.A(net27),
    .B(net62),
    .Y(_06291_));
 sky130_fd_sc_hd__and4_1 _11694_ (.A(net27),
    .B(net26),
    .C(net61),
    .D(net62),
    .X(_06302_));
 sky130_fd_sc_hd__nand2_2 _11695_ (.A(net27),
    .B(net61),
    .Y(_06313_));
 sky130_fd_sc_hd__a22o_1 _11696_ (.A1(net27),
    .A2(net61),
    .B1(net62),
    .B2(net26),
    .X(_06324_));
 sky130_fd_sc_hd__o2bb2ai_1 _11697_ (.A1_N(_05337_),
    .A2_N(_06313_),
    .B1(_06291_),
    .B2(_05315_),
    .Y(_06335_));
 sky130_fd_sc_hd__o221ai_1 _11698_ (.A1(_01802_),
    .A2(_01890_),
    .B1(_05315_),
    .B2(_06291_),
    .C1(_06324_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand3_1 _11699_ (.A(_06335_),
    .B(net63),
    .C(net23),
    .Y(_06357_));
 sky130_fd_sc_hd__o21ai_1 _11700_ (.A1(_01802_),
    .A2(_01890_),
    .B1(_06335_),
    .Y(_06368_));
 sky130_fd_sc_hd__o2111ai_1 _11701_ (.A1(_05315_),
    .A2(_06291_),
    .B1(net23),
    .C1(net63),
    .D1(_06324_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand3_1 _11702_ (.A(_06280_),
    .B(_06346_),
    .C(_06357_),
    .Y(_06390_));
 sky130_fd_sc_hd__nand3_2 _11703_ (.A(_06368_),
    .B(_06379_),
    .C(_06269_),
    .Y(_06401_));
 sky130_fd_sc_hd__and3_1 _11704_ (.A(_05326_),
    .B(net63),
    .C(net12),
    .X(_06412_));
 sky130_fd_sc_hd__a31o_1 _11705_ (.A1(_05326_),
    .A2(net63),
    .A3(net12),
    .B1(_05348_),
    .X(_06423_));
 sky130_fd_sc_hd__a21oi_1 _11706_ (.A1(_06390_),
    .A2(_06401_),
    .B1(_06423_),
    .Y(_06434_));
 sky130_fd_sc_hd__a211o_1 _11707_ (.A1(_06390_),
    .A2(_06401_),
    .B1(_06412_),
    .C1(_05348_),
    .X(_06445_));
 sky130_fd_sc_hd__o21a_1 _11708_ (.A1(_05348_),
    .A2(_06412_),
    .B1(_06390_),
    .X(_06456_));
 sky130_fd_sc_hd__nand3_1 _11709_ (.A(_06390_),
    .B(_06401_),
    .C(_06423_),
    .Y(_06467_));
 sky130_fd_sc_hd__a21oi_1 _11710_ (.A1(_06456_),
    .A2(_06401_),
    .B1(_06434_),
    .Y(_06478_));
 sky130_fd_sc_hd__a21o_1 _11711_ (.A1(_06456_),
    .A2(_06401_),
    .B1(_06434_),
    .X(_06489_));
 sky130_fd_sc_hd__o21ai_1 _11712_ (.A1(_01780_),
    .A2(_01868_),
    .B1(_05578_),
    .Y(_06500_));
 sky130_fd_sc_hd__o21ai_1 _11713_ (.A1(_05534_),
    .A2(_05545_),
    .B1(_05578_),
    .Y(_06511_));
 sky130_fd_sc_hd__o21a_1 _11714_ (.A1(_05534_),
    .A2(_05545_),
    .B1(_05578_),
    .X(_06522_));
 sky130_fd_sc_hd__nand2_1 _11715_ (.A(net55),
    .B(net31),
    .Y(_06533_));
 sky130_fd_sc_hd__a22oi_4 _11716_ (.A1(net33),
    .A2(net2),
    .B1(net32),
    .B2(net44),
    .Y(_06544_));
 sky130_fd_sc_hd__a22o_1 _11717_ (.A1(net33),
    .A2(net2),
    .B1(net32),
    .B2(net44),
    .X(_06555_));
 sky130_fd_sc_hd__and4_1 _11718_ (.A(net33),
    .B(net44),
    .C(net2),
    .D(net32),
    .X(_06566_));
 sky130_fd_sc_hd__nand4_4 _11719_ (.A(net33),
    .B(net44),
    .C(net2),
    .D(net32),
    .Y(_06577_));
 sky130_fd_sc_hd__o211ai_2 _11720_ (.A1(_01780_),
    .A2(_01879_),
    .B1(_06555_),
    .C1(_06577_),
    .Y(_06588_));
 sky130_fd_sc_hd__o21bai_1 _11721_ (.A1(_06544_),
    .A2(_06566_),
    .B1_N(_06533_),
    .Y(_06599_));
 sky130_fd_sc_hd__o22a_2 _11722_ (.A1(_01780_),
    .A2(_01879_),
    .B1(_06544_),
    .B2(_06566_),
    .X(_06609_));
 sky130_fd_sc_hd__o22ai_1 _11723_ (.A1(_01780_),
    .A2(_01879_),
    .B1(_06544_),
    .B2(_06566_),
    .Y(_06620_));
 sky130_fd_sc_hd__nand4_2 _11724_ (.A(_06555_),
    .B(_06577_),
    .C(net55),
    .D(net31),
    .Y(_06631_));
 sky130_fd_sc_hd__a22oi_1 _11725_ (.A1(_05556_),
    .A2(_06500_),
    .B1(_06620_),
    .B2(_06631_),
    .Y(_06642_));
 sky130_fd_sc_hd__nand3_4 _11726_ (.A(_06522_),
    .B(_06588_),
    .C(_06599_),
    .Y(_06653_));
 sky130_fd_sc_hd__nand2_2 _11727_ (.A(_06511_),
    .B(_06631_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand3_1 _11728_ (.A(_06620_),
    .B(_06631_),
    .C(_06511_),
    .Y(_06675_));
 sky130_fd_sc_hd__nand2_1 _11729_ (.A(net28),
    .B(net60),
    .Y(_06686_));
 sky130_fd_sc_hd__a22oi_4 _11730_ (.A1(net59),
    .A2(net29),
    .B1(net30),
    .B2(net58),
    .Y(_06697_));
 sky130_fd_sc_hd__a22o_1 _11731_ (.A1(net59),
    .A2(net29),
    .B1(net30),
    .B2(net58),
    .X(_06708_));
 sky130_fd_sc_hd__and4_1 _11732_ (.A(net58),
    .B(net59),
    .C(net29),
    .D(net30),
    .X(_06719_));
 sky130_fd_sc_hd__nand4_2 _11733_ (.A(net58),
    .B(net59),
    .C(net29),
    .D(net30),
    .Y(_06730_));
 sky130_fd_sc_hd__and3_1 _11734_ (.A(_06686_),
    .B(_06708_),
    .C(_06730_),
    .X(_06741_));
 sky130_fd_sc_hd__o211ai_1 _11735_ (.A1(_01748_),
    .A2(_01835_),
    .B1(_06708_),
    .C1(_06730_),
    .Y(_06752_));
 sky130_fd_sc_hd__o211a_1 _11736_ (.A1(_06697_),
    .A2(_06719_),
    .B1(net28),
    .C1(net60),
    .X(_06763_));
 sky130_fd_sc_hd__o21bai_1 _11737_ (.A1(_06697_),
    .A2(_06719_),
    .B1_N(_06686_),
    .Y(_06774_));
 sky130_fd_sc_hd__o22a_1 _11738_ (.A1(_01748_),
    .A2(_01835_),
    .B1(_06697_),
    .B2(_06719_),
    .X(_06785_));
 sky130_fd_sc_hd__o21ai_1 _11739_ (.A1(_06697_),
    .A2(_06719_),
    .B1(_06686_),
    .Y(_06796_));
 sky130_fd_sc_hd__and4_1 _11740_ (.A(_06708_),
    .B(_06730_),
    .C(net28),
    .D(net60),
    .X(_06807_));
 sky130_fd_sc_hd__nand4_1 _11741_ (.A(_06708_),
    .B(_06730_),
    .C(net28),
    .D(net60),
    .Y(_06818_));
 sky130_fd_sc_hd__nand2_1 _11742_ (.A(_06796_),
    .B(_06818_),
    .Y(_06829_));
 sky130_fd_sc_hd__nand2_1 _11743_ (.A(_06752_),
    .B(_06774_),
    .Y(_06840_));
 sky130_fd_sc_hd__o221a_2 _11744_ (.A1(_06741_),
    .A2(_06763_),
    .B1(_06609_),
    .B2(_06664_),
    .C1(_06653_),
    .X(_06851_));
 sky130_fd_sc_hd__o221ai_4 _11745_ (.A1(_06741_),
    .A2(_06763_),
    .B1(_06609_),
    .B2(_06664_),
    .C1(_06653_),
    .Y(_06862_));
 sky130_fd_sc_hd__o2bb2ai_2 _11746_ (.A1_N(_06653_),
    .A2_N(_06675_),
    .B1(_06785_),
    .B2(_06807_),
    .Y(_06873_));
 sky130_fd_sc_hd__o221ai_4 _11747_ (.A1(_06785_),
    .A2(_06807_),
    .B1(_06609_),
    .B2(_06664_),
    .C1(_06653_),
    .Y(_06884_));
 sky130_fd_sc_hd__o2bb2ai_1 _11748_ (.A1_N(_06653_),
    .A2_N(_06675_),
    .B1(_06741_),
    .B2(_06763_),
    .Y(_06895_));
 sky130_fd_sc_hd__a32oi_4 _11749_ (.A1(_05523_),
    .A2(_05589_),
    .A3(_05600_),
    .B1(_05743_),
    .B2(_05765_),
    .Y(_06906_));
 sky130_fd_sc_hd__a2bb2oi_1 _11750_ (.A1_N(_05655_),
    .A2_N(_05611_),
    .B1(_05644_),
    .B2(_05776_),
    .Y(_06917_));
 sky130_fd_sc_hd__nand3_4 _11751_ (.A(_06917_),
    .B(_06895_),
    .C(_06884_),
    .Y(_06928_));
 sky130_fd_sc_hd__o21ai_4 _11752_ (.A1(_05666_),
    .A2(_06906_),
    .B1(_06873_),
    .Y(_06939_));
 sky130_fd_sc_hd__o211a_1 _11753_ (.A1(_05666_),
    .A2(_06906_),
    .B1(_06873_),
    .C1(_06862_),
    .X(_06950_));
 sky130_fd_sc_hd__o211ai_2 _11754_ (.A1(_05666_),
    .A2(_06906_),
    .B1(_06873_),
    .C1(_06862_),
    .Y(_06961_));
 sky130_fd_sc_hd__o211ai_4 _11755_ (.A1(_06851_),
    .A2(_06939_),
    .B1(_06928_),
    .C1(_06489_),
    .Y(_06971_));
 sky130_fd_sc_hd__a21o_1 _11756_ (.A1(_06928_),
    .A2(_06961_),
    .B1(_06489_),
    .X(_06982_));
 sky130_fd_sc_hd__a22o_1 _11757_ (.A1(_06445_),
    .A2(_06467_),
    .B1(_06928_),
    .B2(_06961_),
    .X(_06993_));
 sky130_fd_sc_hd__nand2_1 _11758_ (.A(_06478_),
    .B(_06928_),
    .Y(_07004_));
 sky130_fd_sc_hd__o221ai_4 _11759_ (.A1(_06950_),
    .A2(_07004_),
    .B1(_05853_),
    .B2(_05918_),
    .C1(_06993_),
    .Y(_07015_));
 sky130_fd_sc_hd__o2111a_1 _11760_ (.A1(_05874_),
    .A2(_05502_),
    .B1(_05864_),
    .C1(_06971_),
    .D1(_06982_),
    .X(_07026_));
 sky130_fd_sc_hd__o2111ai_4 _11761_ (.A1(_05874_),
    .A2(_05502_),
    .B1(_05864_),
    .C1(_06971_),
    .D1(_06982_),
    .Y(_07037_));
 sky130_fd_sc_hd__a22oi_2 _11762_ (.A1(net12),
    .A2(net64),
    .B1(net34),
    .B2(net1),
    .Y(_07048_));
 sky130_fd_sc_hd__and4_2 _11763_ (.A(net12),
    .B(net1),
    .C(net64),
    .D(net34),
    .X(_07059_));
 sky130_fd_sc_hd__nand4_1 _11764_ (.A(net12),
    .B(net1),
    .C(net64),
    .D(net34),
    .Y(_07070_));
 sky130_fd_sc_hd__nor2_1 _11765_ (.A(_07048_),
    .B(_07059_),
    .Y(_07081_));
 sky130_fd_sc_hd__a31o_1 _11766_ (.A1(_05304_),
    .A2(_05381_),
    .A3(_05403_),
    .B1(_05480_),
    .X(_07092_));
 sky130_fd_sc_hd__o21a_1 _11767_ (.A1(_05436_),
    .A2(_05480_),
    .B1(_07081_),
    .X(_07103_));
 sky130_fd_sc_hd__o211a_1 _11768_ (.A1(_07048_),
    .A2(_07059_),
    .B1(_05425_),
    .C1(_05491_),
    .X(_07114_));
 sky130_fd_sc_hd__o22a_1 _11769_ (.A1(_05436_),
    .A2(_05480_),
    .B1(_07048_),
    .B2(_07059_),
    .X(_07125_));
 sky130_fd_sc_hd__and3_1 _11770_ (.A(_05425_),
    .B(_05491_),
    .C(_07081_),
    .X(_07136_));
 sky130_fd_sc_hd__nor2_1 _11771_ (.A(_07125_),
    .B(_07136_),
    .Y(_07147_));
 sky130_fd_sc_hd__o2bb2ai_2 _11772_ (.A1_N(_07015_),
    .A2_N(_07037_),
    .B1(_07125_),
    .B2(_07136_),
    .Y(_07158_));
 sky130_fd_sc_hd__o211ai_4 _11773_ (.A1(_07103_),
    .A2(_07114_),
    .B1(_07015_),
    .C1(_07037_),
    .Y(_07169_));
 sky130_fd_sc_hd__o2bb2ai_1 _11774_ (.A1_N(_07015_),
    .A2_N(_07037_),
    .B1(_07103_),
    .B2(_07114_),
    .Y(_07180_));
 sky130_fd_sc_hd__o21ai_1 _11775_ (.A1(_07125_),
    .A2(_07136_),
    .B1(_07037_),
    .Y(_07191_));
 sky130_fd_sc_hd__o211ai_1 _11776_ (.A1(_07125_),
    .A2(_07136_),
    .B1(_07015_),
    .C1(_07037_),
    .Y(_07202_));
 sky130_fd_sc_hd__and3_2 _11777_ (.A(_07180_),
    .B(_07202_),
    .C(_06236_),
    .X(_07213_));
 sky130_fd_sc_hd__nand3_2 _11778_ (.A(_07180_),
    .B(_07202_),
    .C(_06236_),
    .Y(_07224_));
 sky130_fd_sc_hd__nand3_4 _11779_ (.A(_06247_),
    .B(_07158_),
    .C(_07169_),
    .Y(_07235_));
 sky130_fd_sc_hd__a31oi_1 _11780_ (.A1(_06247_),
    .A2(_07158_),
    .A3(_07169_),
    .B1(_05227_),
    .Y(_07246_));
 sky130_fd_sc_hd__a31o_1 _11781_ (.A1(_06247_),
    .A2(_07158_),
    .A3(_07169_),
    .B1(_05227_),
    .X(_07257_));
 sky130_fd_sc_hd__nand3b_1 _11782_ (.A_N(_05227_),
    .B(_07224_),
    .C(_07235_),
    .Y(_07268_));
 sky130_fd_sc_hd__o2bb2ai_2 _11783_ (.A1_N(_07224_),
    .A2_N(_07235_),
    .B1(_05205_),
    .B2(_05216_),
    .Y(_07279_));
 sky130_fd_sc_hd__a21o_1 _11784_ (.A1(_07224_),
    .A2(_07235_),
    .B1(_05227_),
    .X(_07290_));
 sky130_fd_sc_hd__o211ai_2 _11785_ (.A1(_05205_),
    .A2(_05216_),
    .B1(_07224_),
    .C1(_07235_),
    .Y(_07301_));
 sky130_fd_sc_hd__o211a_1 _11786_ (.A1(_07213_),
    .A2(_07257_),
    .B1(_06061_),
    .C1(_07279_),
    .X(_07312_));
 sky130_fd_sc_hd__o211ai_4 _11787_ (.A1(_07213_),
    .A2(_07257_),
    .B1(_07279_),
    .C1(_06061_),
    .Y(_07323_));
 sky130_fd_sc_hd__a2bb2oi_2 _11788_ (.A1_N(_06017_),
    .A2_N(_06050_),
    .B1(_07268_),
    .B2(_07279_),
    .Y(_07334_));
 sky130_fd_sc_hd__o211ai_2 _11789_ (.A1(_06050_),
    .A2(_06017_),
    .B1(_07301_),
    .C1(_07290_),
    .Y(_07344_));
 sky130_fd_sc_hd__nand2_1 _11790_ (.A(_07323_),
    .B(_07344_),
    .Y(_07355_));
 sky130_fd_sc_hd__o2111a_1 _11791_ (.A1(_05108_),
    .A2(_06094_),
    .B1(_06127_),
    .C1(_07323_),
    .D1(_07344_),
    .X(_07366_));
 sky130_fd_sc_hd__o2111ai_1 _11792_ (.A1(_05108_),
    .A2(_06094_),
    .B1(_06127_),
    .C1(_07323_),
    .D1(_07344_),
    .Y(_07377_));
 sky130_fd_sc_hd__o22a_1 _11793_ (.A1(_06116_),
    .A2(_06193_),
    .B1(_07312_),
    .B2(_07334_),
    .X(_07388_));
 sky130_fd_sc_hd__o22ai_1 _11794_ (.A1(_06116_),
    .A2(_06193_),
    .B1(_07312_),
    .B2(_07334_),
    .Y(_07399_));
 sky130_fd_sc_hd__o21ai_1 _11795_ (.A1(_07366_),
    .A2(_07388_),
    .B1(_06204_),
    .Y(_07410_));
 sky130_fd_sc_hd__o211a_1 _11796_ (.A1(_05141_),
    .A2(_06149_),
    .B1(_07377_),
    .C1(_07399_),
    .X(_07421_));
 sky130_fd_sc_hd__o211ai_1 _11797_ (.A1(_05141_),
    .A2(_06149_),
    .B1(_07377_),
    .C1(_07399_),
    .Y(_07432_));
 sky130_fd_sc_hd__o2bb2a_1 _11798_ (.A1_N(_07410_),
    .A2_N(_07432_),
    .B1(_05152_),
    .B2(_06215_),
    .X(_07443_));
 sky130_fd_sc_hd__nand2_1 _11799_ (.A(_07432_),
    .B(_06225_),
    .Y(_07454_));
 sky130_fd_sc_hd__a21oi_1 _11800_ (.A1(_06225_),
    .A2(_07432_),
    .B1(_07443_),
    .Y(net66));
 sky130_fd_sc_hd__or3_1 _11801_ (.A(_05108_),
    .B(_06094_),
    .C(_07334_),
    .X(_07475_));
 sky130_fd_sc_hd__o21ai_1 _11802_ (.A1(_05205_),
    .A2(_05216_),
    .B1(_07224_),
    .Y(_07486_));
 sky130_fd_sc_hd__a32oi_2 _11803_ (.A1(_06258_),
    .A2(_06971_),
    .A3(_06982_),
    .B1(_07015_),
    .B2(_07147_),
    .Y(_07497_));
 sky130_fd_sc_hd__o21ai_2 _11804_ (.A1(_06533_),
    .A2(_06544_),
    .B1(_06577_),
    .Y(_07508_));
 sky130_fd_sc_hd__o21a_1 _11805_ (.A1(_06533_),
    .A2(_06544_),
    .B1(_06577_),
    .X(_07519_));
 sky130_fd_sc_hd__nand2_1 _11806_ (.A(net55),
    .B(net32),
    .Y(_07530_));
 sky130_fd_sc_hd__a22oi_4 _11807_ (.A1(net44),
    .A2(net2),
    .B1(net3),
    .B2(net33),
    .Y(_07541_));
 sky130_fd_sc_hd__a22o_1 _11808_ (.A1(net44),
    .A2(net2),
    .B1(net3),
    .B2(net33),
    .X(_07552_));
 sky130_fd_sc_hd__and4_1 _11809_ (.A(net33),
    .B(net44),
    .C(net2),
    .D(net3),
    .X(_07563_));
 sky130_fd_sc_hd__nand4_4 _11810_ (.A(net33),
    .B(net44),
    .C(net2),
    .D(net3),
    .Y(_07574_));
 sky130_fd_sc_hd__o211ai_2 _11811_ (.A1(_01780_),
    .A2(_01912_),
    .B1(_07552_),
    .C1(_07574_),
    .Y(_07585_));
 sky130_fd_sc_hd__o21bai_1 _11812_ (.A1(_07541_),
    .A2(_07563_),
    .B1_N(_07530_),
    .Y(_07596_));
 sky130_fd_sc_hd__o22a_2 _11813_ (.A1(_01780_),
    .A2(_01912_),
    .B1(_07541_),
    .B2(_07563_),
    .X(_07607_));
 sky130_fd_sc_hd__o21ai_1 _11814_ (.A1(_07541_),
    .A2(_07563_),
    .B1(_07530_),
    .Y(_07618_));
 sky130_fd_sc_hd__nand4_2 _11815_ (.A(_07552_),
    .B(_07574_),
    .C(net55),
    .D(net32),
    .Y(_07629_));
 sky130_fd_sc_hd__a21oi_1 _11816_ (.A1(_07618_),
    .A2(_07629_),
    .B1(_07508_),
    .Y(_07640_));
 sky130_fd_sc_hd__nand3_4 _11817_ (.A(_07519_),
    .B(_07585_),
    .C(_07596_),
    .Y(_07651_));
 sky130_fd_sc_hd__nand2_2 _11818_ (.A(_07508_),
    .B(_07629_),
    .Y(_07661_));
 sky130_fd_sc_hd__nand3_2 _11819_ (.A(_07618_),
    .B(_07629_),
    .C(_07508_),
    .Y(_07672_));
 sky130_fd_sc_hd__and4_1 _11820_ (.A(net58),
    .B(net59),
    .C(net30),
    .D(net31),
    .X(_07683_));
 sky130_fd_sc_hd__nand4_2 _11821_ (.A(net58),
    .B(net59),
    .C(net30),
    .D(net31),
    .Y(_07694_));
 sky130_fd_sc_hd__a22oi_2 _11822_ (.A1(net59),
    .A2(net30),
    .B1(net31),
    .B2(net58),
    .Y(_07705_));
 sky130_fd_sc_hd__a22o_1 _11823_ (.A1(net59),
    .A2(net30),
    .B1(net31),
    .B2(net58),
    .X(_07716_));
 sky130_fd_sc_hd__o211a_1 _11824_ (.A1(_01835_),
    .A2(_01857_),
    .B1(_07694_),
    .C1(_07716_),
    .X(_07727_));
 sky130_fd_sc_hd__o211a_1 _11825_ (.A1(_07683_),
    .A2(_07705_),
    .B1(net60),
    .C1(net29),
    .X(_07738_));
 sky130_fd_sc_hd__o22a_1 _11826_ (.A1(_01835_),
    .A2(_01857_),
    .B1(_07683_),
    .B2(_07705_),
    .X(_07749_));
 sky130_fd_sc_hd__a22o_1 _11827_ (.A1(net60),
    .A2(net29),
    .B1(_07694_),
    .B2(_07716_),
    .X(_07760_));
 sky130_fd_sc_hd__and4_1 _11828_ (.A(_07716_),
    .B(net29),
    .C(net60),
    .D(_07694_),
    .X(_07771_));
 sky130_fd_sc_hd__nand4_1 _11829_ (.A(_07716_),
    .B(net29),
    .C(net60),
    .D(_07694_),
    .Y(_07782_));
 sky130_fd_sc_hd__nand2_1 _11830_ (.A(_07760_),
    .B(_07782_),
    .Y(_07793_));
 sky130_fd_sc_hd__o2bb2ai_2 _11831_ (.A1_N(_07651_),
    .A2_N(_07672_),
    .B1(_07727_),
    .B2(_07738_),
    .Y(_07804_));
 sky130_fd_sc_hd__o221ai_4 _11832_ (.A1(_07749_),
    .A2(_07771_),
    .B1(_07607_),
    .B2(_07661_),
    .C1(_07651_),
    .Y(_07815_));
 sky130_fd_sc_hd__o2bb2ai_1 _11833_ (.A1_N(_07651_),
    .A2_N(_07672_),
    .B1(_07749_),
    .B2(_07771_),
    .Y(_07826_));
 sky130_fd_sc_hd__nand4_2 _11834_ (.A(_07651_),
    .B(_07672_),
    .C(_07760_),
    .D(_07782_),
    .Y(_07837_));
 sky130_fd_sc_hd__a21boi_2 _11835_ (.A1(_06653_),
    .A2(_06840_),
    .B1_N(_06675_),
    .Y(_07848_));
 sky130_fd_sc_hd__o22ai_2 _11836_ (.A1(_06609_),
    .A2(_06664_),
    .B1(_06829_),
    .B2(_06642_),
    .Y(_07859_));
 sky130_fd_sc_hd__and3_1 _11837_ (.A(_07804_),
    .B(_07848_),
    .C(_07815_),
    .X(_07870_));
 sky130_fd_sc_hd__nand3_2 _11838_ (.A(_07804_),
    .B(_07848_),
    .C(_07815_),
    .Y(_07881_));
 sky130_fd_sc_hd__nand3_4 _11839_ (.A(_07826_),
    .B(_07837_),
    .C(_07859_),
    .Y(_07892_));
 sky130_fd_sc_hd__a31o_2 _11840_ (.A1(_06324_),
    .A2(net63),
    .A3(net23),
    .B1(_06302_),
    .X(_07903_));
 sky130_fd_sc_hd__a31o_1 _11841_ (.A1(_06708_),
    .A2(net60),
    .A3(net28),
    .B1(_06719_),
    .X(_07914_));
 sky130_fd_sc_hd__o21a_1 _11842_ (.A1(_06686_),
    .A2(_06697_),
    .B1(_06730_),
    .X(_07925_));
 sky130_fd_sc_hd__nand2_2 _11843_ (.A(net28),
    .B(net62),
    .Y(_07936_));
 sky130_fd_sc_hd__and4_1 _11844_ (.A(net28),
    .B(net27),
    .C(net61),
    .D(net62),
    .X(_07947_));
 sky130_fd_sc_hd__nand2_2 _11845_ (.A(net28),
    .B(net61),
    .Y(_07958_));
 sky130_fd_sc_hd__a22o_1 _11846_ (.A1(net28),
    .A2(net61),
    .B1(net62),
    .B2(net27),
    .X(_07969_));
 sky130_fd_sc_hd__o2bb2ai_1 _11847_ (.A1_N(_06291_),
    .A2_N(_07958_),
    .B1(_07936_),
    .B2(_06313_),
    .Y(_07980_));
 sky130_fd_sc_hd__o221ai_2 _11848_ (.A1(_01791_),
    .A2(_01890_),
    .B1(_06313_),
    .B2(_07936_),
    .C1(_07969_),
    .Y(_07991_));
 sky130_fd_sc_hd__nand3_1 _11849_ (.A(_07980_),
    .B(net63),
    .C(net26),
    .Y(_08001_));
 sky130_fd_sc_hd__o2111ai_4 _11850_ (.A1(_06313_),
    .A2(_07936_),
    .B1(net26),
    .C1(net63),
    .D1(_07969_),
    .Y(_08012_));
 sky130_fd_sc_hd__o21ai_2 _11851_ (.A1(_01791_),
    .A2(_01890_),
    .B1(_07980_),
    .Y(_08023_));
 sky130_fd_sc_hd__and3_1 _11852_ (.A(_07914_),
    .B(_08012_),
    .C(_08023_),
    .X(_08034_));
 sky130_fd_sc_hd__nand3_1 _11853_ (.A(_07914_),
    .B(_08012_),
    .C(_08023_),
    .Y(_08045_));
 sky130_fd_sc_hd__nand3_2 _11854_ (.A(_07925_),
    .B(_07991_),
    .C(_08001_),
    .Y(_08056_));
 sky130_fd_sc_hd__nand2_1 _11855_ (.A(_08056_),
    .B(_07903_),
    .Y(_08067_));
 sky130_fd_sc_hd__and3_1 _11856_ (.A(_08045_),
    .B(_08056_),
    .C(_07903_),
    .X(_08078_));
 sky130_fd_sc_hd__a21oi_1 _11857_ (.A1(_08045_),
    .A2(_08056_),
    .B1(_07903_),
    .Y(_08089_));
 sky130_fd_sc_hd__a21o_1 _11858_ (.A1(_08045_),
    .A2(_08056_),
    .B1(_07903_),
    .X(_08100_));
 sky130_fd_sc_hd__o21ai_2 _11859_ (.A1(_08034_),
    .A2(_08067_),
    .B1(_08100_),
    .Y(_08111_));
 sky130_fd_sc_hd__a21o_1 _11860_ (.A1(_07881_),
    .A2(_07892_),
    .B1(_08111_),
    .X(_08122_));
 sky130_fd_sc_hd__o211ai_2 _11861_ (.A1(_08078_),
    .A2(_08089_),
    .B1(_07881_),
    .C1(_07892_),
    .Y(_08133_));
 sky130_fd_sc_hd__o2bb2ai_1 _11862_ (.A1_N(_07881_),
    .A2_N(_07892_),
    .B1(_08078_),
    .B2(_08089_),
    .Y(_08144_));
 sky130_fd_sc_hd__o2111ai_1 _11863_ (.A1(_08034_),
    .A2(_08067_),
    .B1(_08100_),
    .C1(_07892_),
    .D1(_07881_),
    .Y(_08155_));
 sky130_fd_sc_hd__a2bb2oi_2 _11864_ (.A1_N(_06851_),
    .A2_N(_06939_),
    .B1(_06928_),
    .B2(_06478_),
    .Y(_08166_));
 sky130_fd_sc_hd__o2bb2ai_1 _11865_ (.A1_N(_06478_),
    .A2_N(_06928_),
    .B1(_06939_),
    .B2(_06851_),
    .Y(_08177_));
 sky130_fd_sc_hd__nand3_4 _11866_ (.A(_08122_),
    .B(_08166_),
    .C(_08133_),
    .Y(_08188_));
 sky130_fd_sc_hd__a21oi_1 _11867_ (.A1(_08122_),
    .A2(_08133_),
    .B1(_08166_),
    .Y(_08199_));
 sky130_fd_sc_hd__nand3_2 _11868_ (.A(_08144_),
    .B(_08155_),
    .C(_08177_),
    .Y(_08210_));
 sky130_fd_sc_hd__nand2_1 _11869_ (.A(_06401_),
    .B(_06467_),
    .Y(_08221_));
 sky130_fd_sc_hd__inv_2 _11870_ (.A(_08221_),
    .Y(_08232_));
 sky130_fd_sc_hd__nand2_1 _11871_ (.A(net1),
    .B(net35),
    .Y(_08243_));
 sky130_fd_sc_hd__nand4_2 _11872_ (.A(net23),
    .B(net12),
    .C(net64),
    .D(net34),
    .Y(_08254_));
 sky130_fd_sc_hd__a22oi_1 _11873_ (.A1(net23),
    .A2(net64),
    .B1(net34),
    .B2(net12),
    .Y(_08265_));
 sky130_fd_sc_hd__a22o_1 _11874_ (.A1(net23),
    .A2(net64),
    .B1(net34),
    .B2(net12),
    .X(_08276_));
 sky130_fd_sc_hd__a22o_1 _11875_ (.A1(net1),
    .A2(net35),
    .B1(_08254_),
    .B2(_08276_),
    .X(_08287_));
 sky130_fd_sc_hd__nand4_2 _11876_ (.A(_08276_),
    .B(net35),
    .C(net1),
    .D(_08254_),
    .Y(_08298_));
 sky130_fd_sc_hd__nand2_1 _11877_ (.A(_08287_),
    .B(_08298_),
    .Y(_08309_));
 sky130_fd_sc_hd__a21o_1 _11878_ (.A1(_08287_),
    .A2(_08298_),
    .B1(_07059_),
    .X(_08320_));
 sky130_fd_sc_hd__nand3_2 _11879_ (.A(_08287_),
    .B(_08298_),
    .C(_07059_),
    .Y(_08330_));
 sky130_fd_sc_hd__nand2_1 _11880_ (.A(_08320_),
    .B(_08330_),
    .Y(_08341_));
 sky130_fd_sc_hd__and3_2 _11881_ (.A(_08221_),
    .B(_08320_),
    .C(_08330_),
    .X(_08352_));
 sky130_fd_sc_hd__and3_1 _11882_ (.A(_06401_),
    .B(_06467_),
    .C(_08341_),
    .X(_08363_));
 sky130_fd_sc_hd__a21oi_1 _11883_ (.A1(_08320_),
    .A2(_08330_),
    .B1(_08232_),
    .Y(_08374_));
 sky130_fd_sc_hd__and3_1 _11884_ (.A(_08232_),
    .B(_08320_),
    .C(_08330_),
    .X(_08385_));
 sky130_fd_sc_hd__nor2_1 _11885_ (.A(_08352_),
    .B(_08363_),
    .Y(_08396_));
 sky130_fd_sc_hd__o2bb2ai_2 _11886_ (.A1_N(_08188_),
    .A2_N(_08210_),
    .B1(_08374_),
    .B2(_08385_),
    .Y(_08407_));
 sky130_fd_sc_hd__o211ai_4 _11887_ (.A1(_08352_),
    .A2(_08363_),
    .B1(_08188_),
    .C1(_08210_),
    .Y(_08418_));
 sky130_fd_sc_hd__o2bb2ai_1 _11888_ (.A1_N(_08188_),
    .A2_N(_08210_),
    .B1(_08352_),
    .B2(_08363_),
    .Y(_08429_));
 sky130_fd_sc_hd__o21ai_1 _11889_ (.A1(_08374_),
    .A2(_08385_),
    .B1(_08188_),
    .Y(_08440_));
 sky130_fd_sc_hd__a22oi_2 _11890_ (.A1(_07015_),
    .A2(_07191_),
    .B1(_08407_),
    .B2(_08418_),
    .Y(_08451_));
 sky130_fd_sc_hd__o211ai_2 _11891_ (.A1(_08199_),
    .A2(_08440_),
    .B1(_08429_),
    .C1(_07497_),
    .Y(_08462_));
 sky130_fd_sc_hd__o2111ai_4 _11892_ (.A1(_07147_),
    .A2(_07026_),
    .B1(_07015_),
    .C1(_08418_),
    .D1(_08407_),
    .Y(_08473_));
 sky130_fd_sc_hd__inv_2 _11893_ (.A(_08473_),
    .Y(_08484_));
 sky130_fd_sc_hd__a21oi_1 _11894_ (.A1(_08462_),
    .A2(_08473_),
    .B1(_07103_),
    .Y(_08495_));
 sky130_fd_sc_hd__a22o_1 _11895_ (.A1(_07081_),
    .A2(_07092_),
    .B1(_08462_),
    .B2(_08473_),
    .X(_08506_));
 sky130_fd_sc_hd__nand2_1 _11896_ (.A(_08473_),
    .B(_07103_),
    .Y(_08517_));
 sky130_fd_sc_hd__o2111a_1 _11897_ (.A1(_05436_),
    .A2(_05480_),
    .B1(_08473_),
    .C1(_07081_),
    .D1(_08462_),
    .X(_08528_));
 sky130_fd_sc_hd__o2bb2ai_4 _11898_ (.A1_N(_07235_),
    .A2_N(_07486_),
    .B1(_08495_),
    .B2(_08528_),
    .Y(_08539_));
 sky130_fd_sc_hd__o221a_1 _11899_ (.A1(_07213_),
    .A2(_07246_),
    .B1(_08451_),
    .B2(_08517_),
    .C1(_08506_),
    .X(_08550_));
 sky130_fd_sc_hd__o221ai_1 _11900_ (.A1(_08451_),
    .A2(_08517_),
    .B1(_07213_),
    .B2(_07246_),
    .C1(_08506_),
    .Y(_08561_));
 sky130_fd_sc_hd__nand2_1 _11901_ (.A(_08539_),
    .B(_08561_),
    .Y(_08572_));
 sky130_fd_sc_hd__a31o_1 _11902_ (.A1(_06072_),
    .A2(_07290_),
    .A3(_07301_),
    .B1(_06127_),
    .X(_08583_));
 sky130_fd_sc_hd__o21ai_2 _11903_ (.A1(_06127_),
    .A2(_07334_),
    .B1(_07323_),
    .Y(_08594_));
 sky130_fd_sc_hd__and3_1 _11904_ (.A(_07344_),
    .B(_08539_),
    .C(_06116_),
    .X(_08605_));
 sky130_fd_sc_hd__nand2_1 _11905_ (.A(_07312_),
    .B(_08539_),
    .Y(_08616_));
 sky130_fd_sc_hd__o211ai_1 _11906_ (.A1(_07334_),
    .A2(_06127_),
    .B1(_07323_),
    .C1(_08572_),
    .Y(_08627_));
 sky130_fd_sc_hd__o211ai_2 _11907_ (.A1(_08572_),
    .A2(_08583_),
    .B1(_08616_),
    .C1(_08627_),
    .Y(_08637_));
 sky130_fd_sc_hd__o31a_1 _11908_ (.A1(_05108_),
    .A2(_06149_),
    .A3(_07355_),
    .B1(_08637_),
    .X(_08648_));
 sky130_fd_sc_hd__nand2_1 _11909_ (.A(_07475_),
    .B(_08637_),
    .Y(_08659_));
 sky130_fd_sc_hd__or4_1 _11910_ (.A(_05108_),
    .B(_06149_),
    .C(_07355_),
    .D(_08637_),
    .X(_08670_));
 sky130_fd_sc_hd__o21a_1 _11911_ (.A1(_05152_),
    .A2(_06215_),
    .B1(_07410_),
    .X(_08681_));
 sky130_fd_sc_hd__o2bb2ai_1 _11912_ (.A1_N(_08659_),
    .A2_N(_08670_),
    .B1(_08681_),
    .B2(_07421_),
    .Y(_08692_));
 sky130_fd_sc_hd__o31a_1 _11913_ (.A1(_07421_),
    .A2(_08648_),
    .A3(_08681_),
    .B1(_08692_),
    .X(net67));
 sky130_fd_sc_hd__o211ai_2 _11914_ (.A1(_07475_),
    .A2(_08637_),
    .B1(_07410_),
    .C1(_07454_),
    .Y(_08713_));
 sky130_fd_sc_hd__o31ai_1 _11915_ (.A1(_07421_),
    .A2(_08648_),
    .A3(_08681_),
    .B1(_08670_),
    .Y(_08724_));
 sky130_fd_sc_hd__o21a_1 _11916_ (.A1(_08078_),
    .A2(_08089_),
    .B1(_07892_),
    .X(_08735_));
 sky130_fd_sc_hd__a32oi_4 _11917_ (.A1(_07804_),
    .A2(_07848_),
    .A3(_07815_),
    .B1(_08111_),
    .B2(_07892_),
    .Y(_08746_));
 sky130_fd_sc_hd__a31o_1 _11918_ (.A1(_07716_),
    .A2(net29),
    .A3(net60),
    .B1(_07683_),
    .X(_08757_));
 sky130_fd_sc_hd__o31a_1 _11919_ (.A1(_01835_),
    .A2(_01857_),
    .A3(_07705_),
    .B1(_07694_),
    .X(_08768_));
 sky130_fd_sc_hd__nor2_1 _11920_ (.A(_01769_),
    .B(_01890_),
    .Y(_08779_));
 sky130_fd_sc_hd__nand2_2 _11921_ (.A(net29),
    .B(net62),
    .Y(_08790_));
 sky130_fd_sc_hd__and4_1 _11922_ (.A(net28),
    .B(net29),
    .C(net61),
    .D(net62),
    .X(_08801_));
 sky130_fd_sc_hd__nand4_1 _11923_ (.A(net28),
    .B(net29),
    .C(net61),
    .D(net62),
    .Y(_08812_));
 sky130_fd_sc_hd__nand2_1 _11924_ (.A(net29),
    .B(net61),
    .Y(_08823_));
 sky130_fd_sc_hd__a22oi_4 _11925_ (.A1(net29),
    .A2(net61),
    .B1(net62),
    .B2(net28),
    .Y(_08834_));
 sky130_fd_sc_hd__a22o_1 _11926_ (.A1(net29),
    .A2(net61),
    .B1(net62),
    .B2(net28),
    .X(_08845_));
 sky130_fd_sc_hd__o221ai_4 _11927_ (.A1(_01769_),
    .A2(_01890_),
    .B1(_07958_),
    .B2(_08790_),
    .C1(_08845_),
    .Y(_08856_));
 sky130_fd_sc_hd__o21ai_1 _11928_ (.A1(_08801_),
    .A2(_08834_),
    .B1(_08779_),
    .Y(_08867_));
 sky130_fd_sc_hd__and4_1 _11929_ (.A(_08845_),
    .B(net63),
    .C(net27),
    .D(_08812_),
    .X(_08878_));
 sky130_fd_sc_hd__o2111ai_1 _11930_ (.A1(_07958_),
    .A2(_08790_),
    .B1(net27),
    .C1(net63),
    .D1(_08845_),
    .Y(_08889_));
 sky130_fd_sc_hd__a22o_1 _11931_ (.A1(net27),
    .A2(net63),
    .B1(_08812_),
    .B2(_08845_),
    .X(_08900_));
 sky130_fd_sc_hd__nand2_1 _11932_ (.A(_08757_),
    .B(_08900_),
    .Y(_08911_));
 sky130_fd_sc_hd__nand3_2 _11933_ (.A(_08900_),
    .B(_08757_),
    .C(_08889_),
    .Y(_08922_));
 sky130_fd_sc_hd__nand3_4 _11934_ (.A(_08768_),
    .B(_08856_),
    .C(_08867_),
    .Y(_08933_));
 sky130_fd_sc_hd__a31o_2 _11935_ (.A1(_07969_),
    .A2(net63),
    .A3(net26),
    .B1(_07947_),
    .X(_08943_));
 sky130_fd_sc_hd__a21oi_2 _11936_ (.A1(_08922_),
    .A2(_08933_),
    .B1(_08943_),
    .Y(_08954_));
 sky130_fd_sc_hd__a21o_1 _11937_ (.A1(_08922_),
    .A2(_08933_),
    .B1(_08943_),
    .X(_08965_));
 sky130_fd_sc_hd__and3_1 _11938_ (.A(_08922_),
    .B(_08933_),
    .C(_08943_),
    .X(_08976_));
 sky130_fd_sc_hd__o211ai_4 _11939_ (.A1(_08878_),
    .A2(_08911_),
    .B1(_08933_),
    .C1(_08943_),
    .Y(_08987_));
 sky130_fd_sc_hd__nand2_2 _11940_ (.A(_08965_),
    .B(_08987_),
    .Y(_08998_));
 sky130_fd_sc_hd__o21ai_2 _11941_ (.A1(_07530_),
    .A2(_07541_),
    .B1(_07574_),
    .Y(_09009_));
 sky130_fd_sc_hd__o21a_1 _11942_ (.A1(_07530_),
    .A2(_07541_),
    .B1(_07574_),
    .X(_09020_));
 sky130_fd_sc_hd__nand2_1 _11943_ (.A(net55),
    .B(net2),
    .Y(_09031_));
 sky130_fd_sc_hd__a22oi_4 _11944_ (.A1(net44),
    .A2(net3),
    .B1(net4),
    .B2(net33),
    .Y(_09042_));
 sky130_fd_sc_hd__a22o_1 _11945_ (.A1(net44),
    .A2(net3),
    .B1(net4),
    .B2(net33),
    .X(_09053_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(net44),
    .B(net4),
    .Y(_09064_));
 sky130_fd_sc_hd__and4_2 _11947_ (.A(net33),
    .B(net44),
    .C(net3),
    .D(net4),
    .X(_09075_));
 sky130_fd_sc_hd__nand4_2 _11948_ (.A(net33),
    .B(net44),
    .C(net3),
    .D(net4),
    .Y(_09086_));
 sky130_fd_sc_hd__o211ai_4 _11949_ (.A1(_01780_),
    .A2(_01901_),
    .B1(_09053_),
    .C1(_09086_),
    .Y(_09097_));
 sky130_fd_sc_hd__o21bai_4 _11950_ (.A1(_09042_),
    .A2(_09075_),
    .B1_N(_09031_),
    .Y(_09108_));
 sky130_fd_sc_hd__a22o_1 _11951_ (.A1(net55),
    .A2(net2),
    .B1(_09053_),
    .B2(_09086_),
    .X(_09119_));
 sky130_fd_sc_hd__a41o_1 _11952_ (.A1(net33),
    .A2(net44),
    .A3(net3),
    .A4(net4),
    .B1(_09031_),
    .X(_09130_));
 sky130_fd_sc_hd__nand3_4 _11953_ (.A(_09020_),
    .B(_09097_),
    .C(_09108_),
    .Y(_09141_));
 sky130_fd_sc_hd__o211a_2 _11954_ (.A1(_09042_),
    .A2(_09130_),
    .B1(_09009_),
    .C1(_09119_),
    .X(_09152_));
 sky130_fd_sc_hd__o211ai_4 _11955_ (.A1(_09042_),
    .A2(_09130_),
    .B1(_09009_),
    .C1(_09119_),
    .Y(_09163_));
 sky130_fd_sc_hd__nand2_1 _11956_ (.A(net60),
    .B(net30),
    .Y(_09174_));
 sky130_fd_sc_hd__a22oi_2 _11957_ (.A1(net59),
    .A2(net31),
    .B1(net32),
    .B2(net58),
    .Y(_09185_));
 sky130_fd_sc_hd__a22o_2 _11958_ (.A1(net59),
    .A2(net31),
    .B1(net32),
    .B2(net58),
    .X(_09196_));
 sky130_fd_sc_hd__and4_1 _11959_ (.A(net58),
    .B(net59),
    .C(net31),
    .D(net32),
    .X(_09207_));
 sky130_fd_sc_hd__nand4_2 _11960_ (.A(net58),
    .B(net59),
    .C(net31),
    .D(net32),
    .Y(_09218_));
 sky130_fd_sc_hd__and3_1 _11961_ (.A(_09174_),
    .B(_09196_),
    .C(_09218_),
    .X(_09229_));
 sky130_fd_sc_hd__o211ai_2 _11962_ (.A1(_01835_),
    .A2(_01868_),
    .B1(_09196_),
    .C1(_09218_),
    .Y(_09240_));
 sky130_fd_sc_hd__o211a_1 _11963_ (.A1(_09185_),
    .A2(_09207_),
    .B1(net60),
    .C1(net30),
    .X(_09250_));
 sky130_fd_sc_hd__a21o_1 _11964_ (.A1(_09196_),
    .A2(_09218_),
    .B1(_09174_),
    .X(_09261_));
 sky130_fd_sc_hd__o22a_1 _11965_ (.A1(_01835_),
    .A2(_01868_),
    .B1(_09185_),
    .B2(_09207_),
    .X(_09272_));
 sky130_fd_sc_hd__and4_1 _11966_ (.A(_09196_),
    .B(_09218_),
    .C(net60),
    .D(net30),
    .X(_09283_));
 sky130_fd_sc_hd__nand2_1 _11967_ (.A(_09240_),
    .B(_09261_),
    .Y(_09294_));
 sky130_fd_sc_hd__o2bb2ai_4 _11968_ (.A1_N(_09141_),
    .A2_N(_09163_),
    .B1(_09272_),
    .B2(_09283_),
    .Y(_09305_));
 sky130_fd_sc_hd__a32oi_4 _11969_ (.A1(_09020_),
    .A2(_09097_),
    .A3(_09108_),
    .B1(_09240_),
    .B2(_09261_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21ai_2 _11970_ (.A1(_09229_),
    .A2(_09250_),
    .B1(_09141_),
    .Y(_09327_));
 sky130_fd_sc_hd__o211ai_4 _11971_ (.A1(_09229_),
    .A2(_09250_),
    .B1(_09141_),
    .C1(_09163_),
    .Y(_09338_));
 sky130_fd_sc_hd__inv_2 _11972_ (.A(_09338_),
    .Y(_09349_));
 sky130_fd_sc_hd__o22ai_4 _11973_ (.A1(_07607_),
    .A2(_07661_),
    .B1(_07793_),
    .B2(_07640_),
    .Y(_09360_));
 sky130_fd_sc_hd__a21oi_4 _11974_ (.A1(_09305_),
    .A2(_09338_),
    .B1(_09360_),
    .Y(_09371_));
 sky130_fd_sc_hd__a21o_1 _11975_ (.A1(_09305_),
    .A2(_09338_),
    .B1(_09360_),
    .X(_09382_));
 sky130_fd_sc_hd__nand2_2 _11976_ (.A(_09305_),
    .B(_09360_),
    .Y(_09393_));
 sky130_fd_sc_hd__o211a_1 _11977_ (.A1(_09152_),
    .A2(_09327_),
    .B1(_09360_),
    .C1(_09305_),
    .X(_09404_));
 sky130_fd_sc_hd__o211ai_4 _11978_ (.A1(_09152_),
    .A2(_09327_),
    .B1(_09360_),
    .C1(_09305_),
    .Y(_09415_));
 sky130_fd_sc_hd__nand3_2 _11979_ (.A(_08965_),
    .B(_08987_),
    .C(_09415_),
    .Y(_09426_));
 sky130_fd_sc_hd__o22ai_2 _11980_ (.A1(_08954_),
    .A2(_08976_),
    .B1(_09371_),
    .B2(_09404_),
    .Y(_09437_));
 sky130_fd_sc_hd__o221ai_4 _11981_ (.A1(_08954_),
    .A2(_08976_),
    .B1(_09349_),
    .B2(_09393_),
    .C1(_09382_),
    .Y(_09448_));
 sky130_fd_sc_hd__o21bai_2 _11982_ (.A1(_09371_),
    .A2(_09404_),
    .B1_N(_08998_),
    .Y(_09459_));
 sky130_fd_sc_hd__o211a_1 _11983_ (.A1(_09371_),
    .A2(_09426_),
    .B1(_08746_),
    .C1(_09437_),
    .X(_09470_));
 sky130_fd_sc_hd__o211ai_4 _11984_ (.A1(_09371_),
    .A2(_09426_),
    .B1(_08746_),
    .C1(_09437_),
    .Y(_09481_));
 sky130_fd_sc_hd__o211ai_4 _11985_ (.A1(_07870_),
    .A2(_08735_),
    .B1(_09448_),
    .C1(_09459_),
    .Y(_09492_));
 sky130_fd_sc_hd__and4_1 _11986_ (.A(net26),
    .B(net23),
    .C(net64),
    .D(net34),
    .X(_09503_));
 sky130_fd_sc_hd__nand4_1 _11987_ (.A(net26),
    .B(net23),
    .C(net64),
    .D(net34),
    .Y(_09514_));
 sky130_fd_sc_hd__a22o_1 _11988_ (.A1(net26),
    .A2(net64),
    .B1(net34),
    .B2(net23),
    .X(_09525_));
 sky130_fd_sc_hd__o2bb2ai_1 _11989_ (.A1_N(_09514_),
    .A2_N(_09525_),
    .B1(_01824_),
    .B2(_01934_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand4_2 _11990_ (.A(_09525_),
    .B(net35),
    .C(net12),
    .D(_09514_),
    .Y(_09546_));
 sky130_fd_sc_hd__o21ai_1 _11991_ (.A1(_08243_),
    .A2(_08265_),
    .B1(_08254_),
    .Y(_09557_));
 sky130_fd_sc_hd__a21oi_1 _11992_ (.A1(_09535_),
    .A2(_09546_),
    .B1(_09557_),
    .Y(_09568_));
 sky130_fd_sc_hd__a21o_1 _11993_ (.A1(_09535_),
    .A2(_09546_),
    .B1(_09557_),
    .X(_09579_));
 sky130_fd_sc_hd__and3_1 _11994_ (.A(_09535_),
    .B(_09546_),
    .C(_09557_),
    .X(_09590_));
 sky130_fd_sc_hd__nand3_1 _11995_ (.A(_09535_),
    .B(_09546_),
    .C(_09557_),
    .Y(_09601_));
 sky130_fd_sc_hd__nand2_1 _11996_ (.A(net1),
    .B(net36),
    .Y(_09612_));
 sky130_fd_sc_hd__o21ai_1 _11997_ (.A1(_09568_),
    .A2(_09590_),
    .B1(_09612_),
    .Y(_09623_));
 sky130_fd_sc_hd__nand4_1 _11998_ (.A(_09579_),
    .B(_09601_),
    .C(net1),
    .D(net36),
    .Y(_09634_));
 sky130_fd_sc_hd__o21bai_1 _11999_ (.A1(_09568_),
    .A2(_09590_),
    .B1_N(_09612_),
    .Y(_09645_));
 sky130_fd_sc_hd__nand3_1 _12000_ (.A(_09579_),
    .B(_09601_),
    .C(_09612_),
    .Y(_09656_));
 sky130_fd_sc_hd__a32oi_4 _12001_ (.A1(_07914_),
    .A2(_08012_),
    .A3(_08023_),
    .B1(_08056_),
    .B2(_07903_),
    .Y(_09667_));
 sky130_fd_sc_hd__a32o_1 _12002_ (.A1(_07914_),
    .A2(_08012_),
    .A3(_08023_),
    .B1(_08056_),
    .B2(_07903_),
    .X(_09678_));
 sky130_fd_sc_hd__nand3_2 _12003_ (.A(_09645_),
    .B(_09656_),
    .C(_09667_),
    .Y(_09689_));
 sky130_fd_sc_hd__inv_2 _12004_ (.A(_09689_),
    .Y(_09700_));
 sky130_fd_sc_hd__nand3_2 _12005_ (.A(_09623_),
    .B(_09634_),
    .C(_09678_),
    .Y(_09711_));
 sky130_fd_sc_hd__inv_2 _12006_ (.A(_09711_),
    .Y(_09722_));
 sky130_fd_sc_hd__o2bb2a_1 _12007_ (.A1_N(_09689_),
    .A2_N(_09711_),
    .B1(_07070_),
    .B2(_08309_),
    .X(_09733_));
 sky130_fd_sc_hd__a2bb2o_1 _12008_ (.A1_N(_07070_),
    .A2_N(_08309_),
    .B1(_09689_),
    .B2(_09711_),
    .X(_09744_));
 sky130_fd_sc_hd__and4_1 _12009_ (.A(_08287_),
    .B(_08298_),
    .C(_09689_),
    .D(_07059_),
    .X(_09755_));
 sky130_fd_sc_hd__and4b_1 _12010_ (.A_N(_08309_),
    .B(_09689_),
    .C(_09711_),
    .D(_07059_),
    .X(_09766_));
 sky130_fd_sc_hd__nand3b_1 _12011_ (.A_N(_08330_),
    .B(_09689_),
    .C(_09711_),
    .Y(_09777_));
 sky130_fd_sc_hd__and3_1 _12012_ (.A(_08330_),
    .B(_09689_),
    .C(_09711_),
    .X(_09788_));
 sky130_fd_sc_hd__a21oi_1 _12013_ (.A1(_09689_),
    .A2(_09711_),
    .B1(_08330_),
    .Y(_09799_));
 sky130_fd_sc_hd__nand2_1 _12014_ (.A(_09744_),
    .B(_09777_),
    .Y(_09810_));
 sky130_fd_sc_hd__o2bb2ai_1 _12015_ (.A1_N(_09481_),
    .A2_N(_09492_),
    .B1(_09788_),
    .B2(_09799_),
    .Y(_09821_));
 sky130_fd_sc_hd__o211ai_2 _12016_ (.A1(_09733_),
    .A2(_09766_),
    .B1(_09481_),
    .C1(_09492_),
    .Y(_09832_));
 sky130_fd_sc_hd__o2bb2ai_1 _12017_ (.A1_N(_09481_),
    .A2_N(_09492_),
    .B1(_09733_),
    .B2(_09766_),
    .Y(_09842_));
 sky130_fd_sc_hd__o21a_1 _12018_ (.A1(_09788_),
    .A2(_09799_),
    .B1(_09492_),
    .X(_09853_));
 sky130_fd_sc_hd__o211ai_1 _12019_ (.A1(_09788_),
    .A2(_09799_),
    .B1(_09481_),
    .C1(_09492_),
    .Y(_09864_));
 sky130_fd_sc_hd__a21o_1 _12020_ (.A1(_08188_),
    .A2(_08396_),
    .B1(_08199_),
    .X(_09875_));
 sky130_fd_sc_hd__a21oi_1 _12021_ (.A1(_08188_),
    .A2(_08396_),
    .B1(_08199_),
    .Y(_09886_));
 sky130_fd_sc_hd__nand3_2 _12022_ (.A(_09821_),
    .B(_09832_),
    .C(_09886_),
    .Y(_09897_));
 sky130_fd_sc_hd__and3_1 _12023_ (.A(_09875_),
    .B(_09864_),
    .C(_09842_),
    .X(_09908_));
 sky130_fd_sc_hd__nand3_1 _12024_ (.A(_09875_),
    .B(_09864_),
    .C(_09842_),
    .Y(_09919_));
 sky130_fd_sc_hd__o2bb2ai_2 _12025_ (.A1_N(_09897_),
    .A2_N(_09919_),
    .B1(_08232_),
    .B2(_08341_),
    .Y(_09930_));
 sky130_fd_sc_hd__a311oi_2 _12026_ (.A1(_09821_),
    .A2(_09832_),
    .A3(_09886_),
    .B1(_08341_),
    .C1(_08232_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand3_2 _12027_ (.A(_09919_),
    .B(_08352_),
    .C(_09897_),
    .Y(_09952_));
 sky130_fd_sc_hd__a21oi_1 _12028_ (.A1(_07081_),
    .A2(_07092_),
    .B1(_08451_),
    .Y(_09963_));
 sky130_fd_sc_hd__a31o_1 _12029_ (.A1(_08473_),
    .A2(_07081_),
    .A3(_07092_),
    .B1(_08451_),
    .X(_09974_));
 sky130_fd_sc_hd__o2bb2ai_2 _12030_ (.A1_N(_09930_),
    .A2_N(_09952_),
    .B1(_09963_),
    .B2(_08484_),
    .Y(_09985_));
 sky130_fd_sc_hd__and3_1 _12031_ (.A(_09974_),
    .B(_09952_),
    .C(_09930_),
    .X(_09996_));
 sky130_fd_sc_hd__nand3_2 _12032_ (.A(_09974_),
    .B(_09952_),
    .C(_09930_),
    .Y(_10007_));
 sky130_fd_sc_hd__a21oi_1 _12033_ (.A1(_09985_),
    .A2(_10007_),
    .B1(_08550_),
    .Y(_10018_));
 sky130_fd_sc_hd__a21o_1 _12034_ (.A1(_09985_),
    .A2(_10007_),
    .B1(_08550_),
    .X(_10029_));
 sky130_fd_sc_hd__nand3_2 _12035_ (.A(_08550_),
    .B(_09985_),
    .C(_10007_),
    .Y(_10040_));
 sky130_fd_sc_hd__a22oi_2 _12036_ (.A1(_08539_),
    .A2(_08594_),
    .B1(_10029_),
    .B2(_10040_),
    .Y(_10051_));
 sky130_fd_sc_hd__or2_1 _12037_ (.A(_08616_),
    .B(_10018_),
    .X(_10062_));
 sky130_fd_sc_hd__and3_1 _12038_ (.A(_08605_),
    .B(_10029_),
    .C(_10040_),
    .X(_10073_));
 sky130_fd_sc_hd__a41oi_4 _12039_ (.A1(_08539_),
    .A2(_08594_),
    .A3(_10029_),
    .A4(_10040_),
    .B1(_10051_),
    .Y(_10084_));
 sky130_fd_sc_hd__xor2_1 _12040_ (.A(_08724_),
    .B(_10084_),
    .X(net68));
 sky130_fd_sc_hd__a21oi_1 _12041_ (.A1(_08352_),
    .A2(_09897_),
    .B1(_09908_),
    .Y(_10105_));
 sky130_fd_sc_hd__o21a_1 _12042_ (.A1(_07070_),
    .A2(_08309_),
    .B1(_09711_),
    .X(_10115_));
 sky130_fd_sc_hd__o2bb2ai_1 _12043_ (.A1_N(_08943_),
    .A2_N(_08933_),
    .B1(_08878_),
    .B2(_08911_),
    .Y(_10126_));
 sky130_fd_sc_hd__a31oi_1 _12044_ (.A1(_09525_),
    .A2(net35),
    .A3(net12),
    .B1(_09503_),
    .Y(_10137_));
 sky130_fd_sc_hd__a31o_1 _12045_ (.A1(_09525_),
    .A2(net35),
    .A3(net12),
    .B1(_09503_),
    .X(_10148_));
 sky130_fd_sc_hd__nand2_1 _12046_ (.A(net23),
    .B(net35),
    .Y(_10159_));
 sky130_fd_sc_hd__nand4_4 _12047_ (.A(net27),
    .B(net26),
    .C(net64),
    .D(net34),
    .Y(_10170_));
 sky130_fd_sc_hd__a22oi_1 _12048_ (.A1(net27),
    .A2(net64),
    .B1(net34),
    .B2(net26),
    .Y(_10181_));
 sky130_fd_sc_hd__a22o_2 _12049_ (.A1(net27),
    .A2(net64),
    .B1(net34),
    .B2(net26),
    .X(_10192_));
 sky130_fd_sc_hd__o211ai_1 _12050_ (.A1(_01802_),
    .A2(_01934_),
    .B1(_10170_),
    .C1(_10192_),
    .Y(_10203_));
 sky130_fd_sc_hd__a21o_1 _12051_ (.A1(_10170_),
    .A2(_10192_),
    .B1(_10159_),
    .X(_10214_));
 sky130_fd_sc_hd__a22o_1 _12052_ (.A1(net23),
    .A2(net35),
    .B1(_10170_),
    .B2(_10192_),
    .X(_10225_));
 sky130_fd_sc_hd__nand4_1 _12053_ (.A(_10192_),
    .B(net35),
    .C(net23),
    .D(_10170_),
    .Y(_10236_));
 sky130_fd_sc_hd__and3_1 _12054_ (.A(_10214_),
    .B(_10137_),
    .C(_10203_),
    .X(_10247_));
 sky130_fd_sc_hd__nand3_1 _12055_ (.A(_10214_),
    .B(_10137_),
    .C(_10203_),
    .Y(_10258_));
 sky130_fd_sc_hd__nand3_2 _12056_ (.A(_10148_),
    .B(_10225_),
    .C(_10236_),
    .Y(_10269_));
 sky130_fd_sc_hd__nand2_1 _12057_ (.A(net12),
    .B(net36),
    .Y(_10280_));
 sky130_fd_sc_hd__and4_1 _12058_ (.A(net12),
    .B(net1),
    .C(net36),
    .D(net37),
    .X(_10291_));
 sky130_fd_sc_hd__nand4_2 _12059_ (.A(net12),
    .B(net1),
    .C(net36),
    .D(net37),
    .Y(_10302_));
 sky130_fd_sc_hd__a22oi_2 _12060_ (.A1(net12),
    .A2(net36),
    .B1(net37),
    .B2(net1),
    .Y(_10313_));
 sky130_fd_sc_hd__a21oi_1 _12061_ (.A1(net1),
    .A2(net37),
    .B1(_10280_),
    .Y(_10324_));
 sky130_fd_sc_hd__and3_1 _12062_ (.A(_10280_),
    .B(net37),
    .C(net1),
    .X(_10335_));
 sky130_fd_sc_hd__o2bb2ai_1 _12063_ (.A1_N(_10258_),
    .A2_N(_10269_),
    .B1(_10291_),
    .B2(_10313_),
    .Y(_10346_));
 sky130_fd_sc_hd__o211ai_1 _12064_ (.A1(_10324_),
    .A2(_10335_),
    .B1(_10258_),
    .C1(_10269_),
    .Y(_10357_));
 sky130_fd_sc_hd__o2bb2ai_1 _12065_ (.A1_N(_10258_),
    .A2_N(_10269_),
    .B1(_10324_),
    .B2(_10335_),
    .Y(_10368_));
 sky130_fd_sc_hd__o211ai_1 _12066_ (.A1(_10291_),
    .A2(_10313_),
    .B1(_10258_),
    .C1(_10269_),
    .Y(_10378_));
 sky130_fd_sc_hd__nand4_1 _12067_ (.A(_08922_),
    .B(_08987_),
    .C(_10368_),
    .D(_10378_),
    .Y(_10389_));
 sky130_fd_sc_hd__nand3_2 _12068_ (.A(_10126_),
    .B(_10346_),
    .C(_10357_),
    .Y(_10400_));
 sky130_fd_sc_hd__a31o_1 _12069_ (.A1(_09579_),
    .A2(net36),
    .A3(net1),
    .B1(_09590_),
    .X(_10411_));
 sky130_fd_sc_hd__a21o_1 _12070_ (.A1(_10389_),
    .A2(_10400_),
    .B1(_10411_),
    .X(_10422_));
 sky130_fd_sc_hd__nand3_2 _12071_ (.A(_10389_),
    .B(_10400_),
    .C(_10411_),
    .Y(_10433_));
 sky130_fd_sc_hd__nand2_2 _12072_ (.A(_10422_),
    .B(_10433_),
    .Y(_10444_));
 sky130_fd_sc_hd__o22ai_2 _12073_ (.A1(_09349_),
    .A2(_09393_),
    .B1(_09371_),
    .B2(_08998_),
    .Y(_10455_));
 sky130_fd_sc_hd__o32a_1 _12074_ (.A1(_08954_),
    .A2(_08976_),
    .A3(_09371_),
    .B1(_09393_),
    .B2(_09349_),
    .X(_10466_));
 sky130_fd_sc_hd__nand2_2 _12075_ (.A(net61),
    .B(net30),
    .Y(_10477_));
 sky130_fd_sc_hd__a22oi_2 _12076_ (.A1(net61),
    .A2(net30),
    .B1(net62),
    .B2(net29),
    .Y(_10488_));
 sky130_fd_sc_hd__a22o_1 _12077_ (.A1(net61),
    .A2(net30),
    .B1(net62),
    .B2(net29),
    .X(_10499_));
 sky130_fd_sc_hd__nand2_2 _12078_ (.A(net30),
    .B(net62),
    .Y(_10510_));
 sky130_fd_sc_hd__and4_1 _12079_ (.A(net29),
    .B(net61),
    .C(net30),
    .D(net62),
    .X(_10521_));
 sky130_fd_sc_hd__or2_1 _12080_ (.A(_08790_),
    .B(_10477_),
    .X(_10532_));
 sky130_fd_sc_hd__o2111ai_4 _12081_ (.A1(_08823_),
    .A2(_10510_),
    .B1(net28),
    .C1(net63),
    .D1(_10499_),
    .Y(_10543_));
 sky130_fd_sc_hd__o22ai_4 _12082_ (.A1(_01748_),
    .A2(_01890_),
    .B1(_10488_),
    .B2(_10521_),
    .Y(_10554_));
 sky130_fd_sc_hd__o21a_1 _12083_ (.A1(_01835_),
    .A2(_01868_),
    .B1(_09218_),
    .X(_10565_));
 sky130_fd_sc_hd__o21ai_1 _12084_ (.A1(_01835_),
    .A2(_01868_),
    .B1(_09218_),
    .Y(_10576_));
 sky130_fd_sc_hd__o2bb2ai_2 _12085_ (.A1_N(_10543_),
    .A2_N(_10554_),
    .B1(_10565_),
    .B2(_09185_),
    .Y(_10587_));
 sky130_fd_sc_hd__nand4_4 _12086_ (.A(_09196_),
    .B(_10543_),
    .C(_10554_),
    .D(_10576_),
    .Y(_10598_));
 sky130_fd_sc_hd__o22a_1 _12087_ (.A1(_01769_),
    .A2(_01890_),
    .B1(_07958_),
    .B2(_08790_),
    .X(_10609_));
 sky130_fd_sc_hd__a31o_1 _12088_ (.A1(_08845_),
    .A2(net63),
    .A3(net27),
    .B1(_08801_),
    .X(_10620_));
 sky130_fd_sc_hd__o2bb2ai_4 _12089_ (.A1_N(_10587_),
    .A2_N(_10598_),
    .B1(_10609_),
    .B2(_08834_),
    .Y(_10631_));
 sky130_fd_sc_hd__nand3_2 _12090_ (.A(_10587_),
    .B(_10598_),
    .C(_10620_),
    .Y(_10641_));
 sky130_fd_sc_hd__nand2_1 _12091_ (.A(_10631_),
    .B(_10641_),
    .Y(_10652_));
 sky130_fd_sc_hd__a21oi_2 _12092_ (.A1(_09141_),
    .A2(_09294_),
    .B1(_09152_),
    .Y(_10663_));
 sky130_fd_sc_hd__nor2_1 _12093_ (.A(_09031_),
    .B(_09042_),
    .Y(_10674_));
 sky130_fd_sc_hd__o32a_1 _12094_ (.A1(_01737_),
    .A2(_01923_),
    .A3(_09064_),
    .B1(_09042_),
    .B2(_09031_),
    .X(_10685_));
 sky130_fd_sc_hd__nand2_1 _12095_ (.A(net55),
    .B(net3),
    .Y(_10696_));
 sky130_fd_sc_hd__nand2_1 _12096_ (.A(net33),
    .B(net5),
    .Y(_10707_));
 sky130_fd_sc_hd__and4_2 _12097_ (.A(net33),
    .B(net44),
    .C(net4),
    .D(net5),
    .X(_10718_));
 sky130_fd_sc_hd__nand4_2 _12098_ (.A(net33),
    .B(net44),
    .C(net4),
    .D(net5),
    .Y(_10729_));
 sky130_fd_sc_hd__a22oi_4 _12099_ (.A1(net44),
    .A2(net4),
    .B1(net5),
    .B2(net33),
    .Y(_10740_));
 sky130_fd_sc_hd__a22o_1 _12100_ (.A1(net44),
    .A2(net4),
    .B1(net5),
    .B2(net33),
    .X(_10751_));
 sky130_fd_sc_hd__o211ai_2 _12101_ (.A1(_01780_),
    .A2(_01923_),
    .B1(_10729_),
    .C1(_10751_),
    .Y(_10762_));
 sky130_fd_sc_hd__o21bai_2 _12102_ (.A1(_10718_),
    .A2(_10740_),
    .B1_N(_10696_),
    .Y(_10773_));
 sky130_fd_sc_hd__a22o_1 _12103_ (.A1(net55),
    .A2(net3),
    .B1(_10729_),
    .B2(_10751_),
    .X(_10784_));
 sky130_fd_sc_hd__a41o_1 _12104_ (.A1(net33),
    .A2(net44),
    .A3(net4),
    .A4(net5),
    .B1(_10696_),
    .X(_10795_));
 sky130_fd_sc_hd__nand3_4 _12105_ (.A(_10685_),
    .B(_10762_),
    .C(_10773_),
    .Y(_10806_));
 sky130_fd_sc_hd__a2bb2oi_1 _12106_ (.A1_N(_09075_),
    .A2_N(_10674_),
    .B1(_10762_),
    .B2(_10773_),
    .Y(_10817_));
 sky130_fd_sc_hd__o221ai_4 _12107_ (.A1(_09075_),
    .A2(_10674_),
    .B1(_10740_),
    .B2(_10795_),
    .C1(_10784_),
    .Y(_10828_));
 sky130_fd_sc_hd__nand2_1 _12108_ (.A(net60),
    .B(net31),
    .Y(_10839_));
 sky130_fd_sc_hd__a22oi_2 _12109_ (.A1(net58),
    .A2(net2),
    .B1(net32),
    .B2(net59),
    .Y(_10850_));
 sky130_fd_sc_hd__a22o_1 _12110_ (.A1(net58),
    .A2(net2),
    .B1(net32),
    .B2(net59),
    .X(_10861_));
 sky130_fd_sc_hd__and4_1 _12111_ (.A(net58),
    .B(net59),
    .C(net2),
    .D(net32),
    .X(_10872_));
 sky130_fd_sc_hd__nand4_2 _12112_ (.A(net58),
    .B(net59),
    .C(net2),
    .D(net32),
    .Y(_10882_));
 sky130_fd_sc_hd__and3_1 _12113_ (.A(_10839_),
    .B(_10861_),
    .C(_10882_),
    .X(_10893_));
 sky130_fd_sc_hd__o211ai_1 _12114_ (.A1(_01835_),
    .A2(_01879_),
    .B1(_10861_),
    .C1(_10882_),
    .Y(_10904_));
 sky130_fd_sc_hd__o211a_1 _12115_ (.A1(_10850_),
    .A2(_10872_),
    .B1(net60),
    .C1(net31),
    .X(_10915_));
 sky130_fd_sc_hd__a21o_1 _12116_ (.A1(_10861_),
    .A2(_10882_),
    .B1(_10839_),
    .X(_10926_));
 sky130_fd_sc_hd__o22a_1 _12117_ (.A1(_01835_),
    .A2(_01879_),
    .B1(_10850_),
    .B2(_10872_),
    .X(_10937_));
 sky130_fd_sc_hd__and4_1 _12118_ (.A(_10861_),
    .B(_10882_),
    .C(net60),
    .D(net31),
    .X(_10948_));
 sky130_fd_sc_hd__nand2_1 _12119_ (.A(_10904_),
    .B(_10926_),
    .Y(_10959_));
 sky130_fd_sc_hd__o211ai_2 _12120_ (.A1(_10893_),
    .A2(_10915_),
    .B1(_10806_),
    .C1(_10828_),
    .Y(_10970_));
 sky130_fd_sc_hd__o2bb2ai_2 _12121_ (.A1_N(_10806_),
    .A2_N(_10828_),
    .B1(_10937_),
    .B2(_10948_),
    .Y(_10981_));
 sky130_fd_sc_hd__o211ai_4 _12122_ (.A1(_10937_),
    .A2(_10948_),
    .B1(_10806_),
    .C1(_10828_),
    .Y(_10992_));
 sky130_fd_sc_hd__o2bb2ai_2 _12123_ (.A1_N(_10806_),
    .A2_N(_10828_),
    .B1(_10893_),
    .B2(_10915_),
    .Y(_11003_));
 sky130_fd_sc_hd__nand3_4 _12124_ (.A(_11003_),
    .B(_10663_),
    .C(_10992_),
    .Y(_11014_));
 sky130_fd_sc_hd__o211a_2 _12125_ (.A1(_09152_),
    .A2(_09316_),
    .B1(_10970_),
    .C1(_10981_),
    .X(_11025_));
 sky130_fd_sc_hd__o211ai_4 _12126_ (.A1(_09152_),
    .A2(_09316_),
    .B1(_10970_),
    .C1(_10981_),
    .Y(_11036_));
 sky130_fd_sc_hd__nand3_2 _12127_ (.A(_10652_),
    .B(_11014_),
    .C(_11036_),
    .Y(_11047_));
 sky130_fd_sc_hd__a21o_2 _12128_ (.A1(_11014_),
    .A2(_11036_),
    .B1(_10652_),
    .X(_11058_));
 sky130_fd_sc_hd__a22o_1 _12129_ (.A1(_10631_),
    .A2(_10641_),
    .B1(_11014_),
    .B2(_11036_),
    .X(_11069_));
 sky130_fd_sc_hd__a31oi_2 _12130_ (.A1(_10663_),
    .A2(_10992_),
    .A3(_11003_),
    .B1(_10652_),
    .Y(_11080_));
 sky130_fd_sc_hd__nand4_2 _12131_ (.A(_10631_),
    .B(_10641_),
    .C(_11014_),
    .D(_11036_),
    .Y(_11091_));
 sky130_fd_sc_hd__o2111ai_4 _12132_ (.A1(_08998_),
    .A2(_09371_),
    .B1(_09415_),
    .C1(_11047_),
    .D1(_11058_),
    .Y(_11101_));
 sky130_fd_sc_hd__nand3_4 _12133_ (.A(_11069_),
    .B(_11091_),
    .C(_10455_),
    .Y(_11112_));
 sky130_fd_sc_hd__a22o_1 _12134_ (.A1(_10422_),
    .A2(_10433_),
    .B1(_11101_),
    .B2(_11112_),
    .X(_11123_));
 sky130_fd_sc_hd__nand4_1 _12135_ (.A(_10422_),
    .B(_10433_),
    .C(_11101_),
    .D(_11112_),
    .Y(_11134_));
 sky130_fd_sc_hd__nand3_1 _12136_ (.A(_10444_),
    .B(_11101_),
    .C(_11112_),
    .Y(_11145_));
 sky130_fd_sc_hd__a21o_1 _12137_ (.A1(_11101_),
    .A2(_11112_),
    .B1(_10444_),
    .X(_11156_));
 sky130_fd_sc_hd__a31oi_1 _12138_ (.A1(_09492_),
    .A2(_09744_),
    .A3(_09777_),
    .B1(_09470_),
    .Y(_11167_));
 sky130_fd_sc_hd__a21boi_1 _12139_ (.A1(_09481_),
    .A2(_09810_),
    .B1_N(_09492_),
    .Y(_11178_));
 sky130_fd_sc_hd__a2bb2oi_1 _12140_ (.A1_N(_09470_),
    .A2_N(_09853_),
    .B1(_11145_),
    .B2(_11156_),
    .Y(_11189_));
 sky130_fd_sc_hd__nand3_2 _12141_ (.A(_11123_),
    .B(_11134_),
    .C(_11178_),
    .Y(_11200_));
 sky130_fd_sc_hd__a21oi_1 _12142_ (.A1(_11123_),
    .A2(_11134_),
    .B1(_11178_),
    .Y(_11211_));
 sky130_fd_sc_hd__nand3_1 _12143_ (.A(_11145_),
    .B(_11156_),
    .C(_11167_),
    .Y(_11222_));
 sky130_fd_sc_hd__o211a_2 _12144_ (.A1(_09722_),
    .A2(_09755_),
    .B1(_11200_),
    .C1(_11222_),
    .X(_11233_));
 sky130_fd_sc_hd__o211ai_2 _12145_ (.A1(_09722_),
    .A2(_09755_),
    .B1(_11200_),
    .C1(_11222_),
    .Y(_11244_));
 sky130_fd_sc_hd__a2bb2oi_1 _12146_ (.A1_N(_09700_),
    .A2_N(_10115_),
    .B1(_11200_),
    .B2(_11222_),
    .Y(_11255_));
 sky130_fd_sc_hd__o22ai_2 _12147_ (.A1(_09700_),
    .A2(_10115_),
    .B1(_11189_),
    .B2(_11211_),
    .Y(_11266_));
 sky130_fd_sc_hd__o21ai_2 _12148_ (.A1(_09908_),
    .A2(_09941_),
    .B1(_11266_),
    .Y(_00000_));
 sky130_fd_sc_hd__o211ai_1 _12149_ (.A1(_09908_),
    .A2(_09941_),
    .B1(_11244_),
    .C1(_11266_),
    .Y(_00011_));
 sky130_fd_sc_hd__o21ai_2 _12150_ (.A1(_11233_),
    .A2(_11255_),
    .B1(_10105_),
    .Y(_00022_));
 sky130_fd_sc_hd__o211a_1 _12151_ (.A1(_11233_),
    .A2(_00000_),
    .B1(_09996_),
    .C1(_00022_),
    .X(_00032_));
 sky130_fd_sc_hd__o211ai_4 _12152_ (.A1(_11233_),
    .A2(_00000_),
    .B1(_09996_),
    .C1(_00022_),
    .Y(_00043_));
 sky130_fd_sc_hd__a21oi_1 _12153_ (.A1(_00011_),
    .A2(_00022_),
    .B1(_09996_),
    .Y(_00054_));
 sky130_fd_sc_hd__a32o_1 _12154_ (.A1(_09930_),
    .A2(_09974_),
    .A3(_09952_),
    .B1(_00022_),
    .B2(_00011_),
    .X(_00065_));
 sky130_fd_sc_hd__nand2_1 _12155_ (.A(_00043_),
    .B(_00065_),
    .Y(_00076_));
 sky130_fd_sc_hd__o21ai_1 _12156_ (.A1(_08616_),
    .A2(_10018_),
    .B1(_10040_),
    .Y(_00087_));
 sky130_fd_sc_hd__a21o_1 _12157_ (.A1(_00043_),
    .A2(_00065_),
    .B1(_00087_),
    .X(_00098_));
 sky130_fd_sc_hd__o2111ai_1 _12158_ (.A1(_08616_),
    .A2(_10018_),
    .B1(_10040_),
    .C1(_00043_),
    .D1(_00065_),
    .Y(_00109_));
 sky130_fd_sc_hd__o21ai_1 _12159_ (.A1(_00032_),
    .A2(_00054_),
    .B1(_00087_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand4_2 _12160_ (.A(_09985_),
    .B(_10007_),
    .C(_00065_),
    .D(_08550_),
    .Y(_00131_));
 sky130_fd_sc_hd__nand2_1 _12161_ (.A(_00109_),
    .B(_00120_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand4_1 _12162_ (.A(_00142_),
    .B(_08713_),
    .C(_08659_),
    .D(_10084_),
    .Y(_00153_));
 sky130_fd_sc_hd__a31o_1 _12163_ (.A1(_08659_),
    .A2(_08713_),
    .A3(_10084_),
    .B1(_00142_),
    .X(_00164_));
 sky130_fd_sc_hd__o21ai_1 _12164_ (.A1(_10073_),
    .A2(_00164_),
    .B1(_00153_),
    .Y(_00175_));
 sky130_fd_sc_hd__a21oi_1 _12165_ (.A1(_10073_),
    .A2(_00142_),
    .B1(_00175_),
    .Y(net69));
 sky130_fd_sc_hd__a2bb2oi_1 _12166_ (.A1_N(_10062_),
    .A2_N(_00076_),
    .B1(_10073_),
    .B2(_00098_),
    .Y(_00195_));
 sky130_fd_sc_hd__and2_1 _12167_ (.A(_00195_),
    .B(_00153_),
    .X(_00206_));
 sky130_fd_sc_hd__and2_1 _12168_ (.A(_10400_),
    .B(_10433_),
    .X(_00217_));
 sky130_fd_sc_hd__a21oi_2 _12169_ (.A1(_10400_),
    .A2(_10433_),
    .B1(_10302_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _12170_ (.A(_00217_),
    .B(_10302_),
    .Y(_00239_));
 sky130_fd_sc_hd__and2b_1 _12171_ (.A_N(_00228_),
    .B(_00239_),
    .X(_00250_));
 sky130_fd_sc_hd__nand2b_2 _12172_ (.A_N(_00228_),
    .B(_00239_),
    .Y(_00261_));
 sky130_fd_sc_hd__a31o_1 _12173_ (.A1(_10499_),
    .A2(net63),
    .A3(net28),
    .B1(_10521_),
    .X(_00272_));
 sky130_fd_sc_hd__o21ai_1 _12174_ (.A1(_10839_),
    .A2(_10850_),
    .B1(_10882_),
    .Y(_00283_));
 sky130_fd_sc_hd__o21a_1 _12175_ (.A1(_10839_),
    .A2(_10850_),
    .B1(_10882_),
    .X(_00294_));
 sky130_fd_sc_hd__nand2_2 _12176_ (.A(net62),
    .B(net31),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_4 _12177_ (.A(net61),
    .B(net31),
    .Y(_00316_));
 sky130_fd_sc_hd__a22oi_2 _12178_ (.A1(net30),
    .A2(net62),
    .B1(net31),
    .B2(net61),
    .Y(_00327_));
 sky130_fd_sc_hd__a22o_1 _12179_ (.A1(net30),
    .A2(net62),
    .B1(net31),
    .B2(net61),
    .X(_00338_));
 sky130_fd_sc_hd__o2bb2ai_1 _12180_ (.A1_N(_10510_),
    .A2_N(_00316_),
    .B1(_00305_),
    .B2(_10477_),
    .Y(_00348_));
 sky130_fd_sc_hd__o221ai_4 _12181_ (.A1(_01857_),
    .A2(_01890_),
    .B1(_10477_),
    .B2(_00305_),
    .C1(_00338_),
    .Y(_00359_));
 sky130_fd_sc_hd__nand3_1 _12182_ (.A(_00348_),
    .B(net63),
    .C(net29),
    .Y(_00370_));
 sky130_fd_sc_hd__o21ai_1 _12183_ (.A1(_01857_),
    .A2(_01890_),
    .B1(_00348_),
    .Y(_00381_));
 sky130_fd_sc_hd__o2111ai_1 _12184_ (.A1(_10477_),
    .A2(_00305_),
    .B1(net29),
    .C1(net63),
    .D1(_00338_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand3_2 _12185_ (.A(_00294_),
    .B(_00359_),
    .C(_00370_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand3_2 _12186_ (.A(_00381_),
    .B(_00392_),
    .C(_00283_),
    .Y(_00414_));
 sky130_fd_sc_hd__inv_2 _12187_ (.A(_00414_),
    .Y(_00425_));
 sky130_fd_sc_hd__a22oi_4 _12188_ (.A1(_10532_),
    .A2(_10543_),
    .B1(_00403_),
    .B2(_00414_),
    .Y(_00436_));
 sky130_fd_sc_hd__and4_2 _12189_ (.A(_10532_),
    .B(_10543_),
    .C(_00403_),
    .D(_00414_),
    .X(_00447_));
 sky130_fd_sc_hd__a21o_1 _12190_ (.A1(_00403_),
    .A2(_00414_),
    .B1(_00272_),
    .X(_00458_));
 sky130_fd_sc_hd__a32o_1 _12191_ (.A1(_00294_),
    .A2(_00359_),
    .A3(_00370_),
    .B1(_10543_),
    .B2(_10532_),
    .X(_00469_));
 sky130_fd_sc_hd__o21ai_4 _12192_ (.A1(_00425_),
    .A2(_00469_),
    .B1(_00458_),
    .Y(_00480_));
 sky130_fd_sc_hd__a21oi_2 _12193_ (.A1(_10806_),
    .A2(_10959_),
    .B1(_10817_),
    .Y(_00490_));
 sky130_fd_sc_hd__a21o_2 _12194_ (.A1(_10806_),
    .A2(_10959_),
    .B1(_10817_),
    .X(_00501_));
 sky130_fd_sc_hd__nand2_1 _12195_ (.A(net60),
    .B(net32),
    .Y(_00512_));
 sky130_fd_sc_hd__nand2_1 _12196_ (.A(net58),
    .B(net3),
    .Y(_00523_));
 sky130_fd_sc_hd__a22oi_1 _12197_ (.A1(net59),
    .A2(net2),
    .B1(net3),
    .B2(net58),
    .Y(_00534_));
 sky130_fd_sc_hd__a22o_1 _12198_ (.A1(net59),
    .A2(net2),
    .B1(net3),
    .B2(net58),
    .X(_00545_));
 sky130_fd_sc_hd__nand4_4 _12199_ (.A(net58),
    .B(net59),
    .C(net2),
    .D(net3),
    .Y(_00556_));
 sky130_fd_sc_hd__o211ai_4 _12200_ (.A1(_01835_),
    .A2(_01912_),
    .B1(_00545_),
    .C1(_00556_),
    .Y(_00567_));
 sky130_fd_sc_hd__a21o_1 _12201_ (.A1(_00545_),
    .A2(_00556_),
    .B1(_00512_),
    .X(_00578_));
 sky130_fd_sc_hd__o2bb2a_2 _12202_ (.A1_N(_00545_),
    .A2_N(_00556_),
    .B1(_01835_),
    .B2(_01912_),
    .X(_00589_));
 sky130_fd_sc_hd__and4_2 _12203_ (.A(_00545_),
    .B(_00556_),
    .C(net60),
    .D(net32),
    .X(_00600_));
 sky130_fd_sc_hd__nand2_1 _12204_ (.A(_00567_),
    .B(_00578_),
    .Y(_00611_));
 sky130_fd_sc_hd__a21oi_2 _12205_ (.A1(_09064_),
    .A2(_10707_),
    .B1(_10696_),
    .Y(_00622_));
 sky130_fd_sc_hd__o21ai_2 _12206_ (.A1(_10696_),
    .A2(_10740_),
    .B1(_10729_),
    .Y(_00633_));
 sky130_fd_sc_hd__o31a_2 _12207_ (.A1(_01780_),
    .A2(_01923_),
    .A3(_10740_),
    .B1(_10729_),
    .X(_00643_));
 sky130_fd_sc_hd__nand2_1 _12208_ (.A(net55),
    .B(net4),
    .Y(_00654_));
 sky130_fd_sc_hd__a22oi_4 _12209_ (.A1(net44),
    .A2(net5),
    .B1(net6),
    .B2(net33),
    .Y(_00665_));
 sky130_fd_sc_hd__a22o_1 _12210_ (.A1(net44),
    .A2(net5),
    .B1(net6),
    .B2(net33),
    .X(_00676_));
 sky130_fd_sc_hd__and4_1 _12211_ (.A(net33),
    .B(net44),
    .C(net5),
    .D(net6),
    .X(_00687_));
 sky130_fd_sc_hd__nand4_4 _12212_ (.A(net33),
    .B(net44),
    .C(net5),
    .D(net6),
    .Y(_00698_));
 sky130_fd_sc_hd__o211ai_1 _12213_ (.A1(_01780_),
    .A2(_01945_),
    .B1(_00676_),
    .C1(_00698_),
    .Y(_00709_));
 sky130_fd_sc_hd__a21o_1 _12214_ (.A1(_00676_),
    .A2(_00698_),
    .B1(_00654_),
    .X(_00720_));
 sky130_fd_sc_hd__o22ai_4 _12215_ (.A1(_01780_),
    .A2(_01945_),
    .B1(_00665_),
    .B2(_00687_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand3_2 _12216_ (.A(_00698_),
    .B(net4),
    .C(net55),
    .Y(_00742_));
 sky130_fd_sc_hd__nand4_2 _12217_ (.A(_00676_),
    .B(_00698_),
    .C(net55),
    .D(net4),
    .Y(_00753_));
 sky130_fd_sc_hd__o21ai_2 _12218_ (.A1(_00665_),
    .A2(_00742_),
    .B1(_00731_),
    .Y(_00764_));
 sky130_fd_sc_hd__o221a_4 _12219_ (.A1(_00665_),
    .A2(_00742_),
    .B1(_10718_),
    .B2(_00622_),
    .C1(_00731_),
    .X(_00775_));
 sky130_fd_sc_hd__o221ai_4 _12220_ (.A1(_10718_),
    .A2(_00622_),
    .B1(_00665_),
    .B2(_00742_),
    .C1(_00731_),
    .Y(_00785_));
 sky130_fd_sc_hd__a21oi_2 _12221_ (.A1(_00731_),
    .A2(_00753_),
    .B1(_00633_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand3_2 _12222_ (.A(_00643_),
    .B(_00709_),
    .C(_00720_),
    .Y(_00807_));
 sky130_fd_sc_hd__o2bb2ai_2 _12223_ (.A1_N(_00567_),
    .A2_N(_00578_),
    .B1(_00775_),
    .B2(_00796_),
    .Y(_00818_));
 sky130_fd_sc_hd__o211ai_4 _12224_ (.A1(_00589_),
    .A2(_00600_),
    .B1(_00785_),
    .C1(_00807_),
    .Y(_00829_));
 sky130_fd_sc_hd__a22oi_4 _12225_ (.A1(_00567_),
    .A2(_00578_),
    .B1(_00764_),
    .B2(_00643_),
    .Y(_00840_));
 sky130_fd_sc_hd__o21ai_4 _12226_ (.A1(_00643_),
    .A2(_00764_),
    .B1(_00840_),
    .Y(_00851_));
 sky130_fd_sc_hd__o22ai_4 _12227_ (.A1(_00589_),
    .A2(_00600_),
    .B1(_00775_),
    .B2(_00796_),
    .Y(_00862_));
 sky130_fd_sc_hd__a21oi_2 _12228_ (.A1(_00818_),
    .A2(_00829_),
    .B1(_00490_),
    .Y(_00873_));
 sky130_fd_sc_hd__nand3_2 _12229_ (.A(_00501_),
    .B(_00851_),
    .C(_00862_),
    .Y(_00884_));
 sky130_fd_sc_hd__a21oi_4 _12230_ (.A1(_00851_),
    .A2(_00862_),
    .B1(_00501_),
    .Y(_00895_));
 sky130_fd_sc_hd__nand3_2 _12231_ (.A(_00490_),
    .B(_00818_),
    .C(_00829_),
    .Y(_00906_));
 sky130_fd_sc_hd__a21boi_2 _12232_ (.A1(_00884_),
    .A2(_00906_),
    .B1_N(_00480_),
    .Y(_00917_));
 sky130_fd_sc_hd__o21ai_2 _12233_ (.A1(_00873_),
    .A2(_00895_),
    .B1(_00480_),
    .Y(_00927_));
 sky130_fd_sc_hd__o21ai_2 _12234_ (.A1(_00436_),
    .A2(_00447_),
    .B1(_00906_),
    .Y(_00938_));
 sky130_fd_sc_hd__o211a_1 _12235_ (.A1(_00436_),
    .A2(_00447_),
    .B1(_00884_),
    .C1(_00906_),
    .X(_00949_));
 sky130_fd_sc_hd__a311oi_4 _12236_ (.A1(_00501_),
    .A2(_00851_),
    .A3(_00862_),
    .B1(_00447_),
    .C1(_00436_),
    .Y(_00960_));
 sky130_fd_sc_hd__o21ai_4 _12237_ (.A1(_00480_),
    .A2(_00895_),
    .B1(_00884_),
    .Y(_00971_));
 sky130_fd_sc_hd__a32o_1 _12238_ (.A1(_00490_),
    .A2(_00818_),
    .A3(_00829_),
    .B1(_00884_),
    .B2(_00480_),
    .X(_00982_));
 sky130_fd_sc_hd__nor2_1 _12239_ (.A(_00917_),
    .B(_00949_),
    .Y(_00993_));
 sky130_fd_sc_hd__o21ai_1 _12240_ (.A1(_00873_),
    .A2(_00938_),
    .B1(_00927_),
    .Y(_01004_));
 sky130_fd_sc_hd__a31oi_4 _12241_ (.A1(_10631_),
    .A2(_10641_),
    .A3(_11014_),
    .B1(_11025_),
    .Y(_01015_));
 sky130_fd_sc_hd__inv_2 _12242_ (.A(_01015_),
    .Y(_01026_));
 sky130_fd_sc_hd__o21ai_4 _12243_ (.A1(_00917_),
    .A2(_00949_),
    .B1(_01015_),
    .Y(_01037_));
 sky130_fd_sc_hd__o221a_2 _12244_ (.A1(_00873_),
    .A2(_00938_),
    .B1(_11025_),
    .B2(_11080_),
    .C1(_00927_),
    .X(_01047_));
 sky130_fd_sc_hd__o221ai_4 _12245_ (.A1(_11025_),
    .A2(_11080_),
    .B1(_00873_),
    .B2(_00938_),
    .C1(_00927_),
    .Y(_01058_));
 sky130_fd_sc_hd__a21boi_1 _12246_ (.A1(_10587_),
    .A2(_10620_),
    .B1_N(_10598_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_1 _12247_ (.A(_10598_),
    .B(_10641_),
    .Y(_01080_));
 sky130_fd_sc_hd__o21ai_1 _12248_ (.A1(_01802_),
    .A2(_01934_),
    .B1(_10170_),
    .Y(_01091_));
 sky130_fd_sc_hd__o31a_1 _12249_ (.A1(_01802_),
    .A2(_01934_),
    .A3(_10181_),
    .B1(_10170_),
    .X(_01102_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(net26),
    .B(net35),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _12251_ (.A(net28),
    .B(net64),
    .Y(_01124_));
 sky130_fd_sc_hd__nand4_4 _12252_ (.A(net28),
    .B(net27),
    .C(net64),
    .D(net34),
    .Y(_01135_));
 sky130_fd_sc_hd__a22oi_4 _12253_ (.A1(net28),
    .A2(net64),
    .B1(net34),
    .B2(net27),
    .Y(_01146_));
 sky130_fd_sc_hd__a22o_1 _12254_ (.A1(net28),
    .A2(net64),
    .B1(net34),
    .B2(net27),
    .X(_01157_));
 sky130_fd_sc_hd__o211ai_1 _12255_ (.A1(_01791_),
    .A2(_01934_),
    .B1(_01135_),
    .C1(_01157_),
    .Y(_01167_));
 sky130_fd_sc_hd__a21o_1 _12256_ (.A1(_01135_),
    .A2(_01157_),
    .B1(_01113_),
    .X(_01178_));
 sky130_fd_sc_hd__o2bb2ai_1 _12257_ (.A1_N(_01135_),
    .A2_N(_01157_),
    .B1(_01791_),
    .B2(_01934_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand4_2 _12258_ (.A(_01157_),
    .B(net35),
    .C(net26),
    .D(_01135_),
    .Y(_01200_));
 sky130_fd_sc_hd__and3_2 _12259_ (.A(_01102_),
    .B(_01167_),
    .C(_01178_),
    .X(_01211_));
 sky130_fd_sc_hd__nand3_1 _12260_ (.A(_01102_),
    .B(_01167_),
    .C(_01178_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand4_4 _12261_ (.A(_10192_),
    .B(_01091_),
    .C(_01189_),
    .D(_01200_),
    .Y(_01233_));
 sky130_fd_sc_hd__a22oi_1 _12262_ (.A1(net23),
    .A2(net36),
    .B1(net37),
    .B2(net12),
    .Y(_01244_));
 sky130_fd_sc_hd__a22o_1 _12263_ (.A1(net23),
    .A2(net36),
    .B1(net37),
    .B2(net12),
    .X(_01255_));
 sky130_fd_sc_hd__and4_1 _12264_ (.A(net23),
    .B(net12),
    .C(net36),
    .D(net37),
    .X(_01265_));
 sky130_fd_sc_hd__and4b_1 _12265_ (.A_N(_01265_),
    .B(net38),
    .C(net1),
    .D(_01255_),
    .X(_01276_));
 sky130_fd_sc_hd__nand4b_1 _12266_ (.A_N(_01265_),
    .B(net38),
    .C(net1),
    .D(_01255_),
    .Y(_01287_));
 sky130_fd_sc_hd__o2bb2a_1 _12267_ (.A1_N(net1),
    .A2_N(net38),
    .B1(_01244_),
    .B2(_01265_),
    .X(_01298_));
 sky130_fd_sc_hd__o2bb2ai_1 _12268_ (.A1_N(net1),
    .A2_N(net38),
    .B1(_01244_),
    .B2(_01265_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _12269_ (.A(_01287_),
    .B(_01309_),
    .Y(_01320_));
 sky130_fd_sc_hd__o2bb2ai_1 _12270_ (.A1_N(_01222_),
    .A2_N(_01233_),
    .B1(_01276_),
    .B2(_01298_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand4_1 _12271_ (.A(_01222_),
    .B(_01233_),
    .C(_01287_),
    .D(_01309_),
    .Y(_01342_));
 sky130_fd_sc_hd__a21o_1 _12272_ (.A1(_01222_),
    .A2(_01233_),
    .B1(_01320_),
    .X(_01352_));
 sky130_fd_sc_hd__o211ai_1 _12273_ (.A1(_01276_),
    .A2(_01298_),
    .B1(_01222_),
    .C1(_01233_),
    .Y(_01363_));
 sky130_fd_sc_hd__nand3_2 _12274_ (.A(_01352_),
    .B(_01363_),
    .C(_01069_),
    .Y(_01374_));
 sky130_fd_sc_hd__and3_2 _12275_ (.A(_01080_),
    .B(_01331_),
    .C(_01342_),
    .X(_01385_));
 sky130_fd_sc_hd__nand3_2 _12276_ (.A(_01080_),
    .B(_01331_),
    .C(_01342_),
    .Y(_01396_));
 sky130_fd_sc_hd__o21a_1 _12277_ (.A1(_10291_),
    .A2(_10313_),
    .B1(_10269_),
    .X(_01407_));
 sky130_fd_sc_hd__nor2_1 _12278_ (.A(_10247_),
    .B(_01407_),
    .Y(_01418_));
 sky130_fd_sc_hd__o2bb2ai_2 _12279_ (.A1_N(_01374_),
    .A2_N(_01396_),
    .B1(_01407_),
    .B2(_10247_),
    .Y(_01428_));
 sky130_fd_sc_hd__inv_2 _12280_ (.A(_01428_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_2 _12281_ (.A(_01374_),
    .B(_01418_),
    .Y(_01450_));
 sky130_fd_sc_hd__and3_2 _12282_ (.A(_01374_),
    .B(_01396_),
    .C(_01418_),
    .X(_01461_));
 sky130_fd_sc_hd__o21ai_2 _12283_ (.A1(_01385_),
    .A2(_01450_),
    .B1(_01428_),
    .Y(_01472_));
 sky130_fd_sc_hd__a21oi_2 _12284_ (.A1(_01004_),
    .A2(_01015_),
    .B1(_01472_),
    .Y(_01482_));
 sky130_fd_sc_hd__o211ai_2 _12285_ (.A1(_01385_),
    .A2(_01450_),
    .B1(_01428_),
    .C1(_01037_),
    .Y(_01493_));
 sky130_fd_sc_hd__o21ai_1 _12286_ (.A1(_01004_),
    .A2(_01015_),
    .B1(_01482_),
    .Y(_01504_));
 sky130_fd_sc_hd__o2bb2ai_2 _12287_ (.A1_N(_01037_),
    .A2_N(_01058_),
    .B1(_01439_),
    .B2(_01461_),
    .Y(_01515_));
 sky130_fd_sc_hd__a21o_1 _12288_ (.A1(_01037_),
    .A2(_01058_),
    .B1(_01472_),
    .X(_01526_));
 sky130_fd_sc_hd__o211ai_4 _12289_ (.A1(_01439_),
    .A2(_01461_),
    .B1(_01037_),
    .C1(_01058_),
    .Y(_01536_));
 sky130_fd_sc_hd__a32oi_4 _12290_ (.A1(_10466_),
    .A2(_11047_),
    .A3(_11058_),
    .B1(_11112_),
    .B2(_10444_),
    .Y(_01547_));
 sky130_fd_sc_hd__a32o_1 _12291_ (.A1(_10466_),
    .A2(_11047_),
    .A3(_11058_),
    .B1(_11112_),
    .B2(_10444_),
    .X(_01558_));
 sky130_fd_sc_hd__and3_1 _12292_ (.A(_01526_),
    .B(_01536_),
    .C(_01558_),
    .X(_01569_));
 sky130_fd_sc_hd__nand3_2 _12293_ (.A(_01526_),
    .B(_01536_),
    .C(_01558_),
    .Y(_01579_));
 sky130_fd_sc_hd__o211ai_4 _12294_ (.A1(_01047_),
    .A2(_01493_),
    .B1(_01547_),
    .C1(_01515_),
    .Y(_01590_));
 sky130_fd_sc_hd__a21o_1 _12295_ (.A1(_01579_),
    .A2(_01590_),
    .B1(_00250_),
    .X(_01595_));
 sky130_fd_sc_hd__nand3_1 _12296_ (.A(_01579_),
    .B(_01590_),
    .C(_00250_),
    .Y(_01596_));
 sky130_fd_sc_hd__nand3_1 _12297_ (.A(_00261_),
    .B(_01579_),
    .C(_01590_),
    .Y(_01597_));
 sky130_fd_sc_hd__a21o_1 _12298_ (.A1(_01579_),
    .A2(_01590_),
    .B1(_00261_),
    .X(_01598_));
 sky130_fd_sc_hd__nand4_1 _12299_ (.A(_11200_),
    .B(_11244_),
    .C(_01597_),
    .D(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__o211a_1 _12300_ (.A1(_11189_),
    .A2(_11233_),
    .B1(_01595_),
    .C1(_01596_),
    .X(_01600_));
 sky130_fd_sc_hd__o211ai_1 _12301_ (.A1(_11189_),
    .A2(_11233_),
    .B1(_01595_),
    .C1(_01596_),
    .Y(_01601_));
 sky130_fd_sc_hd__o2bb2a_2 _12302_ (.A1_N(_01599_),
    .A2_N(_01601_),
    .B1(_11233_),
    .B2(_00000_),
    .X(_01602_));
 sky130_fd_sc_hd__and4b_4 _12303_ (.A_N(_00000_),
    .B(_01599_),
    .C(_01601_),
    .D(_11244_),
    .X(_01603_));
 sky130_fd_sc_hd__nor2_1 _12304_ (.A(_01602_),
    .B(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__o2bb2a_1 _12305_ (.A1_N(_00043_),
    .A2_N(_00131_),
    .B1(_01602_),
    .B2(_01603_),
    .X(_01605_));
 sky130_fd_sc_hd__and3_1 _12306_ (.A(_01604_),
    .B(_00131_),
    .C(_00043_),
    .X(_01606_));
 sky130_fd_sc_hd__or2_1 _12307_ (.A(_01605_),
    .B(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__o2bb2ai_1 _12308_ (.A1_N(_00153_),
    .A2_N(_00195_),
    .B1(_01605_),
    .B2(_01606_),
    .Y(_01608_));
 sky130_fd_sc_hd__xnor2_1 _12309_ (.A(_00206_),
    .B(_01607_),
    .Y(net70));
 sky130_fd_sc_hd__o31ai_4 _12310_ (.A1(_00131_),
    .A2(_01602_),
    .A3(_01603_),
    .B1(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__a31oi_2 _12311_ (.A1(_01504_),
    .A2(_01515_),
    .A3(_01547_),
    .B1(_00250_),
    .Y(_01610_));
 sky130_fd_sc_hd__a32oi_4 _12312_ (.A1(_01526_),
    .A2(_01536_),
    .A3(_01558_),
    .B1(_01590_),
    .B2(_00261_),
    .Y(_01611_));
 sky130_fd_sc_hd__a21oi_1 _12313_ (.A1(_01374_),
    .A2(_01418_),
    .B1(_01385_),
    .Y(_01612_));
 sky130_fd_sc_hd__a31o_1 _12314_ (.A1(_01255_),
    .A2(net38),
    .A3(net1),
    .B1(_01265_),
    .X(_01613_));
 sky130_fd_sc_hd__and3_2 _12315_ (.A(_01613_),
    .B(net39),
    .C(net1),
    .X(_01614_));
 sky130_fd_sc_hd__o211ai_2 _12316_ (.A1(_01265_),
    .A2(_01276_),
    .B1(net1),
    .C1(net39),
    .Y(_01615_));
 sky130_fd_sc_hd__a21oi_1 _12317_ (.A1(net1),
    .A2(net39),
    .B1(_01613_),
    .Y(_01616_));
 sky130_fd_sc_hd__or2_2 _12318_ (.A(_01614_),
    .B(_01616_),
    .X(_01617_));
 sky130_fd_sc_hd__inv_2 _12319_ (.A(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__and3_1 _12320_ (.A(_01396_),
    .B(_01450_),
    .C(_01617_),
    .X(_01619_));
 sky130_fd_sc_hd__a211o_1 _12321_ (.A1(_01374_),
    .A2(_01418_),
    .B1(_01618_),
    .C1(_01385_),
    .X(_01620_));
 sky130_fd_sc_hd__a21oi_4 _12322_ (.A1(_01396_),
    .A2(_01450_),
    .B1(_01617_),
    .Y(_01621_));
 sky130_fd_sc_hd__inv_2 _12323_ (.A(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__nor2_1 _12324_ (.A(_01619_),
    .B(_01621_),
    .Y(_01623_));
 sky130_fd_sc_hd__nand2_1 _12325_ (.A(_01620_),
    .B(_01622_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_1 _12326_ (.A(_01058_),
    .B(_01472_),
    .Y(_01625_));
 sky130_fd_sc_hd__o21ai_2 _12327_ (.A1(_00993_),
    .A2(_01026_),
    .B1(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _12328_ (.A(_00414_),
    .B(_00469_),
    .Y(_01627_));
 sky130_fd_sc_hd__a21oi_2 _12329_ (.A1(_00272_),
    .A2(_00403_),
    .B1(_00425_),
    .Y(_01628_));
 sky130_fd_sc_hd__o21a_1 _12330_ (.A1(_01791_),
    .A2(_01934_),
    .B1(_01135_),
    .X(_01629_));
 sky130_fd_sc_hd__o21ai_1 _12331_ (.A1(_01113_),
    .A2(_01146_),
    .B1(_01135_),
    .Y(_01630_));
 sky130_fd_sc_hd__o21a_1 _12332_ (.A1(_01113_),
    .A2(_01146_),
    .B1(_01135_),
    .X(_01631_));
 sky130_fd_sc_hd__a22oi_1 _12333_ (.A1(net29),
    .A2(net64),
    .B1(net34),
    .B2(net28),
    .Y(_01632_));
 sky130_fd_sc_hd__a22o_2 _12334_ (.A1(net29),
    .A2(net64),
    .B1(net34),
    .B2(net28),
    .X(_01633_));
 sky130_fd_sc_hd__nand2_1 _12335_ (.A(net29),
    .B(net34),
    .Y(_01634_));
 sky130_fd_sc_hd__and4_1 _12336_ (.A(net28),
    .B(net29),
    .C(net64),
    .D(net34),
    .X(_01635_));
 sky130_fd_sc_hd__nand4_2 _12337_ (.A(net28),
    .B(net29),
    .C(net64),
    .D(net34),
    .Y(_01636_));
 sky130_fd_sc_hd__a22oi_4 _12338_ (.A1(net27),
    .A2(net35),
    .B1(_01633_),
    .B2(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__a22o_1 _12339_ (.A1(net27),
    .A2(net35),
    .B1(_01633_),
    .B2(_01636_),
    .X(_01638_));
 sky130_fd_sc_hd__o2111a_1 _12340_ (.A1(_01124_),
    .A2(_01634_),
    .B1(net27),
    .C1(net35),
    .D1(_01633_),
    .X(_01639_));
 sky130_fd_sc_hd__o2111ai_1 _12341_ (.A1(_01124_),
    .A2(_01634_),
    .B1(net27),
    .C1(net35),
    .D1(_01633_),
    .Y(_01640_));
 sky130_fd_sc_hd__o22ai_4 _12342_ (.A1(_01146_),
    .A2(_01629_),
    .B1(_01637_),
    .B2(_01639_),
    .Y(_01641_));
 sky130_fd_sc_hd__inv_2 _12343_ (.A(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__and3_1 _12344_ (.A(_01638_),
    .B(_01640_),
    .C(_01630_),
    .X(_01643_));
 sky130_fd_sc_hd__nand3_1 _12345_ (.A(_01638_),
    .B(_01640_),
    .C(_01630_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _12346_ (.A(net12),
    .B(net38),
    .Y(_01645_));
 sky130_fd_sc_hd__a22oi_2 _12347_ (.A1(net26),
    .A2(net36),
    .B1(net37),
    .B2(net23),
    .Y(_01646_));
 sky130_fd_sc_hd__and4_1 _12348_ (.A(net26),
    .B(net23),
    .C(net36),
    .D(net37),
    .X(_01647_));
 sky130_fd_sc_hd__nand4_1 _12349_ (.A(net26),
    .B(net23),
    .C(net36),
    .D(net37),
    .Y(_01648_));
 sky130_fd_sc_hd__nor3_1 _12350_ (.A(_01645_),
    .B(_01646_),
    .C(_01647_),
    .Y(_01649_));
 sky130_fd_sc_hd__o21a_1 _12351_ (.A1(_01646_),
    .A2(_01647_),
    .B1(_01645_),
    .X(_01650_));
 sky130_fd_sc_hd__nor2_1 _12352_ (.A(_01649_),
    .B(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__a21oi_2 _12353_ (.A1(_01641_),
    .A2(_01644_),
    .B1(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__o311a_1 _12354_ (.A1(_01631_),
    .A2(_01637_),
    .A3(_01639_),
    .B1(_01641_),
    .C1(_01651_),
    .X(_01653_));
 sky130_fd_sc_hd__nand3_1 _12355_ (.A(_01651_),
    .B(_01644_),
    .C(_01641_),
    .Y(_01654_));
 sky130_fd_sc_hd__o21ai_4 _12356_ (.A1(_01652_),
    .A2(_01653_),
    .B1(_01628_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand3b_4 _12357_ (.A_N(_01652_),
    .B(_01654_),
    .C(_01627_),
    .Y(_01656_));
 sky130_fd_sc_hd__o21a_1 _12358_ (.A1(_01276_),
    .A2(_01298_),
    .B1(_01233_),
    .X(_01657_));
 sky130_fd_sc_hd__a21oi_4 _12359_ (.A1(_01233_),
    .A2(_01320_),
    .B1(_01211_),
    .Y(_01658_));
 sky130_fd_sc_hd__o2bb2ai_4 _12360_ (.A1_N(_01655_),
    .A2_N(_01656_),
    .B1(_01657_),
    .B2(_01211_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand3_4 _12361_ (.A(_01655_),
    .B(_01656_),
    .C(_01658_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_2 _12362_ (.A(_01659_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__o21ai_1 _12363_ (.A1(_00512_),
    .A2(_00534_),
    .B1(_00556_),
    .Y(_01662_));
 sky130_fd_sc_hd__o21a_1 _12364_ (.A1(_00512_),
    .A2(_00534_),
    .B1(_00556_),
    .X(_01663_));
 sky130_fd_sc_hd__and2_1 _12365_ (.A(net30),
    .B(net63),
    .X(_01664_));
 sky130_fd_sc_hd__nand2_2 _12366_ (.A(net62),
    .B(net32),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_4 _12367_ (.A(net61),
    .B(net32),
    .Y(_01666_));
 sky130_fd_sc_hd__a22o_1 _12368_ (.A1(net62),
    .A2(net31),
    .B1(net32),
    .B2(net61),
    .X(_01667_));
 sky130_fd_sc_hd__o2bb2ai_1 _12369_ (.A1_N(_00305_),
    .A2_N(_01666_),
    .B1(_01665_),
    .B2(_00316_),
    .Y(_01668_));
 sky130_fd_sc_hd__o221ai_4 _12370_ (.A1(_01868_),
    .A2(_01890_),
    .B1(_00316_),
    .B2(_01665_),
    .C1(_01667_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand2_1 _12371_ (.A(_01668_),
    .B(_01664_),
    .Y(_01670_));
 sky130_fd_sc_hd__o21ai_1 _12372_ (.A1(_01868_),
    .A2(_01890_),
    .B1(_01668_),
    .Y(_01671_));
 sky130_fd_sc_hd__o211a_1 _12373_ (.A1(_00316_),
    .A2(_01665_),
    .B1(_01664_),
    .C1(_01667_),
    .X(_01672_));
 sky130_fd_sc_hd__o2111ai_1 _12374_ (.A1(_00316_),
    .A2(_01665_),
    .B1(net30),
    .C1(net63),
    .D1(_01667_),
    .Y(_01673_));
 sky130_fd_sc_hd__nand3_4 _12375_ (.A(_01663_),
    .B(_01669_),
    .C(_01670_),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_1 _12376_ (.A(_01671_),
    .B(_01662_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand3_2 _12377_ (.A(_01671_),
    .B(_01673_),
    .C(_01662_),
    .Y(_01676_));
 sky130_fd_sc_hd__o22a_2 _12378_ (.A1(_01857_),
    .A2(_01890_),
    .B1(_10477_),
    .B2(_00305_),
    .X(_01677_));
 sky130_fd_sc_hd__a21oi_4 _12379_ (.A1(_10510_),
    .A2(_00316_),
    .B1(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__o2bb2a_2 _12380_ (.A1_N(_01674_),
    .A2_N(_01676_),
    .B1(_01677_),
    .B2(_00327_),
    .X(_01679_));
 sky130_fd_sc_hd__o2bb2ai_4 _12381_ (.A1_N(_01674_),
    .A2_N(_01676_),
    .B1(_01677_),
    .B2(_00327_),
    .Y(_01680_));
 sky130_fd_sc_hd__and3_2 _12382_ (.A(_01674_),
    .B(_01676_),
    .C(_01678_),
    .X(_01681_));
 sky130_fd_sc_hd__o211ai_4 _12383_ (.A1(_01672_),
    .A2(_01675_),
    .B1(_01678_),
    .C1(_01674_),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _12384_ (.A(_01680_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__a32o_4 _12385_ (.A1(_00633_),
    .A2(_00731_),
    .A3(_00753_),
    .B1(_00807_),
    .B2(_00611_),
    .X(_01684_));
 sky130_fd_sc_hd__nand2_1 _12386_ (.A(net60),
    .B(net2),
    .Y(_01685_));
 sky130_fd_sc_hd__nand2_1 _12387_ (.A(net59),
    .B(net4),
    .Y(_01686_));
 sky130_fd_sc_hd__nand2_2 _12388_ (.A(net58),
    .B(net4),
    .Y(_01687_));
 sky130_fd_sc_hd__nand4_2 _12389_ (.A(net58),
    .B(net59),
    .C(net3),
    .D(net4),
    .Y(_01688_));
 sky130_fd_sc_hd__a22o_2 _12390_ (.A1(net59),
    .A2(net3),
    .B1(net4),
    .B2(net58),
    .X(_01689_));
 sky130_fd_sc_hd__o221a_2 _12391_ (.A1(_01835_),
    .A2(_01901_),
    .B1(_00523_),
    .B2(_01686_),
    .C1(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__a21oi_2 _12392_ (.A1(_01688_),
    .A2(_01689_),
    .B1(_01685_),
    .Y(_01691_));
 sky130_fd_sc_hd__a2bb2oi_2 _12393_ (.A1_N(_01835_),
    .A2_N(_01901_),
    .B1(_01688_),
    .B2(_01689_),
    .Y(_01692_));
 sky130_fd_sc_hd__o2111a_1 _12394_ (.A1(_00523_),
    .A2(_01686_),
    .B1(net60),
    .C1(net2),
    .D1(_01689_),
    .X(_01693_));
 sky130_fd_sc_hd__nor2_1 _12395_ (.A(_01692_),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__o21ai_4 _12396_ (.A1(_00654_),
    .A2(_00665_),
    .B1(_00698_),
    .Y(_01695_));
 sky130_fd_sc_hd__o21a_2 _12397_ (.A1(_00654_),
    .A2(_00665_),
    .B1(_00698_),
    .X(_01696_));
 sky130_fd_sc_hd__nand2_2 _12398_ (.A(net55),
    .B(net5),
    .Y(_01697_));
 sky130_fd_sc_hd__a22oi_4 _12399_ (.A1(net44),
    .A2(net6),
    .B1(net7),
    .B2(net33),
    .Y(_01698_));
 sky130_fd_sc_hd__a22o_1 _12400_ (.A1(net44),
    .A2(net6),
    .B1(net7),
    .B2(net33),
    .X(_01699_));
 sky130_fd_sc_hd__and4_1 _12401_ (.A(net33),
    .B(net44),
    .C(net6),
    .D(net7),
    .X(_01700_));
 sky130_fd_sc_hd__nand4_4 _12402_ (.A(net33),
    .B(net44),
    .C(net6),
    .D(net7),
    .Y(_01701_));
 sky130_fd_sc_hd__o211ai_1 _12403_ (.A1(_01780_),
    .A2(_01956_),
    .B1(_01699_),
    .C1(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__o21bai_1 _12404_ (.A1(_01698_),
    .A2(_01700_),
    .B1_N(_01697_),
    .Y(_01703_));
 sky130_fd_sc_hd__o22a_1 _12405_ (.A1(_01780_),
    .A2(_01956_),
    .B1(_01698_),
    .B2(_01700_),
    .X(_01704_));
 sky130_fd_sc_hd__o22ai_4 _12406_ (.A1(_01780_),
    .A2(_01956_),
    .B1(_01698_),
    .B2(_01700_),
    .Y(_01705_));
 sky130_fd_sc_hd__a41o_2 _12407_ (.A1(net33),
    .A2(net44),
    .A3(net6),
    .A4(net7),
    .B1(_01697_),
    .X(_01706_));
 sky130_fd_sc_hd__nand4_1 _12408_ (.A(_01699_),
    .B(_01701_),
    .C(net55),
    .D(net5),
    .Y(_01707_));
 sky130_fd_sc_hd__o21ai_2 _12409_ (.A1(_01698_),
    .A2(_01706_),
    .B1(_01705_),
    .Y(_01708_));
 sky130_fd_sc_hd__o21ai_1 _12410_ (.A1(_01698_),
    .A2(_01706_),
    .B1(_01695_),
    .Y(_01709_));
 sky130_fd_sc_hd__o211a_4 _12411_ (.A1(_01698_),
    .A2(_01706_),
    .B1(_01695_),
    .C1(_01705_),
    .X(_01710_));
 sky130_fd_sc_hd__o211ai_4 _12412_ (.A1(_01698_),
    .A2(_01706_),
    .B1(_01695_),
    .C1(_01705_),
    .Y(_01711_));
 sky130_fd_sc_hd__a21oi_1 _12413_ (.A1(_01705_),
    .A2(_01707_),
    .B1(_01695_),
    .Y(_01712_));
 sky130_fd_sc_hd__nand3_2 _12414_ (.A(_01696_),
    .B(_01702_),
    .C(_01703_),
    .Y(_01713_));
 sky130_fd_sc_hd__a2bb2oi_4 _12415_ (.A1_N(_01690_),
    .A2_N(_01691_),
    .B1(_01696_),
    .B2(_01708_),
    .Y(_01714_));
 sky130_fd_sc_hd__o21ai_4 _12416_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01713_),
    .Y(_01715_));
 sky130_fd_sc_hd__o21ai_2 _12417_ (.A1(_01696_),
    .A2(_01708_),
    .B1(_01714_),
    .Y(_01716_));
 sky130_fd_sc_hd__a2bb2oi_1 _12418_ (.A1_N(_01692_),
    .A2_N(_01693_),
    .B1(_01711_),
    .B2(_01713_),
    .Y(_01717_));
 sky130_fd_sc_hd__o22ai_4 _12419_ (.A1(_01692_),
    .A2(_01693_),
    .B1(_01710_),
    .B2(_01712_),
    .Y(_01718_));
 sky130_fd_sc_hd__a21oi_4 _12420_ (.A1(_01711_),
    .A2(_01714_),
    .B1(_01717_),
    .Y(_01719_));
 sky130_fd_sc_hd__a21oi_4 _12421_ (.A1(_01716_),
    .A2(_01718_),
    .B1(_01684_),
    .Y(_01720_));
 sky130_fd_sc_hd__a21o_1 _12422_ (.A1(_01716_),
    .A2(_01718_),
    .B1(_01684_),
    .X(_01721_));
 sky130_fd_sc_hd__o221a_4 _12423_ (.A1(_01710_),
    .A2(_01715_),
    .B1(_00775_),
    .B2(_00840_),
    .C1(_01718_),
    .X(_01722_));
 sky130_fd_sc_hd__o221ai_4 _12424_ (.A1(_01710_),
    .A2(_01715_),
    .B1(_00775_),
    .B2(_00840_),
    .C1(_01718_),
    .Y(_01723_));
 sky130_fd_sc_hd__o211ai_4 _12425_ (.A1(_01679_),
    .A2(_01681_),
    .B1(_01721_),
    .C1(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__o21bai_4 _12426_ (.A1(_01720_),
    .A2(_01722_),
    .B1_N(_01683_),
    .Y(_01725_));
 sky130_fd_sc_hd__o22ai_4 _12427_ (.A1(_01679_),
    .A2(_01681_),
    .B1(_01720_),
    .B2(_01722_),
    .Y(_01726_));
 sky130_fd_sc_hd__o21bai_4 _12428_ (.A1(_01684_),
    .A2(_01719_),
    .B1_N(_01683_),
    .Y(_01727_));
 sky130_fd_sc_hd__o2111ai_4 _12429_ (.A1(_01684_),
    .A2(_01719_),
    .B1(_01723_),
    .C1(_01682_),
    .D1(_01680_),
    .Y(_01728_));
 sky130_fd_sc_hd__o211a_1 _12430_ (.A1(_00895_),
    .A2(_00960_),
    .B1(_01724_),
    .C1(_01725_),
    .X(_01729_));
 sky130_fd_sc_hd__o211ai_4 _12431_ (.A1(_00895_),
    .A2(_00960_),
    .B1(_01724_),
    .C1(_01725_),
    .Y(_01730_));
 sky130_fd_sc_hd__o211ai_4 _12432_ (.A1(_01722_),
    .A2(_01727_),
    .B1(_00971_),
    .C1(_01726_),
    .Y(_01731_));
 sky130_fd_sc_hd__nand4_2 _12433_ (.A(_01659_),
    .B(_01660_),
    .C(_01730_),
    .D(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__a22o_1 _12434_ (.A1(_01659_),
    .A2(_01660_),
    .B1(_01730_),
    .B2(_01731_),
    .X(_01733_));
 sky130_fd_sc_hd__a21o_1 _12435_ (.A1(_01730_),
    .A2(_01731_),
    .B1(_01661_),
    .X(_01734_));
 sky130_fd_sc_hd__nand3_2 _12436_ (.A(_01661_),
    .B(_01730_),
    .C(_01731_),
    .Y(_01735_));
 sky130_fd_sc_hd__o211a_1 _12437_ (.A1(_01047_),
    .A2(_01482_),
    .B1(_01732_),
    .C1(_01733_),
    .X(_01736_));
 sky130_fd_sc_hd__o211ai_4 _12438_ (.A1(_01047_),
    .A2(_01482_),
    .B1(_01732_),
    .C1(_01733_),
    .Y(_01738_));
 sky130_fd_sc_hd__nand3_2 _12439_ (.A(_01734_),
    .B(_01735_),
    .C(_01626_),
    .Y(_01739_));
 sky130_fd_sc_hd__a31o_1 _12440_ (.A1(_01626_),
    .A2(_01734_),
    .A3(_01735_),
    .B1(_01624_),
    .X(_01740_));
 sky130_fd_sc_hd__nand4_1 _12441_ (.A(_01620_),
    .B(_01622_),
    .C(_01738_),
    .D(_01739_),
    .Y(_01741_));
 sky130_fd_sc_hd__a22o_1 _12442_ (.A1(_01620_),
    .A2(_01622_),
    .B1(_01738_),
    .B2(_01739_),
    .X(_01742_));
 sky130_fd_sc_hd__o211ai_2 _12443_ (.A1(_01619_),
    .A2(_01621_),
    .B1(_01738_),
    .C1(_01739_),
    .Y(_01743_));
 sky130_fd_sc_hd__a21o_1 _12444_ (.A1(_01738_),
    .A2(_01739_),
    .B1(_01624_),
    .X(_01744_));
 sky130_fd_sc_hd__and3_1 _12445_ (.A(_01742_),
    .B(_01611_),
    .C(_01741_),
    .X(_01745_));
 sky130_fd_sc_hd__o211ai_2 _12446_ (.A1(_01736_),
    .A2(_01740_),
    .B1(_01611_),
    .C1(_01742_),
    .Y(_01746_));
 sky130_fd_sc_hd__o211ai_4 _12447_ (.A1(_01569_),
    .A2(_01610_),
    .B1(_01743_),
    .C1(_01744_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_1 _12448_ (.A(_01747_),
    .B(_00228_),
    .Y(_01749_));
 sky130_fd_sc_hd__nand3_1 _12449_ (.A(_01747_),
    .B(_00228_),
    .C(_01746_),
    .Y(_01750_));
 sky130_fd_sc_hd__o2bb2ai_2 _12450_ (.A1_N(_01746_),
    .A2_N(_01747_),
    .B1(_10302_),
    .B2(_00217_),
    .Y(_01751_));
 sky130_fd_sc_hd__o21ai_1 _12451_ (.A1(_01745_),
    .A2(_01749_),
    .B1(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__and3_1 _12452_ (.A(_01751_),
    .B(_01600_),
    .C(_01750_),
    .X(_01753_));
 sky130_fd_sc_hd__o211ai_1 _12453_ (.A1(_01745_),
    .A2(_01749_),
    .B1(_01600_),
    .C1(_01751_),
    .Y(_01754_));
 sky130_fd_sc_hd__a21oi_1 _12454_ (.A1(_01750_),
    .A2(_01751_),
    .B1(_01600_),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_2 _12455_ (.A(_01753_),
    .B(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__or2_2 _12456_ (.A(_01753_),
    .B(_01755_),
    .X(_01757_));
 sky130_fd_sc_hd__or3_2 _12457_ (.A(_00043_),
    .B(_01602_),
    .C(_01603_),
    .X(_01758_));
 sky130_fd_sc_hd__o21ba_1 _12458_ (.A1(_00043_),
    .A2(_01602_),
    .B1_N(_01603_),
    .X(_01760_));
 sky130_fd_sc_hd__xnor2_4 _12459_ (.A(_01756_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__xor2_1 _12460_ (.A(_01609_),
    .B(_01761_),
    .X(net71));
 sky130_fd_sc_hd__a2bb2oi_4 _12461_ (.A1_N(_01757_),
    .A2_N(_01758_),
    .B1(_01761_),
    .B2(_01609_),
    .Y(_01762_));
 sky130_fd_sc_hd__o2bb2ai_4 _12462_ (.A1_N(_01609_),
    .A2_N(_01761_),
    .B1(_01758_),
    .B2(_01757_),
    .Y(_01763_));
 sky130_fd_sc_hd__a31o_1 _12463_ (.A1(_01742_),
    .A2(_01611_),
    .A3(_01741_),
    .B1(_00228_),
    .X(_01764_));
 sky130_fd_sc_hd__a21oi_1 _12464_ (.A1(_00228_),
    .A2(_01747_),
    .B1(_01745_),
    .Y(_01765_));
 sky130_fd_sc_hd__a32oi_4 _12465_ (.A1(_01626_),
    .A2(_01734_),
    .A3(_01735_),
    .B1(_01738_),
    .B2(_01624_),
    .Y(_01766_));
 sky130_fd_sc_hd__a21oi_2 _12466_ (.A1(_01739_),
    .A2(_01623_),
    .B1(_01736_),
    .Y(_01767_));
 sky130_fd_sc_hd__a21boi_4 _12467_ (.A1(_01655_),
    .A2(_01658_),
    .B1_N(_01656_),
    .Y(_01768_));
 sky130_fd_sc_hd__a22o_1 _12468_ (.A1(net12),
    .A2(net39),
    .B1(net40),
    .B2(net1),
    .X(_01770_));
 sky130_fd_sc_hd__and4_1 _12469_ (.A(net12),
    .B(net1),
    .C(net39),
    .D(net40),
    .X(_01771_));
 sky130_fd_sc_hd__nand4_4 _12470_ (.A(net12),
    .B(net1),
    .C(net39),
    .D(net40),
    .Y(_01772_));
 sky130_fd_sc_hd__o21ai_2 _12471_ (.A1(_01645_),
    .A2(_01646_),
    .B1(_01648_),
    .Y(_01773_));
 sky130_fd_sc_hd__a21oi_1 _12472_ (.A1(_01770_),
    .A2(_01772_),
    .B1(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__and3_2 _12473_ (.A(_01770_),
    .B(_01772_),
    .C(_01773_),
    .X(_01775_));
 sky130_fd_sc_hd__nand3_2 _12474_ (.A(_01770_),
    .B(_01772_),
    .C(_01773_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor2_2 _12475_ (.A(_01774_),
    .B(_01775_),
    .Y(_01777_));
 sky130_fd_sc_hd__inv_2 _12476_ (.A(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__or3_2 _12477_ (.A(_01774_),
    .B(_01775_),
    .C(_01615_),
    .X(_01779_));
 sky130_fd_sc_hd__a31o_1 _12478_ (.A1(net1),
    .A2(net39),
    .A3(_01613_),
    .B1(_01777_),
    .X(_01781_));
 sky130_fd_sc_hd__nand2_2 _12479_ (.A(_01779_),
    .B(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__a21oi_4 _12480_ (.A1(_01656_),
    .A2(_01660_),
    .B1(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__o311a_2 _12481_ (.A1(_01628_),
    .A2(_01652_),
    .A3(_01653_),
    .B1(_01660_),
    .C1(_01782_),
    .X(_01784_));
 sky130_fd_sc_hd__a21oi_2 _12482_ (.A1(_01779_),
    .A2(_01781_),
    .B1(_01768_),
    .Y(_01785_));
 sky130_fd_sc_hd__and3_1 _12483_ (.A(_01768_),
    .B(_01779_),
    .C(_01781_),
    .X(_01786_));
 sky130_fd_sc_hd__nor2_1 _12484_ (.A(_01783_),
    .B(_01784_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _12485_ (.A(_01785_),
    .B(_01786_),
    .Y(_01788_));
 sky130_fd_sc_hd__a32oi_4 _12486_ (.A1(_00971_),
    .A2(_01726_),
    .A3(_01728_),
    .B1(_01659_),
    .B2(_01660_),
    .Y(_01789_));
 sky130_fd_sc_hd__a32oi_4 _12487_ (.A1(_00982_),
    .A2(_01724_),
    .A3(_01725_),
    .B1(_01731_),
    .B2(_01661_),
    .Y(_01790_));
 sky130_fd_sc_hd__a21boi_4 _12488_ (.A1(_01674_),
    .A2(_01678_),
    .B1_N(_01676_),
    .Y(_01792_));
 sky130_fd_sc_hd__a2bb2o_1 _12489_ (.A1_N(_01672_),
    .A2_N(_01675_),
    .B1(_01678_),
    .B2(_01674_),
    .X(_01793_));
 sky130_fd_sc_hd__a31o_1 _12490_ (.A1(_01633_),
    .A2(net35),
    .A3(net27),
    .B1(_01635_),
    .X(_01794_));
 sky130_fd_sc_hd__o32a_1 _12491_ (.A1(_01769_),
    .A2(_01934_),
    .A3(_01632_),
    .B1(_01634_),
    .B2(_01124_),
    .X(_01795_));
 sky130_fd_sc_hd__nand2_1 _12492_ (.A(net28),
    .B(net35),
    .Y(_01796_));
 sky130_fd_sc_hd__nand4_4 _12493_ (.A(net29),
    .B(net30),
    .C(net64),
    .D(net34),
    .Y(_01797_));
 sky130_fd_sc_hd__a22oi_1 _12494_ (.A1(net30),
    .A2(net64),
    .B1(net34),
    .B2(net29),
    .Y(_01798_));
 sky130_fd_sc_hd__a22o_1 _12495_ (.A1(net30),
    .A2(net64),
    .B1(net34),
    .B2(net29),
    .X(_01799_));
 sky130_fd_sc_hd__o211ai_2 _12496_ (.A1(_01748_),
    .A2(_01934_),
    .B1(_01797_),
    .C1(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__a21o_1 _12497_ (.A1(_01797_),
    .A2(_01799_),
    .B1(_01796_),
    .X(_01801_));
 sky130_fd_sc_hd__a22o_1 _12498_ (.A1(net28),
    .A2(net35),
    .B1(_01797_),
    .B2(_01799_),
    .X(_01803_));
 sky130_fd_sc_hd__nand4_2 _12499_ (.A(_01799_),
    .B(net35),
    .C(net28),
    .D(_01797_),
    .Y(_01804_));
 sky130_fd_sc_hd__nand3_2 _12500_ (.A(_01795_),
    .B(_01800_),
    .C(_01801_),
    .Y(_01805_));
 sky130_fd_sc_hd__nand3_4 _12501_ (.A(_01794_),
    .B(_01803_),
    .C(_01804_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _12502_ (.A(net23),
    .B(net38),
    .Y(_01807_));
 sky130_fd_sc_hd__nand2_1 _12503_ (.A(net27),
    .B(net36),
    .Y(_01808_));
 sky130_fd_sc_hd__a22oi_2 _12504_ (.A1(net27),
    .A2(net36),
    .B1(net37),
    .B2(net26),
    .Y(_01809_));
 sky130_fd_sc_hd__a22o_1 _12505_ (.A1(net27),
    .A2(net36),
    .B1(net37),
    .B2(net26),
    .X(_01810_));
 sky130_fd_sc_hd__and4_1 _12506_ (.A(net27),
    .B(net26),
    .C(net36),
    .D(net37),
    .X(_01811_));
 sky130_fd_sc_hd__nand4_2 _12507_ (.A(net27),
    .B(net26),
    .C(net36),
    .D(net37),
    .Y(_01812_));
 sky130_fd_sc_hd__and3_1 _12508_ (.A(_01807_),
    .B(_01810_),
    .C(_01812_),
    .X(_01814_));
 sky130_fd_sc_hd__a211o_1 _12509_ (.A1(net23),
    .A2(net38),
    .B1(_01809_),
    .C1(_01811_),
    .X(_01815_));
 sky130_fd_sc_hd__o211a_1 _12510_ (.A1(_01809_),
    .A2(_01811_),
    .B1(net23),
    .C1(net38),
    .X(_01816_));
 sky130_fd_sc_hd__a21o_1 _12511_ (.A1(_01810_),
    .A2(_01812_),
    .B1(_01807_),
    .X(_01817_));
 sky130_fd_sc_hd__o2bb2a_1 _12512_ (.A1_N(net23),
    .A2_N(net38),
    .B1(_01809_),
    .B2(_01811_),
    .X(_01818_));
 sky130_fd_sc_hd__and4_1 _12513_ (.A(_01810_),
    .B(_01812_),
    .C(net23),
    .D(net38),
    .X(_01819_));
 sky130_fd_sc_hd__o2bb2ai_2 _12514_ (.A1_N(_01805_),
    .A2_N(_01806_),
    .B1(_01814_),
    .B2(_01816_),
    .Y(_01820_));
 sky130_fd_sc_hd__o211ai_4 _12515_ (.A1(_01818_),
    .A2(_01819_),
    .B1(_01805_),
    .C1(_01806_),
    .Y(_01821_));
 sky130_fd_sc_hd__o2bb2ai_1 _12516_ (.A1_N(_01805_),
    .A2_N(_01806_),
    .B1(_01818_),
    .B2(_01819_),
    .Y(_01822_));
 sky130_fd_sc_hd__a32o_1 _12517_ (.A1(_01795_),
    .A2(_01800_),
    .A3(_01801_),
    .B1(_01815_),
    .B2(_01817_),
    .X(_01823_));
 sky130_fd_sc_hd__o211ai_1 _12518_ (.A1(_01814_),
    .A2(_01816_),
    .B1(_01805_),
    .C1(_01806_),
    .Y(_01825_));
 sky130_fd_sc_hd__nand3_1 _12519_ (.A(_01820_),
    .B(_01821_),
    .C(_01792_),
    .Y(_01826_));
 sky130_fd_sc_hd__a21oi_4 _12520_ (.A1(_01820_),
    .A2(_01821_),
    .B1(_01792_),
    .Y(_01827_));
 sky130_fd_sc_hd__nand3_2 _12521_ (.A(_01793_),
    .B(_01822_),
    .C(_01825_),
    .Y(_01828_));
 sky130_fd_sc_hd__o32a_1 _12522_ (.A1(_01637_),
    .A2(_01639_),
    .A3(_01631_),
    .B1(_01649_),
    .B2(_01650_),
    .X(_01829_));
 sky130_fd_sc_hd__a21o_1 _12523_ (.A1(_01651_),
    .A2(_01641_),
    .B1(_01643_),
    .X(_01830_));
 sky130_fd_sc_hd__a21oi_1 _12524_ (.A1(_01651_),
    .A2(_01641_),
    .B1(_01643_),
    .Y(_01831_));
 sky130_fd_sc_hd__o2bb2a_1 _12525_ (.A1_N(_01826_),
    .A2_N(_01828_),
    .B1(_01829_),
    .B2(_01642_),
    .X(_01832_));
 sky130_fd_sc_hd__o2bb2ai_1 _12526_ (.A1_N(_01826_),
    .A2_N(_01828_),
    .B1(_01829_),
    .B2(_01642_),
    .Y(_01833_));
 sky130_fd_sc_hd__a31oi_2 _12527_ (.A1(_01820_),
    .A2(_01821_),
    .A3(_01792_),
    .B1(_01831_),
    .Y(_01834_));
 sky130_fd_sc_hd__a31o_1 _12528_ (.A1(_01820_),
    .A2(_01821_),
    .A3(_01792_),
    .B1(_01831_),
    .X(_01836_));
 sky130_fd_sc_hd__and3_1 _12529_ (.A(_01826_),
    .B(_01828_),
    .C(_01830_),
    .X(_01837_));
 sky130_fd_sc_hd__o21a_1 _12530_ (.A1(_01827_),
    .A2(_01836_),
    .B1(_01833_),
    .X(_01838_));
 sky130_fd_sc_hd__o21ai_2 _12531_ (.A1(_01827_),
    .A2(_01836_),
    .B1(_01833_),
    .Y(_01839_));
 sky130_fd_sc_hd__a22oi_4 _12532_ (.A1(_01680_),
    .A2(_01682_),
    .B1(_01719_),
    .B2(_01684_),
    .Y(_01840_));
 sky130_fd_sc_hd__a32o_1 _12533_ (.A1(_01684_),
    .A2(_01716_),
    .A3(_01718_),
    .B1(_01682_),
    .B2(_01680_),
    .X(_01841_));
 sky130_fd_sc_hd__a2bb2o_2 _12534_ (.A1_N(_00316_),
    .A2_N(_01665_),
    .B1(_01664_),
    .B2(_01667_),
    .X(_01842_));
 sky130_fd_sc_hd__o2bb2a_1 _12535_ (.A1_N(_01664_),
    .A2_N(_01667_),
    .B1(_01665_),
    .B2(_00316_),
    .X(_01843_));
 sky130_fd_sc_hd__o21ai_2 _12536_ (.A1(_00523_),
    .A2(_01686_),
    .B1(_01685_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_2 _12537_ (.A(_01689_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand2_4 _12538_ (.A(net62),
    .B(net2),
    .Y(_01847_));
 sky130_fd_sc_hd__and4_2 _12539_ (.A(net61),
    .B(net62),
    .C(net2),
    .D(net32),
    .X(_01848_));
 sky130_fd_sc_hd__nand2_2 _12540_ (.A(net61),
    .B(net2),
    .Y(_01849_));
 sky130_fd_sc_hd__a22oi_2 _12541_ (.A1(net61),
    .A2(net2),
    .B1(net32),
    .B2(net62),
    .Y(_01850_));
 sky130_fd_sc_hd__a22o_2 _12542_ (.A1(net61),
    .A2(net2),
    .B1(net32),
    .B2(net62),
    .X(_01851_));
 sky130_fd_sc_hd__o2bb2ai_2 _12543_ (.A1_N(_01665_),
    .A2_N(_01849_),
    .B1(_01847_),
    .B2(_01666_),
    .Y(_01852_));
 sky130_fd_sc_hd__o221ai_4 _12544_ (.A1(_01879_),
    .A2(_01890_),
    .B1(_01666_),
    .B2(_01847_),
    .C1(_01851_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand3_4 _12545_ (.A(_01852_),
    .B(net63),
    .C(net31),
    .Y(_01854_));
 sky130_fd_sc_hd__o2111ai_4 _12546_ (.A1(_01666_),
    .A2(_01847_),
    .B1(net31),
    .C1(net63),
    .D1(_01851_),
    .Y(_01855_));
 sky130_fd_sc_hd__o21ai_1 _12547_ (.A1(_01879_),
    .A2(_01890_),
    .B1(_01852_),
    .Y(_01856_));
 sky130_fd_sc_hd__a21oi_4 _12548_ (.A1(_01853_),
    .A2(_01854_),
    .B1(_01845_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand4_4 _12549_ (.A(_01689_),
    .B(_01844_),
    .C(_01855_),
    .D(_01856_),
    .Y(_01859_));
 sky130_fd_sc_hd__nand3_2 _12550_ (.A(_01845_),
    .B(_01853_),
    .C(_01854_),
    .Y(_01860_));
 sky130_fd_sc_hd__a31oi_4 _12551_ (.A1(_01845_),
    .A2(_01853_),
    .A3(_01854_),
    .B1(_01843_),
    .Y(_01861_));
 sky130_fd_sc_hd__a31o_1 _12552_ (.A1(_01845_),
    .A2(_01853_),
    .A3(_01854_),
    .B1(_01843_),
    .X(_01862_));
 sky130_fd_sc_hd__and3_2 _12553_ (.A(_01859_),
    .B(_01860_),
    .C(_01842_),
    .X(_01863_));
 sky130_fd_sc_hd__a21oi_4 _12554_ (.A1(_01859_),
    .A2(_01860_),
    .B1(_01842_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21o_1 _12555_ (.A1(_01859_),
    .A2(_01860_),
    .B1(_01842_),
    .X(_01865_));
 sky130_fd_sc_hd__a21oi_1 _12556_ (.A1(_01859_),
    .A2(_01861_),
    .B1(_01864_),
    .Y(_01866_));
 sky130_fd_sc_hd__o21ai_4 _12557_ (.A1(_01858_),
    .A2(_01862_),
    .B1(_01865_),
    .Y(_01867_));
 sky130_fd_sc_hd__o21ai_4 _12558_ (.A1(_01697_),
    .A2(_01698_),
    .B1(_01701_),
    .Y(_01869_));
 sky130_fd_sc_hd__o21a_1 _12559_ (.A1(_01697_),
    .A2(_01698_),
    .B1(_01701_),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_1 _12560_ (.A(net55),
    .B(net6),
    .Y(_01871_));
 sky130_fd_sc_hd__a22oi_4 _12561_ (.A1(net44),
    .A2(net7),
    .B1(net8),
    .B2(net33),
    .Y(_01872_));
 sky130_fd_sc_hd__a22o_2 _12562_ (.A1(net44),
    .A2(net7),
    .B1(net8),
    .B2(net33),
    .X(_01873_));
 sky130_fd_sc_hd__and4_1 _12563_ (.A(net33),
    .B(net44),
    .C(net7),
    .D(net8),
    .X(_01874_));
 sky130_fd_sc_hd__nand4_4 _12564_ (.A(net33),
    .B(net44),
    .C(net7),
    .D(net8),
    .Y(_01875_));
 sky130_fd_sc_hd__o211ai_4 _12565_ (.A1(_01780_),
    .A2(_01966_),
    .B1(_01873_),
    .C1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__o21bai_4 _12566_ (.A1(_01872_),
    .A2(_01874_),
    .B1_N(_01871_),
    .Y(_01877_));
 sky130_fd_sc_hd__o22a_2 _12567_ (.A1(_01780_),
    .A2(_01966_),
    .B1(_01872_),
    .B2(_01874_),
    .X(_01878_));
 sky130_fd_sc_hd__a22o_1 _12568_ (.A1(net55),
    .A2(net6),
    .B1(_01873_),
    .B2(_01875_),
    .X(_01880_));
 sky130_fd_sc_hd__a41o_2 _12569_ (.A1(net33),
    .A2(net44),
    .A3(net7),
    .A4(net8),
    .B1(_01871_),
    .X(_01881_));
 sky130_fd_sc_hd__nand3_4 _12570_ (.A(_01870_),
    .B(_01876_),
    .C(_01877_),
    .Y(_01882_));
 sky130_fd_sc_hd__o21ai_4 _12571_ (.A1(_01872_),
    .A2(_01881_),
    .B1(_01869_),
    .Y(_01883_));
 sky130_fd_sc_hd__o211a_1 _12572_ (.A1(_01872_),
    .A2(_01881_),
    .B1(_01869_),
    .C1(_01880_),
    .X(_01884_));
 sky130_fd_sc_hd__o211ai_4 _12573_ (.A1(_01872_),
    .A2(_01881_),
    .B1(_01869_),
    .C1(_01880_),
    .Y(_01885_));
 sky130_fd_sc_hd__nor2_1 _12574_ (.A(_01835_),
    .B(_01923_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _12575_ (.A(net60),
    .B(net3),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_2 _12576_ (.A(net59),
    .B(net5),
    .Y(_01888_));
 sky130_fd_sc_hd__and4_1 _12577_ (.A(net58),
    .B(net59),
    .C(net4),
    .D(net5),
    .X(_01889_));
 sky130_fd_sc_hd__a22oi_4 _12578_ (.A1(net59),
    .A2(net4),
    .B1(net5),
    .B2(net58),
    .Y(_01891_));
 sky130_fd_sc_hd__a22o_1 _12579_ (.A1(net59),
    .A2(net4),
    .B1(net5),
    .B2(net58),
    .X(_01892_));
 sky130_fd_sc_hd__o221a_1 _12580_ (.A1(_01835_),
    .A2(_01923_),
    .B1(_01687_),
    .B2(_01888_),
    .C1(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__o221ai_4 _12581_ (.A1(_01835_),
    .A2(_01923_),
    .B1(_01687_),
    .B2(_01888_),
    .C1(_01892_),
    .Y(_01894_));
 sky130_fd_sc_hd__o211a_1 _12582_ (.A1(_01889_),
    .A2(_01891_),
    .B1(net60),
    .C1(net3),
    .X(_01895_));
 sky130_fd_sc_hd__o21ai_2 _12583_ (.A1(_01889_),
    .A2(_01891_),
    .B1(_01886_),
    .Y(_01896_));
 sky130_fd_sc_hd__o22a_2 _12584_ (.A1(_01835_),
    .A2(_01923_),
    .B1(_01889_),
    .B2(_01891_),
    .X(_01897_));
 sky130_fd_sc_hd__o311a_2 _12585_ (.A1(_01813_),
    .A2(_01956_),
    .A3(_01687_),
    .B1(_01892_),
    .C1(_01886_),
    .X(_01898_));
 sky130_fd_sc_hd__nand2_2 _12586_ (.A(_01894_),
    .B(_01896_),
    .Y(_01899_));
 sky130_fd_sc_hd__o2bb2ai_2 _12587_ (.A1_N(_01882_),
    .A2_N(_01885_),
    .B1(_01893_),
    .B2(_01895_),
    .Y(_01900_));
 sky130_fd_sc_hd__o221ai_4 _12588_ (.A1(_01878_),
    .A2(_01883_),
    .B1(_01897_),
    .B2(_01898_),
    .C1(_01882_),
    .Y(_01902_));
 sky130_fd_sc_hd__o2bb2ai_4 _12589_ (.A1_N(_01882_),
    .A2_N(_01885_),
    .B1(_01897_),
    .B2(_01898_),
    .Y(_01903_));
 sky130_fd_sc_hd__a32oi_4 _12590_ (.A1(_01870_),
    .A2(_01876_),
    .A3(_01877_),
    .B1(_01894_),
    .B2(_01896_),
    .Y(_01904_));
 sky130_fd_sc_hd__o211ai_4 _12591_ (.A1(_01883_),
    .A2(_01878_),
    .B1(_01882_),
    .C1(_01899_),
    .Y(_01905_));
 sky130_fd_sc_hd__a2bb2oi_1 _12592_ (.A1_N(_01704_),
    .A2_N(_01709_),
    .B1(_01713_),
    .B2(_01694_),
    .Y(_01906_));
 sky130_fd_sc_hd__o21ai_1 _12593_ (.A1(_01696_),
    .A2(_01708_),
    .B1(_01715_),
    .Y(_01907_));
 sky130_fd_sc_hd__a22oi_4 _12594_ (.A1(_01711_),
    .A2(_01715_),
    .B1(_01900_),
    .B2(_01902_),
    .Y(_01908_));
 sky130_fd_sc_hd__o211ai_4 _12595_ (.A1(_01710_),
    .A2(_01714_),
    .B1(_01903_),
    .C1(_01905_),
    .Y(_01909_));
 sky130_fd_sc_hd__a21oi_4 _12596_ (.A1(_01903_),
    .A2(_01905_),
    .B1(_01907_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand3_4 _12597_ (.A(_01900_),
    .B(_01906_),
    .C(_01902_),
    .Y(_01911_));
 sky130_fd_sc_hd__a21o_1 _12598_ (.A1(_01909_),
    .A2(_01911_),
    .B1(_01867_),
    .X(_01913_));
 sky130_fd_sc_hd__o211ai_4 _12599_ (.A1(_01863_),
    .A2(_01864_),
    .B1(_01909_),
    .C1(_01911_),
    .Y(_01914_));
 sky130_fd_sc_hd__nand3_2 _12600_ (.A(_01866_),
    .B(_01909_),
    .C(_01911_),
    .Y(_01915_));
 sky130_fd_sc_hd__inv_2 _12601_ (.A(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__o22ai_4 _12602_ (.A1(_01863_),
    .A2(_01864_),
    .B1(_01908_),
    .B2(_01910_),
    .Y(_01917_));
 sky130_fd_sc_hd__o211ai_2 _12603_ (.A1(_01684_),
    .A2(_01719_),
    .B1(_01841_),
    .C1(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__a22oi_4 _12604_ (.A1(_01723_),
    .A2(_01727_),
    .B1(_01913_),
    .B2(_01914_),
    .Y(_01919_));
 sky130_fd_sc_hd__nand4_2 _12605_ (.A(_01721_),
    .B(_01841_),
    .C(_01915_),
    .D(_01917_),
    .Y(_01920_));
 sky130_fd_sc_hd__a2bb2oi_2 _12606_ (.A1_N(_01720_),
    .A2_N(_01840_),
    .B1(_01915_),
    .B2(_01917_),
    .Y(_01921_));
 sky130_fd_sc_hd__o211ai_4 _12607_ (.A1(_01720_),
    .A2(_01840_),
    .B1(_01913_),
    .C1(_01914_),
    .Y(_01922_));
 sky130_fd_sc_hd__nand2_1 _12608_ (.A(_01838_),
    .B(_01922_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand3_4 _12609_ (.A(_01838_),
    .B(_01920_),
    .C(_01922_),
    .Y(_01925_));
 sky130_fd_sc_hd__inv_2 _12610_ (.A(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__o22ai_4 _12611_ (.A1(_01832_),
    .A2(_01837_),
    .B1(_01919_),
    .B2(_01921_),
    .Y(_01927_));
 sky130_fd_sc_hd__nand2_2 _12612_ (.A(_01790_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__o211a_1 _12613_ (.A1(_01919_),
    .A2(_01924_),
    .B1(_01927_),
    .C1(_01790_),
    .X(_01929_));
 sky130_fd_sc_hd__a2bb2oi_4 _12614_ (.A1_N(_01729_),
    .A2_N(_01789_),
    .B1(_01925_),
    .B2(_01927_),
    .Y(_01930_));
 sky130_fd_sc_hd__a21o_1 _12615_ (.A1(_01925_),
    .A2(_01927_),
    .B1(_01790_),
    .X(_01931_));
 sky130_fd_sc_hd__o211ai_2 _12616_ (.A1(_01926_),
    .A2(_01928_),
    .B1(_01787_),
    .C1(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__inv_2 _12617_ (.A(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__o22ai_2 _12618_ (.A1(_01783_),
    .A2(_01784_),
    .B1(_01929_),
    .B2(_01930_),
    .Y(_01935_));
 sky130_fd_sc_hd__o22ai_4 _12619_ (.A1(_01785_),
    .A2(_01786_),
    .B1(_01929_),
    .B2(_01930_),
    .Y(_01936_));
 sky130_fd_sc_hd__o221ai_4 _12620_ (.A1(_01783_),
    .A2(_01784_),
    .B1(_01926_),
    .B2(_01928_),
    .C1(_01931_),
    .Y(_01937_));
 sky130_fd_sc_hd__nand2_1 _12621_ (.A(_01935_),
    .B(_01766_),
    .Y(_01938_));
 sky130_fd_sc_hd__a22oi_4 _12622_ (.A1(_01738_),
    .A2(_01740_),
    .B1(_01936_),
    .B2(_01937_),
    .Y(_01939_));
 sky130_fd_sc_hd__nand3_2 _12623_ (.A(_01935_),
    .B(_01766_),
    .C(_01932_),
    .Y(_01940_));
 sky130_fd_sc_hd__nand3_4 _12624_ (.A(_01767_),
    .B(_01936_),
    .C(_01937_),
    .Y(_01941_));
 sky130_fd_sc_hd__a2bb2oi_1 _12625_ (.A1_N(_01612_),
    .A2_N(_01617_),
    .B1(_01940_),
    .B2(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__o2bb2ai_2 _12626_ (.A1_N(_01940_),
    .A2_N(_01941_),
    .B1(_01612_),
    .B2(_01617_),
    .Y(_01943_));
 sky130_fd_sc_hd__a31oi_4 _12627_ (.A1(_01767_),
    .A2(_01936_),
    .A3(_01937_),
    .B1(_01622_),
    .Y(_01944_));
 sky130_fd_sc_hd__o2111a_1 _12628_ (.A1(_01385_),
    .A2(_01461_),
    .B1(_01618_),
    .C1(_01940_),
    .D1(_01941_),
    .X(_01946_));
 sky130_fd_sc_hd__o2111ai_4 _12629_ (.A1(_01385_),
    .A2(_01461_),
    .B1(_01618_),
    .C1(_01940_),
    .D1(_01941_),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _12630_ (.A(_01943_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__o2bb2a_1 _12631_ (.A1_N(_01747_),
    .A2_N(_01764_),
    .B1(_01942_),
    .B2(_01946_),
    .X(_01949_));
 sky130_fd_sc_hd__o21ai_1 _12632_ (.A1(_01942_),
    .A2(_01946_),
    .B1(_01765_),
    .Y(_01950_));
 sky130_fd_sc_hd__and4_1 _12633_ (.A(_01747_),
    .B(_01764_),
    .C(_01943_),
    .D(_01947_),
    .X(_01951_));
 sky130_fd_sc_hd__nand4_4 _12634_ (.A(_01747_),
    .B(_01764_),
    .C(_01943_),
    .D(_01947_),
    .Y(_01952_));
 sky130_fd_sc_hd__o211ai_1 _12635_ (.A1(_01600_),
    .A2(_01603_),
    .B1(_01750_),
    .C1(_01751_),
    .Y(_01953_));
 sky130_fd_sc_hd__o21ai_1 _12636_ (.A1(_01949_),
    .A2(_01951_),
    .B1(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__a21oi_1 _12637_ (.A1(_01765_),
    .A2(_01948_),
    .B1(_01754_),
    .Y(_01955_));
 sky130_fd_sc_hd__a31o_1 _12638_ (.A1(_01746_),
    .A2(_01749_),
    .A3(_01948_),
    .B1(_01754_),
    .X(_01957_));
 sky130_fd_sc_hd__nand4b_2 _12639_ (.A_N(_01752_),
    .B(_01950_),
    .C(_01952_),
    .D(_01603_),
    .Y(_01958_));
 sky130_fd_sc_hd__and3_1 _12640_ (.A(_01954_),
    .B(_01957_),
    .C(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__xnor2_1 _12641_ (.A(_01762_),
    .B(_01959_),
    .Y(net72));
 sky130_fd_sc_hd__o22ai_4 _12642_ (.A1(_01916_),
    .A2(_01918_),
    .B1(_01839_),
    .B2(_01921_),
    .Y(_01960_));
 sky130_fd_sc_hd__a21oi_2 _12643_ (.A1(_01838_),
    .A2(_01922_),
    .B1(_01919_),
    .Y(_01961_));
 sky130_fd_sc_hd__o21ai_2 _12644_ (.A1(_01796_),
    .A2(_01798_),
    .B1(_01797_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _12645_ (.A(_01857_),
    .B(_01934_),
    .Y(_01963_));
 sky130_fd_sc_hd__a22oi_4 _12646_ (.A1(net31),
    .A2(net64),
    .B1(net34),
    .B2(net30),
    .Y(_01964_));
 sky130_fd_sc_hd__a22o_1 _12647_ (.A1(net31),
    .A2(net64),
    .B1(net34),
    .B2(net30),
    .X(_01965_));
 sky130_fd_sc_hd__and4_1 _12648_ (.A(net30),
    .B(net31),
    .C(net64),
    .D(net34),
    .X(_01967_));
 sky130_fd_sc_hd__nand4_2 _12649_ (.A(net30),
    .B(net31),
    .C(net64),
    .D(net34),
    .Y(_01968_));
 sky130_fd_sc_hd__o211ai_2 _12650_ (.A1(_01857_),
    .A2(_01934_),
    .B1(_01965_),
    .C1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__o21ai_1 _12651_ (.A1(_01964_),
    .A2(_01967_),
    .B1(_01963_),
    .Y(_01970_));
 sky130_fd_sc_hd__a22o_1 _12652_ (.A1(net29),
    .A2(net35),
    .B1(_01965_),
    .B2(_01968_),
    .X(_01971_));
 sky130_fd_sc_hd__nand4_2 _12653_ (.A(_01965_),
    .B(_01968_),
    .C(net29),
    .D(net35),
    .Y(_01972_));
 sky130_fd_sc_hd__nand3b_4 _12654_ (.A_N(_01962_),
    .B(_01969_),
    .C(_01970_),
    .Y(_01973_));
 sky130_fd_sc_hd__and3_1 _12655_ (.A(_01971_),
    .B(_01972_),
    .C(_01962_),
    .X(_01974_));
 sky130_fd_sc_hd__nand3_4 _12656_ (.A(_01971_),
    .B(_01972_),
    .C(_01962_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _12657_ (.A(net26),
    .B(net38),
    .Y(_01976_));
 sky130_fd_sc_hd__a22oi_4 _12658_ (.A1(net28),
    .A2(net36),
    .B1(net37),
    .B2(net27),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _12659_ (.A(net28),
    .B(net37),
    .Y(_01979_));
 sky130_fd_sc_hd__and4_1 _12660_ (.A(net28),
    .B(net27),
    .C(net36),
    .D(net37),
    .X(_01980_));
 sky130_fd_sc_hd__a211oi_2 _12661_ (.A1(net26),
    .A2(net38),
    .B1(_01978_),
    .C1(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__a211o_1 _12662_ (.A1(net26),
    .A2(net38),
    .B1(_01978_),
    .C1(_01980_),
    .X(_01982_));
 sky130_fd_sc_hd__o211a_1 _12663_ (.A1(_01978_),
    .A2(_01980_),
    .B1(net26),
    .C1(net38),
    .X(_01983_));
 sky130_fd_sc_hd__o211ai_1 _12664_ (.A1(_01978_),
    .A2(_01980_),
    .B1(net26),
    .C1(net38),
    .Y(_01984_));
 sky130_fd_sc_hd__o2bb2a_1 _12665_ (.A1_N(net26),
    .A2_N(net38),
    .B1(_01978_),
    .B2(_01980_),
    .X(_01985_));
 sky130_fd_sc_hd__and4bb_1 _12666_ (.A_N(_01978_),
    .B_N(_01980_),
    .C(net26),
    .D(net38),
    .X(_01986_));
 sky130_fd_sc_hd__o2bb2ai_2 _12667_ (.A1_N(_01973_),
    .A2_N(_01975_),
    .B1(_01981_),
    .B2(_01983_),
    .Y(_01987_));
 sky130_fd_sc_hd__nand4_2 _12668_ (.A(_01973_),
    .B(_01975_),
    .C(_01982_),
    .D(_01984_),
    .Y(_01989_));
 sky130_fd_sc_hd__o2bb2ai_1 _12669_ (.A1_N(_01973_),
    .A2_N(_01975_),
    .B1(_01985_),
    .B2(_01986_),
    .Y(_01990_));
 sky130_fd_sc_hd__o21ai_4 _12670_ (.A1(_01981_),
    .A2(_01983_),
    .B1(_01973_),
    .Y(_01991_));
 sky130_fd_sc_hd__a21oi_1 _12671_ (.A1(_01842_),
    .A2(_01860_),
    .B1(_01858_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand3_4 _12672_ (.A(_01987_),
    .B(_01992_),
    .C(_01989_),
    .Y(_01993_));
 sky130_fd_sc_hd__a22oi_2 _12673_ (.A1(_01859_),
    .A2(_01862_),
    .B1(_01987_),
    .B2(_01989_),
    .Y(_01994_));
 sky130_fd_sc_hd__o221ai_4 _12674_ (.A1(_01858_),
    .A2(_01861_),
    .B1(_01974_),
    .B2(_01991_),
    .C1(_01990_),
    .Y(_01995_));
 sky130_fd_sc_hd__nand2_2 _12675_ (.A(_01806_),
    .B(_01823_),
    .Y(_01996_));
 sky130_fd_sc_hd__a21oi_2 _12676_ (.A1(_01993_),
    .A2(_01995_),
    .B1(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__a21o_1 _12677_ (.A1(_01993_),
    .A2(_01995_),
    .B1(_01996_),
    .X(_01998_));
 sky130_fd_sc_hd__and3_1 _12678_ (.A(_01993_),
    .B(_01995_),
    .C(_01996_),
    .X(_02000_));
 sky130_fd_sc_hd__nand3_1 _12679_ (.A(_01993_),
    .B(_01995_),
    .C(_01996_),
    .Y(_02001_));
 sky130_fd_sc_hd__a22oi_4 _12680_ (.A1(_01806_),
    .A2(_01823_),
    .B1(_01993_),
    .B2(_01995_),
    .Y(_02002_));
 sky130_fd_sc_hd__and4_1 _12681_ (.A(_01806_),
    .B(_01823_),
    .C(_01993_),
    .D(_01995_),
    .X(_02003_));
 sky130_fd_sc_hd__nand2_1 _12682_ (.A(_01998_),
    .B(_02001_),
    .Y(_02004_));
 sky130_fd_sc_hd__o21ai_1 _12683_ (.A1(_01780_),
    .A2(_01966_),
    .B1(_01875_),
    .Y(_02005_));
 sky130_fd_sc_hd__o21ai_2 _12684_ (.A1(_01871_),
    .A2(_01872_),
    .B1(_01875_),
    .Y(_02006_));
 sky130_fd_sc_hd__o21a_1 _12685_ (.A1(_01871_),
    .A2(_01872_),
    .B1(_01875_),
    .X(_02007_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(net55),
    .B(net7),
    .Y(_02008_));
 sky130_fd_sc_hd__a22oi_4 _12687_ (.A1(net44),
    .A2(net8),
    .B1(net9),
    .B2(net33),
    .Y(_02009_));
 sky130_fd_sc_hd__a22o_2 _12688_ (.A1(net44),
    .A2(net8),
    .B1(net9),
    .B2(net33),
    .X(_02011_));
 sky130_fd_sc_hd__and4_1 _12689_ (.A(net33),
    .B(net44),
    .C(net8),
    .D(net9),
    .X(_02012_));
 sky130_fd_sc_hd__nand4_4 _12690_ (.A(net33),
    .B(net44),
    .C(net8),
    .D(net9),
    .Y(_02013_));
 sky130_fd_sc_hd__o211ai_2 _12691_ (.A1(_01780_),
    .A2(_01977_),
    .B1(_02011_),
    .C1(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__o21bai_1 _12692_ (.A1(_02009_),
    .A2(_02012_),
    .B1_N(_02008_),
    .Y(_02015_));
 sky130_fd_sc_hd__o22a_2 _12693_ (.A1(_01780_),
    .A2(_01977_),
    .B1(_02009_),
    .B2(_02012_),
    .X(_02016_));
 sky130_fd_sc_hd__o22ai_4 _12694_ (.A1(_01780_),
    .A2(_01977_),
    .B1(_02009_),
    .B2(_02012_),
    .Y(_02017_));
 sky130_fd_sc_hd__a41o_1 _12695_ (.A1(net33),
    .A2(net44),
    .A3(net8),
    .A4(net9),
    .B1(_02008_),
    .X(_02018_));
 sky130_fd_sc_hd__nand4_2 _12696_ (.A(_02011_),
    .B(_02013_),
    .C(net55),
    .D(net7),
    .Y(_02019_));
 sky130_fd_sc_hd__a22oi_4 _12697_ (.A1(_01873_),
    .A2(_02005_),
    .B1(_02017_),
    .B2(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__nand3_4 _12698_ (.A(_02007_),
    .B(_02014_),
    .C(_02015_),
    .Y(_02022_));
 sky130_fd_sc_hd__o21ai_4 _12699_ (.A1(_02009_),
    .A2(_02018_),
    .B1(_02006_),
    .Y(_02023_));
 sky130_fd_sc_hd__o211a_1 _12700_ (.A1(_02009_),
    .A2(_02018_),
    .B1(_02006_),
    .C1(_02017_),
    .X(_02024_));
 sky130_fd_sc_hd__o211ai_2 _12701_ (.A1(_02009_),
    .A2(_02018_),
    .B1(_02006_),
    .C1(_02017_),
    .Y(_02025_));
 sky130_fd_sc_hd__a22oi_2 _12702_ (.A1(net59),
    .A2(net5),
    .B1(net6),
    .B2(net58),
    .Y(_02026_));
 sky130_fd_sc_hd__a22o_2 _12703_ (.A1(net59),
    .A2(net5),
    .B1(net6),
    .B2(net58),
    .X(_02027_));
 sky130_fd_sc_hd__nand4_4 _12704_ (.A(net58),
    .B(net59),
    .C(net5),
    .D(net6),
    .Y(_02028_));
 sky130_fd_sc_hd__a22oi_4 _12705_ (.A1(net60),
    .A2(net4),
    .B1(_02027_),
    .B2(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__a22o_1 _12706_ (.A1(net60),
    .A2(net4),
    .B1(_02027_),
    .B2(_02028_),
    .X(_02030_));
 sky130_fd_sc_hd__and3_1 _12707_ (.A(_02028_),
    .B(net4),
    .C(net60),
    .X(_02031_));
 sky130_fd_sc_hd__and4_1 _12708_ (.A(_02027_),
    .B(_02028_),
    .C(net60),
    .D(net4),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_1 _12709_ (.A(_02031_),
    .B(_02027_),
    .Y(_02034_));
 sky130_fd_sc_hd__a21oi_2 _12710_ (.A1(_02031_),
    .A2(_02027_),
    .B1(_02029_),
    .Y(_02035_));
 sky130_fd_sc_hd__o21ai_4 _12711_ (.A1(_02020_),
    .A2(_02024_),
    .B1(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__o221ai_4 _12712_ (.A1(_02029_),
    .A2(_02033_),
    .B1(_02016_),
    .B2(_02023_),
    .C1(_02022_),
    .Y(_02037_));
 sky130_fd_sc_hd__o2bb2ai_2 _12713_ (.A1_N(_02022_),
    .A2_N(_02025_),
    .B1(_02029_),
    .B2(_02033_),
    .Y(_02038_));
 sky130_fd_sc_hd__nand3_2 _12714_ (.A(_02025_),
    .B(_02030_),
    .C(_02034_),
    .Y(_02039_));
 sky130_fd_sc_hd__o2111ai_2 _12715_ (.A1(_02016_),
    .A2(_02023_),
    .B1(_02030_),
    .C1(_02034_),
    .D1(_02022_),
    .Y(_02040_));
 sky130_fd_sc_hd__a2bb2oi_4 _12716_ (.A1_N(_01883_),
    .A2_N(_01878_),
    .B1(_01882_),
    .B2(_01899_),
    .Y(_02041_));
 sky130_fd_sc_hd__a21boi_2 _12717_ (.A1(_02038_),
    .A2(_02040_),
    .B1_N(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand3_4 _12718_ (.A(_02036_),
    .B(_02037_),
    .C(_02041_),
    .Y(_02044_));
 sky130_fd_sc_hd__o221a_1 _12719_ (.A1(_02020_),
    .A2(_02039_),
    .B1(_01884_),
    .B2(_01904_),
    .C1(_02038_),
    .X(_02045_));
 sky130_fd_sc_hd__o221ai_4 _12720_ (.A1(_02020_),
    .A2(_02039_),
    .B1(_01884_),
    .B2(_01904_),
    .C1(_02038_),
    .Y(_02046_));
 sky130_fd_sc_hd__o22ai_4 _12721_ (.A1(_01687_),
    .A2(_01888_),
    .B1(_01887_),
    .B2(_01891_),
    .Y(_02047_));
 sky130_fd_sc_hd__and2_1 _12722_ (.A(net63),
    .B(net32),
    .X(_02048_));
 sky130_fd_sc_hd__nand2_2 _12723_ (.A(net62),
    .B(net3),
    .Y(_02049_));
 sky130_fd_sc_hd__and4_1 _12724_ (.A(net61),
    .B(net62),
    .C(net2),
    .D(net3),
    .X(_02050_));
 sky130_fd_sc_hd__nand2_2 _12725_ (.A(net61),
    .B(net3),
    .Y(_02051_));
 sky130_fd_sc_hd__a22o_2 _12726_ (.A1(net62),
    .A2(net2),
    .B1(net3),
    .B2(net61),
    .X(_02052_));
 sky130_fd_sc_hd__o2bb2ai_1 _12727_ (.A1_N(_01847_),
    .A2_N(_02051_),
    .B1(_02049_),
    .B2(_01849_),
    .Y(_02053_));
 sky130_fd_sc_hd__o221ai_4 _12728_ (.A1(_01890_),
    .A2(_01912_),
    .B1(_01849_),
    .B2(_02049_),
    .C1(_02052_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _12729_ (.A(_02053_),
    .B(_02048_),
    .Y(_02056_));
 sky130_fd_sc_hd__o21ai_2 _12730_ (.A1(_01890_),
    .A2(_01912_),
    .B1(_02053_),
    .Y(_02057_));
 sky130_fd_sc_hd__o2111ai_4 _12731_ (.A1(_01849_),
    .A2(_02049_),
    .B1(net63),
    .C1(net32),
    .D1(_02052_),
    .Y(_02058_));
 sky130_fd_sc_hd__a21oi_2 _12732_ (.A1(_02057_),
    .A2(_02058_),
    .B1(_02047_),
    .Y(_02059_));
 sky130_fd_sc_hd__nand3b_4 _12733_ (.A_N(_02047_),
    .B(_02055_),
    .C(_02056_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand3_4 _12734_ (.A(_02057_),
    .B(_02058_),
    .C(_02047_),
    .Y(_02061_));
 sky130_fd_sc_hd__o22a_1 _12735_ (.A1(_01879_),
    .A2(_01890_),
    .B1(_01666_),
    .B2(_01847_),
    .X(_02062_));
 sky130_fd_sc_hd__and3_1 _12736_ (.A(_01851_),
    .B(net63),
    .C(net31),
    .X(_02063_));
 sky130_fd_sc_hd__a31oi_2 _12737_ (.A1(_01851_),
    .A2(net63),
    .A3(net31),
    .B1(_01848_),
    .Y(_02064_));
 sky130_fd_sc_hd__o2bb2a_2 _12738_ (.A1_N(_02060_),
    .A2_N(_02061_),
    .B1(_02062_),
    .B2(_01850_),
    .X(_02066_));
 sky130_fd_sc_hd__o2bb2ai_2 _12739_ (.A1_N(_02060_),
    .A2_N(_02061_),
    .B1(_02062_),
    .B2(_01850_),
    .Y(_02067_));
 sky130_fd_sc_hd__o211a_1 _12740_ (.A1(_01848_),
    .A2(_02063_),
    .B1(_02061_),
    .C1(_02060_),
    .X(_02068_));
 sky130_fd_sc_hd__o211ai_4 _12741_ (.A1(_01848_),
    .A2(_02063_),
    .B1(_02061_),
    .C1(_02060_),
    .Y(_02069_));
 sky130_fd_sc_hd__and3_1 _12742_ (.A(_02060_),
    .B(_02061_),
    .C(_02064_),
    .X(_02070_));
 sky130_fd_sc_hd__o2bb2a_1 _12743_ (.A1_N(_02060_),
    .A2_N(_02061_),
    .B1(_02063_),
    .B2(_01848_),
    .X(_02071_));
 sky130_fd_sc_hd__nand2_2 _12744_ (.A(_02067_),
    .B(_02069_),
    .Y(_02072_));
 sky130_fd_sc_hd__o211ai_4 _12745_ (.A1(_02066_),
    .A2(_02068_),
    .B1(_02044_),
    .C1(_02046_),
    .Y(_02073_));
 sky130_fd_sc_hd__o2bb2ai_2 _12746_ (.A1_N(_02044_),
    .A2_N(_02046_),
    .B1(_02070_),
    .B2(_02071_),
    .Y(_02074_));
 sky130_fd_sc_hd__o2bb2ai_4 _12747_ (.A1_N(_02044_),
    .A2_N(_02046_),
    .B1(_02066_),
    .B2(_02068_),
    .Y(_02075_));
 sky130_fd_sc_hd__o211ai_4 _12748_ (.A1(_02070_),
    .A2(_02071_),
    .B1(_02044_),
    .C1(_02046_),
    .Y(_02077_));
 sky130_fd_sc_hd__a21oi_1 _12749_ (.A1(_01866_),
    .A2(_01911_),
    .B1(_01908_),
    .Y(_02078_));
 sky130_fd_sc_hd__o21ai_4 _12750_ (.A1(_01867_),
    .A2(_01910_),
    .B1(_01909_),
    .Y(_02079_));
 sky130_fd_sc_hd__a21oi_4 _12751_ (.A1(_02075_),
    .A2(_02077_),
    .B1(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__o2111ai_4 _12752_ (.A1(_01910_),
    .A2(_01867_),
    .B1(_01909_),
    .C1(_02073_),
    .D1(_02074_),
    .Y(_02081_));
 sky130_fd_sc_hd__a21oi_4 _12753_ (.A1(_02073_),
    .A2(_02074_),
    .B1(_02078_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand3_2 _12754_ (.A(_02075_),
    .B(_02077_),
    .C(_02079_),
    .Y(_02083_));
 sky130_fd_sc_hd__o21ai_2 _12755_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_02081_),
    .Y(_02084_));
 sky130_fd_sc_hd__o22ai_2 _12756_ (.A1(_01997_),
    .A2(_02000_),
    .B1(_02080_),
    .B2(_02082_),
    .Y(_02085_));
 sky130_fd_sc_hd__o22ai_4 _12757_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_02080_),
    .B2(_02082_),
    .Y(_02086_));
 sky130_fd_sc_hd__o211ai_4 _12758_ (.A1(_01997_),
    .A2(_02000_),
    .B1(_02081_),
    .C1(_02083_),
    .Y(_02088_));
 sky130_fd_sc_hd__o211a_1 _12759_ (.A1(_02082_),
    .A2(_02084_),
    .B1(_01960_),
    .C1(_02085_),
    .X(_02089_));
 sky130_fd_sc_hd__o211ai_4 _12760_ (.A1(_02082_),
    .A2(_02084_),
    .B1(_01960_),
    .C1(_02085_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand3_4 _12761_ (.A(_01961_),
    .B(_02086_),
    .C(_02088_),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2_2 _12762_ (.A(net23),
    .B(net39),
    .Y(_02092_));
 sky130_fd_sc_hd__a22oi_2 _12763_ (.A1(net23),
    .A2(net39),
    .B1(net40),
    .B2(net12),
    .Y(_02093_));
 sky130_fd_sc_hd__a22o_1 _12764_ (.A1(net23),
    .A2(net39),
    .B1(net40),
    .B2(net12),
    .X(_02094_));
 sky130_fd_sc_hd__nand2_1 _12765_ (.A(net23),
    .B(net40),
    .Y(_02095_));
 sky130_fd_sc_hd__and4_2 _12766_ (.A(net23),
    .B(net12),
    .C(net39),
    .D(net40),
    .X(_02096_));
 sky130_fd_sc_hd__nand4_1 _12767_ (.A(net23),
    .B(net12),
    .C(net39),
    .D(net40),
    .Y(_02097_));
 sky130_fd_sc_hd__and4_1 _12768_ (.A(_02094_),
    .B(_02097_),
    .C(net1),
    .D(net41),
    .X(_02099_));
 sky130_fd_sc_hd__nand4_2 _12769_ (.A(_02094_),
    .B(_02097_),
    .C(net1),
    .D(net41),
    .Y(_02100_));
 sky130_fd_sc_hd__o22ai_4 _12770_ (.A1(_01846_),
    .A2(_02010_),
    .B1(_02093_),
    .B2(_02096_),
    .Y(_02101_));
 sky130_fd_sc_hd__o21ai_2 _12771_ (.A1(_01807_),
    .A2(_01809_),
    .B1(_01812_),
    .Y(_02102_));
 sky130_fd_sc_hd__a21oi_2 _12772_ (.A1(_02100_),
    .A2(_02101_),
    .B1(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__a21o_1 _12773_ (.A1(_02100_),
    .A2(_02101_),
    .B1(_02102_),
    .X(_02104_));
 sky130_fd_sc_hd__and3_1 _12774_ (.A(_02100_),
    .B(_02101_),
    .C(_02102_),
    .X(_02105_));
 sky130_fd_sc_hd__nand3_2 _12775_ (.A(_02100_),
    .B(_02101_),
    .C(_02102_),
    .Y(_02106_));
 sky130_fd_sc_hd__nor2_1 _12776_ (.A(_02103_),
    .B(_02105_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand2_1 _12777_ (.A(_02104_),
    .B(_02106_),
    .Y(_02108_));
 sky130_fd_sc_hd__o211ai_2 _12778_ (.A1(_01771_),
    .A2(_01775_),
    .B1(_02104_),
    .C1(_02106_),
    .Y(_02110_));
 sky130_fd_sc_hd__o211ai_2 _12779_ (.A1(_02103_),
    .A2(_02105_),
    .B1(_01772_),
    .C1(_01776_),
    .Y(_02111_));
 sky130_fd_sc_hd__and2_1 _12780_ (.A(_02110_),
    .B(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__nand2_1 _12781_ (.A(_02110_),
    .B(_02111_),
    .Y(_02113_));
 sky130_fd_sc_hd__o211a_1 _12782_ (.A1(_01827_),
    .A2(_01834_),
    .B1(_02110_),
    .C1(_02111_),
    .X(_02114_));
 sky130_fd_sc_hd__o21ai_4 _12783_ (.A1(_01827_),
    .A2(_01834_),
    .B1(_02112_),
    .Y(_02115_));
 sky130_fd_sc_hd__and3_1 _12784_ (.A(_01828_),
    .B(_01836_),
    .C(_02113_),
    .X(_02116_));
 sky130_fd_sc_hd__nand3_2 _12785_ (.A(_01828_),
    .B(_01836_),
    .C(_02113_),
    .Y(_02117_));
 sky130_fd_sc_hd__a22oi_2 _12786_ (.A1(_01614_),
    .A2(_01777_),
    .B1(_02115_),
    .B2(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__a22o_1 _12787_ (.A1(_01614_),
    .A2(_01777_),
    .B1(_02115_),
    .B2(_02117_),
    .X(_02119_));
 sky130_fd_sc_hd__and4_2 _12788_ (.A(_02115_),
    .B(_02117_),
    .C(_01614_),
    .D(_01777_),
    .X(_02121_));
 sky130_fd_sc_hd__nand4_2 _12789_ (.A(_02115_),
    .B(_02117_),
    .C(_01614_),
    .D(_01777_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _12790_ (.A(_02118_),
    .B(_02121_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _12791_ (.A(_02119_),
    .B(_02122_),
    .Y(_02124_));
 sky130_fd_sc_hd__a31oi_2 _12792_ (.A1(_01961_),
    .A2(_02086_),
    .A3(_02088_),
    .B1(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand4_4 _12793_ (.A(_02090_),
    .B(_02091_),
    .C(_02119_),
    .D(_02122_),
    .Y(_02126_));
 sky130_fd_sc_hd__o2bb2ai_4 _12794_ (.A1_N(_02090_),
    .A2_N(_02091_),
    .B1(_02118_),
    .B2(_02121_),
    .Y(_02127_));
 sky130_fd_sc_hd__a31oi_2 _12795_ (.A1(_01927_),
    .A2(_01790_),
    .A3(_01925_),
    .B1(_01787_),
    .Y(_02128_));
 sky130_fd_sc_hd__o22ai_2 _12796_ (.A1(_01926_),
    .A2(_01928_),
    .B1(_01788_),
    .B2(_01930_),
    .Y(_02129_));
 sky130_fd_sc_hd__o2bb2ai_4 _12797_ (.A1_N(_02126_),
    .A2_N(_02127_),
    .B1(_02128_),
    .B2(_01930_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand3_4 _12798_ (.A(_02129_),
    .B(_02127_),
    .C(_02126_),
    .Y(_02132_));
 sky130_fd_sc_hd__o2bb2ai_4 _12799_ (.A1_N(_02130_),
    .A2_N(_02132_),
    .B1(_01768_),
    .B2(_01782_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand3_4 _12800_ (.A(_02130_),
    .B(_02132_),
    .C(_01783_),
    .Y(_02134_));
 sky130_fd_sc_hd__a21bo_1 _12801_ (.A1(_02130_),
    .A2(_02132_),
    .B1_N(_01783_),
    .X(_02135_));
 sky130_fd_sc_hd__o211ai_1 _12802_ (.A1(_01782_),
    .A2(_01768_),
    .B1(_02132_),
    .C1(_02130_),
    .Y(_02136_));
 sky130_fd_sc_hd__o2bb2ai_2 _12803_ (.A1_N(_01621_),
    .A2_N(_01941_),
    .B1(_01938_),
    .B2(_01933_),
    .Y(_02137_));
 sky130_fd_sc_hd__a21oi_1 _12804_ (.A1(_01941_),
    .A2(_01621_),
    .B1(_01939_),
    .Y(_02138_));
 sky130_fd_sc_hd__a21oi_2 _12805_ (.A1(_02133_),
    .A2(_02134_),
    .B1(_02137_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand3_1 _12806_ (.A(_02135_),
    .B(_02136_),
    .C(_02138_),
    .Y(_02140_));
 sky130_fd_sc_hd__o211a_1 _12807_ (.A1(_01939_),
    .A2(_01944_),
    .B1(_02133_),
    .C1(_02134_),
    .X(_02141_));
 sky130_fd_sc_hd__o211ai_4 _12808_ (.A1(_01939_),
    .A2(_01944_),
    .B1(_02133_),
    .C1(_02134_),
    .Y(_02143_));
 sky130_fd_sc_hd__nand2_2 _12809_ (.A(_02140_),
    .B(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__o22ai_2 _12810_ (.A1(_01765_),
    .A2(_01948_),
    .B1(_02139_),
    .B2(_02141_),
    .Y(_02145_));
 sky130_fd_sc_hd__xnor2_1 _12811_ (.A(_01952_),
    .B(_02144_),
    .Y(_02146_));
 sky130_fd_sc_hd__mux2_1 _12812_ (.A0(_02146_),
    .A1(_02145_),
    .S(_01955_),
    .X(_02147_));
 sky130_fd_sc_hd__a21bo_1 _12813_ (.A1(_01763_),
    .A2(_01959_),
    .B1_N(_01958_),
    .X(_02148_));
 sky130_fd_sc_hd__xnor2_1 _12814_ (.A(_02147_),
    .B(_02148_),
    .Y(net73));
 sky130_fd_sc_hd__a32oi_1 _12815_ (.A1(_01600_),
    .A2(_01750_),
    .A3(_01751_),
    .B1(_02140_),
    .B2(_02143_),
    .Y(_02149_));
 sky130_fd_sc_hd__o2bb2ai_1 _12816_ (.A1_N(_01955_),
    .A2_N(_02145_),
    .B1(_02149_),
    .B2(_01958_),
    .Y(_02150_));
 sky130_fd_sc_hd__o211a_1 _12817_ (.A1(_01949_),
    .A2(_01953_),
    .B1(_01954_),
    .C1(_02145_),
    .X(_02151_));
 sky130_fd_sc_hd__nand4_1 _12818_ (.A(_01954_),
    .B(_01957_),
    .C(_01958_),
    .D(_02145_),
    .Y(_02153_));
 sky130_fd_sc_hd__a21oi_1 _12819_ (.A1(_01763_),
    .A2(_02151_),
    .B1(_02150_),
    .Y(_02154_));
 sky130_fd_sc_hd__a31o_1 _12820_ (.A1(_02129_),
    .A2(_02127_),
    .A3(_02126_),
    .B1(_01783_),
    .X(_02155_));
 sky130_fd_sc_hd__a21boi_2 _12821_ (.A1(_02130_),
    .A2(_01783_),
    .B1_N(_02132_),
    .Y(_02156_));
 sky130_fd_sc_hd__a21oi_2 _12822_ (.A1(_02091_),
    .A2(_02123_),
    .B1(_02089_),
    .Y(_02157_));
 sky130_fd_sc_hd__a32oi_4 _12823_ (.A1(_02075_),
    .A2(_02077_),
    .A3(_02079_),
    .B1(_02001_),
    .B2(_01998_),
    .Y(_02158_));
 sky130_fd_sc_hd__o21ai_2 _12824_ (.A1(_02004_),
    .A2(_02080_),
    .B1(_02083_),
    .Y(_02159_));
 sky130_fd_sc_hd__o21a_1 _12825_ (.A1(_01857_),
    .A2(_01934_),
    .B1(_01968_),
    .X(_02160_));
 sky130_fd_sc_hd__a31o_1 _12826_ (.A1(_01965_),
    .A2(net35),
    .A3(net29),
    .B1(_01967_),
    .X(_02161_));
 sky130_fd_sc_hd__nand2_1 _12827_ (.A(net30),
    .B(net35),
    .Y(_02162_));
 sky130_fd_sc_hd__and4_1 _12828_ (.A(net31),
    .B(net32),
    .C(net64),
    .D(net34),
    .X(_02164_));
 sky130_fd_sc_hd__nand4_4 _12829_ (.A(net31),
    .B(net32),
    .C(net64),
    .D(net34),
    .Y(_02165_));
 sky130_fd_sc_hd__a22oi_4 _12830_ (.A1(net32),
    .A2(net64),
    .B1(net34),
    .B2(net31),
    .Y(_02166_));
 sky130_fd_sc_hd__a22o_1 _12831_ (.A1(net32),
    .A2(net64),
    .B1(net34),
    .B2(net31),
    .X(_02167_));
 sky130_fd_sc_hd__a2bb2oi_1 _12832_ (.A1_N(_01868_),
    .A2_N(_01934_),
    .B1(_02165_),
    .B2(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__o21ai_1 _12833_ (.A1(_02164_),
    .A2(_02166_),
    .B1(_02162_),
    .Y(_02169_));
 sky130_fd_sc_hd__nor3_1 _12834_ (.A(_02166_),
    .B(_02162_),
    .C(_02164_),
    .Y(_02170_));
 sky130_fd_sc_hd__nand4_2 _12835_ (.A(_02167_),
    .B(net35),
    .C(net30),
    .D(_02165_),
    .Y(_02171_));
 sky130_fd_sc_hd__and3_1 _12836_ (.A(_02161_),
    .B(_02169_),
    .C(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__nand3_2 _12837_ (.A(_02161_),
    .B(_02169_),
    .C(_02171_),
    .Y(_02173_));
 sky130_fd_sc_hd__o22ai_4 _12838_ (.A1(_01964_),
    .A2(_02160_),
    .B1(_02168_),
    .B2(_02170_),
    .Y(_02175_));
 sky130_fd_sc_hd__nand2_1 _12839_ (.A(net27),
    .B(net38),
    .Y(_02176_));
 sky130_fd_sc_hd__a22oi_2 _12840_ (.A1(net29),
    .A2(net36),
    .B1(net37),
    .B2(net28),
    .Y(_02177_));
 sky130_fd_sc_hd__a22o_1 _12841_ (.A1(net29),
    .A2(net36),
    .B1(net37),
    .B2(net28),
    .X(_02178_));
 sky130_fd_sc_hd__and4_1 _12842_ (.A(net28),
    .B(net29),
    .C(net36),
    .D(net37),
    .X(_02179_));
 sky130_fd_sc_hd__nand4_1 _12843_ (.A(net28),
    .B(net29),
    .C(net36),
    .D(net37),
    .Y(_02180_));
 sky130_fd_sc_hd__and3_1 _12844_ (.A(_02176_),
    .B(_02178_),
    .C(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__o211a_1 _12845_ (.A1(_02177_),
    .A2(_02179_),
    .B1(net27),
    .C1(net38),
    .X(_02182_));
 sky130_fd_sc_hd__o2bb2a_1 _12846_ (.A1_N(net27),
    .A2_N(net38),
    .B1(_02177_),
    .B2(_02179_),
    .X(_02183_));
 sky130_fd_sc_hd__and4_1 _12847_ (.A(_02178_),
    .B(_02180_),
    .C(net27),
    .D(net38),
    .X(_02184_));
 sky130_fd_sc_hd__nor2_1 _12848_ (.A(_02183_),
    .B(_02184_),
    .Y(_02186_));
 sky130_fd_sc_hd__o2bb2ai_1 _12849_ (.A1_N(_02173_),
    .A2_N(_02175_),
    .B1(_02181_),
    .B2(_02182_),
    .Y(_02187_));
 sky130_fd_sc_hd__o211ai_2 _12850_ (.A1(_02183_),
    .A2(_02184_),
    .B1(_02173_),
    .C1(_02175_),
    .Y(_02188_));
 sky130_fd_sc_hd__o2bb2ai_1 _12851_ (.A1_N(_02173_),
    .A2_N(_02175_),
    .B1(_02183_),
    .B2(_02184_),
    .Y(_02189_));
 sky130_fd_sc_hd__o211ai_2 _12852_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_02173_),
    .C1(_02175_),
    .Y(_02190_));
 sky130_fd_sc_hd__o21a_1 _12853_ (.A1(_01850_),
    .A2(_02062_),
    .B1(_02061_),
    .X(_02191_));
 sky130_fd_sc_hd__o21ai_2 _12854_ (.A1(_02064_),
    .A2(_02059_),
    .B1(_02061_),
    .Y(_02192_));
 sky130_fd_sc_hd__o211ai_4 _12855_ (.A1(_02059_),
    .A2(_02191_),
    .B1(_02188_),
    .C1(_02187_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand3_4 _12856_ (.A(_02189_),
    .B(_02190_),
    .C(_02192_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_1 _12857_ (.A(_01975_),
    .B(_01991_),
    .Y(_02195_));
 sky130_fd_sc_hd__a22oi_1 _12858_ (.A1(_01975_),
    .A2(_01991_),
    .B1(_02193_),
    .B2(_02194_),
    .Y(_02197_));
 sky130_fd_sc_hd__a22o_2 _12859_ (.A1(_01975_),
    .A2(_01991_),
    .B1(_02193_),
    .B2(_02194_),
    .X(_02198_));
 sky130_fd_sc_hd__and3b_1 _12860_ (.A_N(_02195_),
    .B(_02194_),
    .C(_02193_),
    .X(_02199_));
 sky130_fd_sc_hd__nand4_4 _12861_ (.A(_01975_),
    .B(_01991_),
    .C(_02193_),
    .D(_02194_),
    .Y(_02200_));
 sky130_fd_sc_hd__a21oi_1 _12862_ (.A1(_02193_),
    .A2(_02194_),
    .B1(_02195_),
    .Y(_02201_));
 sky130_fd_sc_hd__and3_1 _12863_ (.A(_02193_),
    .B(_02194_),
    .C(_02195_),
    .X(_02202_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(_02198_),
    .B(_02200_),
    .Y(_02203_));
 sky130_fd_sc_hd__o21ai_1 _12865_ (.A1(_01780_),
    .A2(_01977_),
    .B1(_02013_),
    .Y(_02204_));
 sky130_fd_sc_hd__o21ai_2 _12866_ (.A1(_02008_),
    .A2(_02009_),
    .B1(_02013_),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _12867_ (.A(net55),
    .B(net8),
    .Y(_02206_));
 sky130_fd_sc_hd__a22oi_4 _12868_ (.A1(net44),
    .A2(net9),
    .B1(net10),
    .B2(net33),
    .Y(_02208_));
 sky130_fd_sc_hd__a22o_1 _12869_ (.A1(net44),
    .A2(net9),
    .B1(net10),
    .B2(net33),
    .X(_02209_));
 sky130_fd_sc_hd__and4_1 _12870_ (.A(net33),
    .B(net44),
    .C(net9),
    .D(net10),
    .X(_02210_));
 sky130_fd_sc_hd__nand4_2 _12871_ (.A(net33),
    .B(net44),
    .C(net9),
    .D(net10),
    .Y(_02211_));
 sky130_fd_sc_hd__o211ai_1 _12872_ (.A1(_01780_),
    .A2(_01988_),
    .B1(_02209_),
    .C1(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__o21bai_1 _12873_ (.A1(_02208_),
    .A2(_02210_),
    .B1_N(_02206_),
    .Y(_02213_));
 sky130_fd_sc_hd__o22a_2 _12874_ (.A1(_01780_),
    .A2(_01988_),
    .B1(_02208_),
    .B2(_02210_),
    .X(_02214_));
 sky130_fd_sc_hd__o22ai_2 _12875_ (.A1(_01780_),
    .A2(_01988_),
    .B1(_02208_),
    .B2(_02210_),
    .Y(_02215_));
 sky130_fd_sc_hd__a41o_1 _12876_ (.A1(net33),
    .A2(net44),
    .A3(net9),
    .A4(net10),
    .B1(_02206_),
    .X(_02216_));
 sky130_fd_sc_hd__nand4_2 _12877_ (.A(_02209_),
    .B(_02211_),
    .C(net55),
    .D(net8),
    .Y(_02217_));
 sky130_fd_sc_hd__a22oi_4 _12878_ (.A1(_02011_),
    .A2(_02204_),
    .B1(_02215_),
    .B2(_02217_),
    .Y(_02219_));
 sky130_fd_sc_hd__nand3b_2 _12879_ (.A_N(_02205_),
    .B(_02212_),
    .C(_02213_),
    .Y(_02220_));
 sky130_fd_sc_hd__o21ai_4 _12880_ (.A1(_02208_),
    .A2(_02216_),
    .B1(_02205_),
    .Y(_02221_));
 sky130_fd_sc_hd__o211a_1 _12881_ (.A1(_02208_),
    .A2(_02216_),
    .B1(_02205_),
    .C1(_02215_),
    .X(_02222_));
 sky130_fd_sc_hd__a22oi_4 _12882_ (.A1(net59),
    .A2(net6),
    .B1(net7),
    .B2(net58),
    .Y(_02223_));
 sky130_fd_sc_hd__a22o_1 _12883_ (.A1(net59),
    .A2(net6),
    .B1(net7),
    .B2(net58),
    .X(_02224_));
 sky130_fd_sc_hd__nand4_2 _12884_ (.A(net58),
    .B(net59),
    .C(net6),
    .D(net7),
    .Y(_02225_));
 sky130_fd_sc_hd__nand2_1 _12885_ (.A(net60),
    .B(net5),
    .Y(_02226_));
 sky130_fd_sc_hd__a22oi_1 _12886_ (.A1(net60),
    .A2(net5),
    .B1(_02224_),
    .B2(_02225_),
    .Y(_02227_));
 sky130_fd_sc_hd__a22o_1 _12887_ (.A1(net60),
    .A2(net5),
    .B1(_02224_),
    .B2(_02225_),
    .X(_02228_));
 sky130_fd_sc_hd__and3_1 _12888_ (.A(_02225_),
    .B(net5),
    .C(net60),
    .X(_02230_));
 sky130_fd_sc_hd__a41o_1 _12889_ (.A1(net58),
    .A2(net59),
    .A3(net6),
    .A4(net7),
    .B1(_02226_),
    .X(_02231_));
 sky130_fd_sc_hd__a21oi_2 _12890_ (.A1(_02230_),
    .A2(_02224_),
    .B1(_02227_),
    .Y(_02232_));
 sky130_fd_sc_hd__o21ai_4 _12891_ (.A1(_02223_),
    .A2(_02231_),
    .B1(_02228_),
    .Y(_02233_));
 sky130_fd_sc_hd__o21ai_1 _12892_ (.A1(_02219_),
    .A2(_02222_),
    .B1(_02232_),
    .Y(_02234_));
 sky130_fd_sc_hd__o211ai_2 _12893_ (.A1(_02214_),
    .A2(_02221_),
    .B1(_02233_),
    .C1(_02220_),
    .Y(_02235_));
 sky130_fd_sc_hd__o21ai_2 _12894_ (.A1(_02219_),
    .A2(_02222_),
    .B1(_02233_),
    .Y(_02236_));
 sky130_fd_sc_hd__o211ai_4 _12895_ (.A1(_02214_),
    .A2(_02221_),
    .B1(_02232_),
    .C1(_02220_),
    .Y(_02237_));
 sky130_fd_sc_hd__a21oi_1 _12896_ (.A1(_02022_),
    .A2(_02035_),
    .B1(_02024_),
    .Y(_02238_));
 sky130_fd_sc_hd__o2bb2ai_2 _12897_ (.A1_N(_02035_),
    .A2_N(_02022_),
    .B1(_02016_),
    .B2(_02023_),
    .Y(_02239_));
 sky130_fd_sc_hd__a21oi_2 _12898_ (.A1(_02236_),
    .A2(_02237_),
    .B1(_02239_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand3_4 _12899_ (.A(_02234_),
    .B(_02238_),
    .C(_02235_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand3_4 _12900_ (.A(_02236_),
    .B(_02237_),
    .C(_02239_),
    .Y(_02243_));
 sky130_fd_sc_hd__o31ai_2 _12901_ (.A1(_01835_),
    .A2(_01945_),
    .A3(_02026_),
    .B1(_02028_),
    .Y(_02244_));
 sky130_fd_sc_hd__o31a_1 _12902_ (.A1(_01835_),
    .A2(_01945_),
    .A3(_02026_),
    .B1(_02028_),
    .X(_02245_));
 sky130_fd_sc_hd__nand2_2 _12903_ (.A(net62),
    .B(net4),
    .Y(_02246_));
 sky130_fd_sc_hd__and4_1 _12904_ (.A(net61),
    .B(net62),
    .C(net3),
    .D(net4),
    .X(_02247_));
 sky130_fd_sc_hd__nand2_1 _12905_ (.A(net61),
    .B(net4),
    .Y(_02248_));
 sky130_fd_sc_hd__a22o_1 _12906_ (.A1(net62),
    .A2(net3),
    .B1(net4),
    .B2(net61),
    .X(_02249_));
 sky130_fd_sc_hd__o2bb2ai_1 _12907_ (.A1_N(_02049_),
    .A2_N(_02248_),
    .B1(_02246_),
    .B2(_02051_),
    .Y(_02250_));
 sky130_fd_sc_hd__o221ai_2 _12908_ (.A1(_01890_),
    .A2(_01901_),
    .B1(_02051_),
    .B2(_02246_),
    .C1(_02249_),
    .Y(_02252_));
 sky130_fd_sc_hd__nand3_1 _12909_ (.A(_02250_),
    .B(net2),
    .C(net63),
    .Y(_02253_));
 sky130_fd_sc_hd__o21ai_1 _12910_ (.A1(_01890_),
    .A2(_01901_),
    .B1(_02250_),
    .Y(_02254_));
 sky130_fd_sc_hd__o2111ai_4 _12911_ (.A1(_02051_),
    .A2(_02246_),
    .B1(net63),
    .C1(net2),
    .D1(_02249_),
    .Y(_02255_));
 sky130_fd_sc_hd__nand3_2 _12912_ (.A(_02245_),
    .B(_02252_),
    .C(_02253_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand3_4 _12913_ (.A(_02254_),
    .B(_02255_),
    .C(_02244_),
    .Y(_02257_));
 sky130_fd_sc_hd__and3_1 _12914_ (.A(_02052_),
    .B(net32),
    .C(net63),
    .X(_02258_));
 sky130_fd_sc_hd__a31o_1 _12915_ (.A1(_02052_),
    .A2(net32),
    .A3(net63),
    .B1(_02050_),
    .X(_02259_));
 sky130_fd_sc_hd__o2bb2a_1 _12916_ (.A1_N(_02048_),
    .A2_N(_02052_),
    .B1(_02049_),
    .B2(_01849_),
    .X(_02260_));
 sky130_fd_sc_hd__a31o_2 _12917_ (.A1(_02245_),
    .A2(_02252_),
    .A3(_02253_),
    .B1(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__and3_1 _12918_ (.A(_02256_),
    .B(_02257_),
    .C(_02259_),
    .X(_02262_));
 sky130_fd_sc_hd__a21oi_1 _12919_ (.A1(_02256_),
    .A2(_02257_),
    .B1(_02259_),
    .Y(_02263_));
 sky130_fd_sc_hd__o2bb2a_1 _12920_ (.A1_N(_02256_),
    .A2_N(_02257_),
    .B1(_02258_),
    .B2(_02050_),
    .X(_02264_));
 sky130_fd_sc_hd__o2bb2ai_4 _12921_ (.A1_N(_02256_),
    .A2_N(_02257_),
    .B1(_02258_),
    .B2(_02050_),
    .Y(_02265_));
 sky130_fd_sc_hd__and3_1 _12922_ (.A(_02256_),
    .B(_02257_),
    .C(_02260_),
    .X(_02266_));
 sky130_fd_sc_hd__nand3_2 _12923_ (.A(_02256_),
    .B(_02257_),
    .C(_02260_),
    .Y(_02267_));
 sky130_fd_sc_hd__nand2_1 _12924_ (.A(_02265_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand4_4 _12925_ (.A(_02242_),
    .B(_02243_),
    .C(_02265_),
    .D(_02267_),
    .Y(_02269_));
 sky130_fd_sc_hd__o2bb2ai_4 _12926_ (.A1_N(_02242_),
    .A2_N(_02243_),
    .B1(_02264_),
    .B2(_02266_),
    .Y(_02270_));
 sky130_fd_sc_hd__o2bb2ai_2 _12927_ (.A1_N(_02242_),
    .A2_N(_02243_),
    .B1(_02262_),
    .B2(_02263_),
    .Y(_02271_));
 sky130_fd_sc_hd__nand3_2 _12928_ (.A(_02242_),
    .B(_02268_),
    .C(_02243_),
    .Y(_02273_));
 sky130_fd_sc_hd__a32oi_4 _12929_ (.A1(_02036_),
    .A2(_02037_),
    .A3(_02041_),
    .B1(_02046_),
    .B2(_02072_),
    .Y(_02274_));
 sky130_fd_sc_hd__a31oi_4 _12930_ (.A1(_02044_),
    .A2(_02067_),
    .A3(_02069_),
    .B1(_02045_),
    .Y(_02275_));
 sky130_fd_sc_hd__a21oi_2 _12931_ (.A1(_02269_),
    .A2(_02270_),
    .B1(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__nand3_1 _12932_ (.A(_02271_),
    .B(_02274_),
    .C(_02273_),
    .Y(_02277_));
 sky130_fd_sc_hd__o2111ai_4 _12933_ (.A1(_02072_),
    .A2(_02042_),
    .B1(_02046_),
    .C1(_02269_),
    .D1(_02270_),
    .Y(_02278_));
 sky130_fd_sc_hd__a32oi_4 _12934_ (.A1(_02269_),
    .A2(_02270_),
    .A3(_02275_),
    .B1(_02200_),
    .B2(_02198_),
    .Y(_02279_));
 sky130_fd_sc_hd__a32oi_4 _12935_ (.A1(_02271_),
    .A2(_02274_),
    .A3(_02273_),
    .B1(_02198_),
    .B2(_02200_),
    .Y(_02280_));
 sky130_fd_sc_hd__o211a_1 _12936_ (.A1(_02197_),
    .A2(_02199_),
    .B1(_02277_),
    .C1(_02278_),
    .X(_02281_));
 sky130_fd_sc_hd__nand2_2 _12937_ (.A(_02280_),
    .B(_02278_),
    .Y(_02282_));
 sky130_fd_sc_hd__a2bb2oi_1 _12938_ (.A1_N(_02201_),
    .A2_N(_02202_),
    .B1(_02277_),
    .B2(_02278_),
    .Y(_02284_));
 sky130_fd_sc_hd__a2bb2o_2 _12939_ (.A1_N(_02201_),
    .A2_N(_02202_),
    .B1(_02277_),
    .B2(_02278_),
    .X(_02285_));
 sky130_fd_sc_hd__a21oi_1 _12940_ (.A1(_02203_),
    .A2(_02278_),
    .B1(_02276_),
    .Y(_02286_));
 sky130_fd_sc_hd__a32o_1 _12941_ (.A1(_02271_),
    .A2(_02274_),
    .A3(_02273_),
    .B1(_02203_),
    .B2(_02278_),
    .X(_02287_));
 sky130_fd_sc_hd__a221oi_2 _12942_ (.A1(_02280_),
    .A2(_02278_),
    .B1(_02084_),
    .B2(_02083_),
    .C1(_02284_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand3_2 _12943_ (.A(_02285_),
    .B(_02159_),
    .C(_02282_),
    .Y(_02289_));
 sky130_fd_sc_hd__a2bb2oi_4 _12944_ (.A1_N(_02080_),
    .A2_N(_02158_),
    .B1(_02282_),
    .B2(_02285_),
    .Y(_02290_));
 sky130_fd_sc_hd__o22ai_2 _12945_ (.A1(_02080_),
    .A2(_02158_),
    .B1(_02281_),
    .B2(_02284_),
    .Y(_02291_));
 sky130_fd_sc_hd__a31o_1 _12946_ (.A1(_02094_),
    .A2(net41),
    .A3(net1),
    .B1(_02096_),
    .X(_02292_));
 sky130_fd_sc_hd__o22ai_4 _12947_ (.A1(_01808_),
    .A2(_01979_),
    .B1(_01976_),
    .B2(_01978_),
    .Y(_02293_));
 sky130_fd_sc_hd__nand2_1 _12948_ (.A(net12),
    .B(net41),
    .Y(_02295_));
 sky130_fd_sc_hd__nand2_2 _12949_ (.A(net26),
    .B(net40),
    .Y(_02296_));
 sky130_fd_sc_hd__nand4_1 _12950_ (.A(net26),
    .B(net23),
    .C(net39),
    .D(net40),
    .Y(_02297_));
 sky130_fd_sc_hd__nand2_2 _12951_ (.A(net26),
    .B(net39),
    .Y(_02298_));
 sky130_fd_sc_hd__a22o_1 _12952_ (.A1(net26),
    .A2(net39),
    .B1(net40),
    .B2(net23),
    .X(_02299_));
 sky130_fd_sc_hd__o2bb2ai_1 _12953_ (.A1_N(_02095_),
    .A2_N(_02298_),
    .B1(_02296_),
    .B2(_02092_),
    .Y(_02300_));
 sky130_fd_sc_hd__o221ai_4 _12954_ (.A1(_01824_),
    .A2(_02010_),
    .B1(_02092_),
    .B2(_02296_),
    .C1(_02299_),
    .Y(_02301_));
 sky130_fd_sc_hd__nand3_1 _12955_ (.A(_02300_),
    .B(net41),
    .C(net12),
    .Y(_02302_));
 sky130_fd_sc_hd__o21ai_1 _12956_ (.A1(_01824_),
    .A2(_02010_),
    .B1(_02300_),
    .Y(_02303_));
 sky130_fd_sc_hd__o2111ai_4 _12957_ (.A1(_02092_),
    .A2(_02296_),
    .B1(net12),
    .C1(net41),
    .D1(_02299_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand3b_4 _12958_ (.A_N(_02293_),
    .B(_02301_),
    .C(_02302_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand3_4 _12959_ (.A(_02303_),
    .B(_02304_),
    .C(_02293_),
    .Y(_02307_));
 sky130_fd_sc_hd__inv_2 _12960_ (.A(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__a21oi_1 _12961_ (.A1(_02306_),
    .A2(_02307_),
    .B1(_02292_),
    .Y(_02309_));
 sky130_fd_sc_hd__a21o_1 _12962_ (.A1(_02306_),
    .A2(_02307_),
    .B1(_02292_),
    .X(_02310_));
 sky130_fd_sc_hd__o21a_1 _12963_ (.A1(_02096_),
    .A2(_02099_),
    .B1(_02306_),
    .X(_02311_));
 sky130_fd_sc_hd__o211a_1 _12964_ (.A1(_02096_),
    .A2(_02099_),
    .B1(_02306_),
    .C1(_02307_),
    .X(_02312_));
 sky130_fd_sc_hd__o211ai_4 _12965_ (.A1(_02096_),
    .A2(_02099_),
    .B1(_02306_),
    .C1(_02307_),
    .Y(_02313_));
 sky130_fd_sc_hd__a21oi_4 _12966_ (.A1(_01772_),
    .A2(_02106_),
    .B1(_02103_),
    .Y(_02314_));
 sky130_fd_sc_hd__a21oi_2 _12967_ (.A1(_02310_),
    .A2(_02313_),
    .B1(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__o21bai_2 _12968_ (.A1(_02309_),
    .A2(_02312_),
    .B1_N(_02314_),
    .Y(_02317_));
 sky130_fd_sc_hd__nand3_2 _12969_ (.A(_02310_),
    .B(_02313_),
    .C(_02314_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _12970_ (.A(net1),
    .B(net42),
    .Y(_02319_));
 sky130_fd_sc_hd__a22o_1 _12971_ (.A1(net1),
    .A2(net42),
    .B1(_02317_),
    .B2(_02318_),
    .X(_02320_));
 sky130_fd_sc_hd__nand4_1 _12972_ (.A(_02317_),
    .B(_02318_),
    .C(net1),
    .D(net42),
    .Y(_02321_));
 sky130_fd_sc_hd__a21o_1 _12973_ (.A1(_02317_),
    .A2(_02318_),
    .B1(_02319_),
    .X(_02322_));
 sky130_fd_sc_hd__nand3_1 _12974_ (.A(_02317_),
    .B(_02318_),
    .C(_02319_),
    .Y(_02323_));
 sky130_fd_sc_hd__o21ai_1 _12975_ (.A1(_01996_),
    .A2(_01994_),
    .B1(_01993_),
    .Y(_02324_));
 sky130_fd_sc_hd__o21a_1 _12976_ (.A1(_01996_),
    .A2(_01994_),
    .B1(_01993_),
    .X(_02325_));
 sky130_fd_sc_hd__nand3_2 _12977_ (.A(_02322_),
    .B(_02323_),
    .C(_02324_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand3_2 _12978_ (.A(_02320_),
    .B(_02321_),
    .C(_02325_),
    .Y(_02328_));
 sky130_fd_sc_hd__inv_2 _12979_ (.A(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__o2bb2a_1 _12980_ (.A1_N(_02326_),
    .A2_N(_02328_),
    .B1(_01776_),
    .B2(_02108_),
    .X(_02330_));
 sky130_fd_sc_hd__o2bb2ai_2 _12981_ (.A1_N(_02326_),
    .A2_N(_02328_),
    .B1(_01776_),
    .B2(_02108_),
    .Y(_02331_));
 sky130_fd_sc_hd__nand4_4 _12982_ (.A(_02326_),
    .B(_02328_),
    .C(_01775_),
    .D(_02107_),
    .Y(_02332_));
 sky130_fd_sc_hd__inv_2 _12983_ (.A(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__nand2_1 _12984_ (.A(_02331_),
    .B(_02332_),
    .Y(_02334_));
 sky130_fd_sc_hd__nand3_2 _12985_ (.A(_02289_),
    .B(_02291_),
    .C(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__o21bai_4 _12986_ (.A1(_02288_),
    .A2(_02290_),
    .B1_N(_02334_),
    .Y(_02336_));
 sky130_fd_sc_hd__o2bb2ai_1 _12987_ (.A1_N(_02289_),
    .A2_N(_02291_),
    .B1(_02330_),
    .B2(_02333_),
    .Y(_02337_));
 sky130_fd_sc_hd__nand3_1 _12988_ (.A(_02289_),
    .B(_02331_),
    .C(_02332_),
    .Y(_02339_));
 sky130_fd_sc_hd__o221ai_4 _12989_ (.A1(_02089_),
    .A2(_02125_),
    .B1(_02290_),
    .B2(_02339_),
    .C1(_02337_),
    .Y(_02340_));
 sky130_fd_sc_hd__and3_1 _12990_ (.A(_02336_),
    .B(_02157_),
    .C(_02335_),
    .X(_02341_));
 sky130_fd_sc_hd__nand3_4 _12991_ (.A(_02336_),
    .B(_02157_),
    .C(_02335_),
    .Y(_02342_));
 sky130_fd_sc_hd__o31a_1 _12992_ (.A1(_01615_),
    .A2(_01774_),
    .A3(_01775_),
    .B1(_02115_),
    .X(_02343_));
 sky130_fd_sc_hd__o311a_1 _12993_ (.A1(_01827_),
    .A2(_01837_),
    .A3(_02112_),
    .B1(_01777_),
    .C1(_01614_),
    .X(_02344_));
 sky130_fd_sc_hd__a31o_1 _12994_ (.A1(_01828_),
    .A2(_01836_),
    .A3(_02113_),
    .B1(_02343_),
    .X(_02345_));
 sky130_fd_sc_hd__o2bb2ai_1 _12995_ (.A1_N(_02340_),
    .A2_N(_02342_),
    .B1(_02344_),
    .B2(_02114_),
    .Y(_02346_));
 sky130_fd_sc_hd__o2111ai_2 _12996_ (.A1(_02116_),
    .A2(_01779_),
    .B1(_02115_),
    .C1(_02340_),
    .D1(_02342_),
    .Y(_02347_));
 sky130_fd_sc_hd__o2bb2ai_2 _12997_ (.A1_N(_02340_),
    .A2_N(_02342_),
    .B1(_02343_),
    .B2(_02116_),
    .Y(_02348_));
 sky130_fd_sc_hd__o211ai_4 _12998_ (.A1(_02114_),
    .A2(_02121_),
    .B1(_02340_),
    .C1(_02342_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2_1 _12999_ (.A(_02348_),
    .B(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__a22oi_1 _13000_ (.A1(_02130_),
    .A2(_02155_),
    .B1(_02348_),
    .B2(_02350_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand3_2 _13001_ (.A(_02156_),
    .B(_02346_),
    .C(_02347_),
    .Y(_02353_));
 sky130_fd_sc_hd__a21oi_1 _13002_ (.A1(_02346_),
    .A2(_02347_),
    .B1(_02156_),
    .Y(_02354_));
 sky130_fd_sc_hd__nand4_4 _13003_ (.A(_02130_),
    .B(_02155_),
    .C(_02348_),
    .D(_02350_),
    .Y(_02355_));
 sky130_fd_sc_hd__nand2_1 _13004_ (.A(_02353_),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__a32oi_4 _13005_ (.A1(_02133_),
    .A2(_02137_),
    .A3(_02134_),
    .B1(_02355_),
    .B2(_02353_),
    .Y(_02357_));
 sky130_fd_sc_hd__nor3_1 _13006_ (.A(_02352_),
    .B(_02354_),
    .C(_02143_),
    .Y(_02358_));
 sky130_fd_sc_hd__nand3_2 _13007_ (.A(_02141_),
    .B(_02353_),
    .C(_02355_),
    .Y(_02359_));
 sky130_fd_sc_hd__o22ai_2 _13008_ (.A1(_01952_),
    .A2(_02144_),
    .B1(_02357_),
    .B2(_02358_),
    .Y(_02361_));
 sky130_fd_sc_hd__nor4_1 _13009_ (.A(_01952_),
    .B(_02139_),
    .C(_02141_),
    .D(_02356_),
    .Y(_02362_));
 sky130_fd_sc_hd__o41a_1 _13010_ (.A1(_01952_),
    .A2(_02139_),
    .A3(_02141_),
    .A4(_02357_),
    .B1(_02361_),
    .X(_02363_));
 sky130_fd_sc_hd__o31ai_4 _13011_ (.A1(_01952_),
    .A2(_02144_),
    .A3(_02357_),
    .B1(_02361_),
    .Y(_02364_));
 sky130_fd_sc_hd__xnor2_1 _13012_ (.A(_02154_),
    .B(_02363_),
    .Y(net74));
 sky130_fd_sc_hd__o311a_1 _13013_ (.A1(_01615_),
    .A2(_02116_),
    .A3(_01778_),
    .B1(_02115_),
    .C1(_02340_),
    .X(_02365_));
 sky130_fd_sc_hd__a32oi_4 _13014_ (.A1(_02157_),
    .A2(_02335_),
    .A3(_02336_),
    .B1(_02340_),
    .B2(_02345_),
    .Y(_02366_));
 sky130_fd_sc_hd__a31o_1 _13015_ (.A1(_02320_),
    .A2(_02321_),
    .A3(_02325_),
    .B1(_02333_),
    .X(_02367_));
 sky130_fd_sc_hd__o21ai_1 _13016_ (.A1(_01835_),
    .A2(_01956_),
    .B1(_02225_),
    .Y(_02368_));
 sky130_fd_sc_hd__o21ai_1 _13017_ (.A1(_02226_),
    .A2(_02223_),
    .B1(_02225_),
    .Y(_02369_));
 sky130_fd_sc_hd__a22o_1 _13018_ (.A1(net62),
    .A2(net4),
    .B1(net5),
    .B2(net61),
    .X(_02371_));
 sky130_fd_sc_hd__nand2_1 _13019_ (.A(net62),
    .B(net5),
    .Y(_02372_));
 sky130_fd_sc_hd__and4_1 _13020_ (.A(net61),
    .B(net62),
    .C(net4),
    .D(net5),
    .X(_02373_));
 sky130_fd_sc_hd__nand4_1 _13021_ (.A(net61),
    .B(net62),
    .C(net4),
    .D(net5),
    .Y(_02374_));
 sky130_fd_sc_hd__a22oi_1 _13022_ (.A1(net63),
    .A2(net3),
    .B1(_02371_),
    .B2(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__o2bb2ai_1 _13023_ (.A1_N(_02371_),
    .A2_N(_02374_),
    .B1(_01890_),
    .B2(_01923_),
    .Y(_02376_));
 sky130_fd_sc_hd__o2111a_1 _13024_ (.A1(_02248_),
    .A2(_02372_),
    .B1(net63),
    .C1(net3),
    .D1(_02371_),
    .X(_02377_));
 sky130_fd_sc_hd__o2111ai_1 _13025_ (.A1(_02248_),
    .A2(_02372_),
    .B1(net63),
    .C1(net3),
    .D1(_02371_),
    .Y(_02378_));
 sky130_fd_sc_hd__o2bb2ai_2 _13026_ (.A1_N(_02224_),
    .A2_N(_02368_),
    .B1(_02375_),
    .B2(_02377_),
    .Y(_02379_));
 sky130_fd_sc_hd__nand3_2 _13027_ (.A(_02369_),
    .B(_02376_),
    .C(_02378_),
    .Y(_02380_));
 sky130_fd_sc_hd__a31o_1 _13028_ (.A1(_02249_),
    .A2(net2),
    .A3(net63),
    .B1(_02247_),
    .X(_02382_));
 sky130_fd_sc_hd__a21o_2 _13029_ (.A1(_02379_),
    .A2(_02380_),
    .B1(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__nand3_4 _13030_ (.A(_02379_),
    .B(_02380_),
    .C(_02382_),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _13031_ (.A(_02383_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__o21ai_2 _13032_ (.A1(_02206_),
    .A2(_02208_),
    .B1(_02211_),
    .Y(_02386_));
 sky130_fd_sc_hd__o21a_1 _13033_ (.A1(_02206_),
    .A2(_02208_),
    .B1(_02211_),
    .X(_02387_));
 sky130_fd_sc_hd__nand2_1 _13034_ (.A(net55),
    .B(net9),
    .Y(_02388_));
 sky130_fd_sc_hd__a22oi_4 _13035_ (.A1(net44),
    .A2(net10),
    .B1(net11),
    .B2(net33),
    .Y(_02389_));
 sky130_fd_sc_hd__a22o_1 _13036_ (.A1(net44),
    .A2(net10),
    .B1(net11),
    .B2(net33),
    .X(_02390_));
 sky130_fd_sc_hd__nand2_1 _13037_ (.A(net44),
    .B(net11),
    .Y(_02391_));
 sky130_fd_sc_hd__and4_1 _13038_ (.A(net33),
    .B(net44),
    .C(net10),
    .D(net11),
    .X(_02393_));
 sky130_fd_sc_hd__nand4_4 _13039_ (.A(net33),
    .B(net44),
    .C(net10),
    .D(net11),
    .Y(_02394_));
 sky130_fd_sc_hd__o211ai_2 _13040_ (.A1(_01780_),
    .A2(_01999_),
    .B1(_02390_),
    .C1(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__o21bai_1 _13041_ (.A1(_02389_),
    .A2(_02393_),
    .B1_N(_02388_),
    .Y(_02396_));
 sky130_fd_sc_hd__o22a_2 _13042_ (.A1(_01780_),
    .A2(_01999_),
    .B1(_02389_),
    .B2(_02393_),
    .X(_02397_));
 sky130_fd_sc_hd__o22ai_2 _13043_ (.A1(_01780_),
    .A2(_01999_),
    .B1(_02389_),
    .B2(_02393_),
    .Y(_02398_));
 sky130_fd_sc_hd__nand4_2 _13044_ (.A(_02390_),
    .B(_02394_),
    .C(net55),
    .D(net9),
    .Y(_02399_));
 sky130_fd_sc_hd__a21oi_1 _13045_ (.A1(_02398_),
    .A2(_02399_),
    .B1(_02386_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand3_4 _13046_ (.A(_02387_),
    .B(_02395_),
    .C(_02396_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand2_2 _13047_ (.A(_02386_),
    .B(_02399_),
    .Y(_02402_));
 sky130_fd_sc_hd__nand3_2 _13048_ (.A(_02398_),
    .B(_02399_),
    .C(_02386_),
    .Y(_02404_));
 sky130_fd_sc_hd__a22oi_4 _13049_ (.A1(net59),
    .A2(net7),
    .B1(net8),
    .B2(net58),
    .Y(_02405_));
 sky130_fd_sc_hd__a22o_1 _13050_ (.A1(net59),
    .A2(net7),
    .B1(net8),
    .B2(net58),
    .X(_02406_));
 sky130_fd_sc_hd__nand4_4 _13051_ (.A(net58),
    .B(net59),
    .C(net7),
    .D(net8),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _13052_ (.A(net60),
    .B(net6),
    .Y(_02408_));
 sky130_fd_sc_hd__a22oi_4 _13053_ (.A1(net60),
    .A2(net6),
    .B1(_02406_),
    .B2(_02407_),
    .Y(_02409_));
 sky130_fd_sc_hd__o2bb2ai_2 _13054_ (.A1_N(_02406_),
    .A2_N(_02407_),
    .B1(_01835_),
    .B2(_01966_),
    .Y(_02410_));
 sky130_fd_sc_hd__a41oi_1 _13055_ (.A1(net58),
    .A2(net59),
    .A3(net7),
    .A4(net8),
    .B1(_02408_),
    .Y(_02411_));
 sky130_fd_sc_hd__a41o_1 _13056_ (.A1(net58),
    .A2(net59),
    .A3(net7),
    .A4(net8),
    .B1(_02408_),
    .X(_02412_));
 sky130_fd_sc_hd__and4_2 _13057_ (.A(_02406_),
    .B(_02407_),
    .C(net60),
    .D(net6),
    .X(_02413_));
 sky130_fd_sc_hd__a21oi_1 _13058_ (.A1(_02406_),
    .A2(_02411_),
    .B1(_02409_),
    .Y(_02415_));
 sky130_fd_sc_hd__o21ai_2 _13059_ (.A1(_02405_),
    .A2(_02412_),
    .B1(_02410_),
    .Y(_02416_));
 sky130_fd_sc_hd__a21o_1 _13060_ (.A1(_02401_),
    .A2(_02404_),
    .B1(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__o221ai_4 _13061_ (.A1(_02409_),
    .A2(_02413_),
    .B1(_02397_),
    .B2(_02402_),
    .C1(_02401_),
    .Y(_02418_));
 sky130_fd_sc_hd__o2bb2ai_4 _13062_ (.A1_N(_02401_),
    .A2_N(_02404_),
    .B1(_02409_),
    .B2(_02413_),
    .Y(_02419_));
 sky130_fd_sc_hd__o2111ai_4 _13063_ (.A1(_02405_),
    .A2(_02412_),
    .B1(_02410_),
    .C1(_02401_),
    .D1(_02404_),
    .Y(_02420_));
 sky130_fd_sc_hd__a21oi_1 _13064_ (.A1(_02220_),
    .A2(_02232_),
    .B1(_02222_),
    .Y(_02421_));
 sky130_fd_sc_hd__o22ai_4 _13065_ (.A1(_02214_),
    .A2(_02221_),
    .B1(_02233_),
    .B2(_02219_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21oi_2 _13066_ (.A1(_02419_),
    .A2(_02420_),
    .B1(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__nand3_4 _13067_ (.A(_02417_),
    .B(_02421_),
    .C(_02418_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand3_4 _13068_ (.A(_02419_),
    .B(_02420_),
    .C(_02422_),
    .Y(_02426_));
 sky130_fd_sc_hd__a21o_1 _13069_ (.A1(_02424_),
    .A2(_02426_),
    .B1(_02385_),
    .X(_02427_));
 sky130_fd_sc_hd__nand3_2 _13070_ (.A(_02385_),
    .B(_02424_),
    .C(_02426_),
    .Y(_02428_));
 sky130_fd_sc_hd__a22o_2 _13071_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_02424_),
    .B2(_02426_),
    .X(_02429_));
 sky130_fd_sc_hd__nand4_4 _13072_ (.A(_02383_),
    .B(_02384_),
    .C(_02424_),
    .D(_02426_),
    .Y(_02430_));
 sky130_fd_sc_hd__a31oi_4 _13073_ (.A1(_02243_),
    .A2(_02265_),
    .A3(_02267_),
    .B1(_02241_),
    .Y(_02431_));
 sky130_fd_sc_hd__a21boi_4 _13074_ (.A1(_02242_),
    .A2(_02268_),
    .B1_N(_02243_),
    .Y(_02432_));
 sky130_fd_sc_hd__and3_1 _13075_ (.A(_02427_),
    .B(_02428_),
    .C(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__nand3_4 _13076_ (.A(_02427_),
    .B(_02428_),
    .C(_02432_),
    .Y(_02434_));
 sky130_fd_sc_hd__a21oi_1 _13077_ (.A1(_02427_),
    .A2(_02428_),
    .B1(_02432_),
    .Y(_02435_));
 sky130_fd_sc_hd__nand3_4 _13078_ (.A(_02429_),
    .B(_02431_),
    .C(_02430_),
    .Y(_02437_));
 sky130_fd_sc_hd__o21a_1 _13079_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_02175_),
    .X(_02438_));
 sky130_fd_sc_hd__a32o_2 _13080_ (.A1(_02161_),
    .A2(_02169_),
    .A3(_02171_),
    .B1(_02175_),
    .B2(_02186_),
    .X(_02439_));
 sky130_fd_sc_hd__nand2_1 _13081_ (.A(_02257_),
    .B(_02261_),
    .Y(_02440_));
 sky130_fd_sc_hd__and2_1 _13082_ (.A(net28),
    .B(net38),
    .X(_02441_));
 sky130_fd_sc_hd__nand2_1 _13083_ (.A(net28),
    .B(net38),
    .Y(_02442_));
 sky130_fd_sc_hd__and4_1 _13084_ (.A(net29),
    .B(net30),
    .C(net36),
    .D(net37),
    .X(_02443_));
 sky130_fd_sc_hd__nand4_1 _13085_ (.A(net29),
    .B(net30),
    .C(net36),
    .D(net37),
    .Y(_02444_));
 sky130_fd_sc_hd__a22oi_2 _13086_ (.A1(net30),
    .A2(net36),
    .B1(net37),
    .B2(net29),
    .Y(_02445_));
 sky130_fd_sc_hd__a22o_1 _13087_ (.A1(net30),
    .A2(net36),
    .B1(net37),
    .B2(net29),
    .X(_02446_));
 sky130_fd_sc_hd__and3_1 _13088_ (.A(_02442_),
    .B(_02444_),
    .C(_02446_),
    .X(_02448_));
 sky130_fd_sc_hd__o211a_1 _13089_ (.A1(_02443_),
    .A2(_02445_),
    .B1(net28),
    .C1(net38),
    .X(_02449_));
 sky130_fd_sc_hd__o2bb2a_1 _13090_ (.A1_N(net28),
    .A2_N(net38),
    .B1(_02443_),
    .B2(_02445_),
    .X(_02450_));
 sky130_fd_sc_hd__and3_1 _13091_ (.A(_02446_),
    .B(_02441_),
    .C(_02444_),
    .X(_02451_));
 sky130_fd_sc_hd__nor2_1 _13092_ (.A(_02448_),
    .B(_02449_),
    .Y(_02452_));
 sky130_fd_sc_hd__o21ai_4 _13093_ (.A1(_02162_),
    .A2(_02166_),
    .B1(_02165_),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_1 _13094_ (.A(net31),
    .B(net35),
    .Y(_02454_));
 sky130_fd_sc_hd__a22oi_4 _13095_ (.A1(net2),
    .A2(net64),
    .B1(net34),
    .B2(net32),
    .Y(_02455_));
 sky130_fd_sc_hd__and4_1 _13096_ (.A(net2),
    .B(net32),
    .C(net64),
    .D(net34),
    .X(_02456_));
 sky130_fd_sc_hd__nand4_1 _13097_ (.A(net2),
    .B(net32),
    .C(net64),
    .D(net34),
    .Y(_02457_));
 sky130_fd_sc_hd__a41o_1 _13098_ (.A1(net2),
    .A2(net32),
    .A3(net64),
    .A4(net34),
    .B1(_02454_),
    .X(_02459_));
 sky130_fd_sc_hd__nand4b_1 _13099_ (.A_N(_02455_),
    .B(_02457_),
    .C(net31),
    .D(net35),
    .Y(_02460_));
 sky130_fd_sc_hd__o22ai_4 _13100_ (.A1(_01879_),
    .A2(_01934_),
    .B1(_02455_),
    .B2(_02456_),
    .Y(_02461_));
 sky130_fd_sc_hd__o211a_1 _13101_ (.A1(_02455_),
    .A2(_02459_),
    .B1(_02453_),
    .C1(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__o211ai_4 _13102_ (.A1(_02455_),
    .A2(_02459_),
    .B1(_02453_),
    .C1(_02461_),
    .Y(_02463_));
 sky130_fd_sc_hd__a21oi_2 _13103_ (.A1(_02460_),
    .A2(_02461_),
    .B1(_02453_),
    .Y(_02464_));
 sky130_fd_sc_hd__a21o_1 _13104_ (.A1(_02460_),
    .A2(_02461_),
    .B1(_02453_),
    .X(_02465_));
 sky130_fd_sc_hd__o22ai_4 _13105_ (.A1(_02448_),
    .A2(_02449_),
    .B1(_02462_),
    .B2(_02464_),
    .Y(_02466_));
 sky130_fd_sc_hd__o211ai_4 _13106_ (.A1(_02450_),
    .A2(_02451_),
    .B1(_02463_),
    .C1(_02465_),
    .Y(_02467_));
 sky130_fd_sc_hd__o211ai_2 _13107_ (.A1(_02448_),
    .A2(_02449_),
    .B1(_02463_),
    .C1(_02465_),
    .Y(_02468_));
 sky130_fd_sc_hd__o21ai_1 _13108_ (.A1(_02462_),
    .A2(_02464_),
    .B1(_02452_),
    .Y(_02470_));
 sky130_fd_sc_hd__a22oi_4 _13109_ (.A1(_02257_),
    .A2(_02261_),
    .B1(_02466_),
    .B2(_02467_),
    .Y(_02471_));
 sky130_fd_sc_hd__a22o_2 _13110_ (.A1(_02257_),
    .A2(_02261_),
    .B1(_02466_),
    .B2(_02467_),
    .X(_02472_));
 sky130_fd_sc_hd__a21oi_4 _13111_ (.A1(_02468_),
    .A2(_02470_),
    .B1(_02440_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand4_4 _13112_ (.A(_02257_),
    .B(_02261_),
    .C(_02466_),
    .D(_02467_),
    .Y(_02474_));
 sky130_fd_sc_hd__nor4_1 _13113_ (.A(_02172_),
    .B(_02438_),
    .C(_02471_),
    .D(_02473_),
    .Y(_02475_));
 sky130_fd_sc_hd__nand3b_1 _13114_ (.A_N(_02439_),
    .B(_02472_),
    .C(_02474_),
    .Y(_02476_));
 sky130_fd_sc_hd__o22a_1 _13115_ (.A1(_02172_),
    .A2(_02438_),
    .B1(_02471_),
    .B2(_02473_),
    .X(_02477_));
 sky130_fd_sc_hd__o21ai_1 _13116_ (.A1(_02471_),
    .A2(_02473_),
    .B1(_02439_),
    .Y(_02478_));
 sky130_fd_sc_hd__and3_1 _13117_ (.A(_02439_),
    .B(_02472_),
    .C(_02474_),
    .X(_02479_));
 sky130_fd_sc_hd__o211ai_4 _13118_ (.A1(_02172_),
    .A2(_02438_),
    .B1(_02472_),
    .C1(_02474_),
    .Y(_02481_));
 sky130_fd_sc_hd__a21oi_1 _13119_ (.A1(_02472_),
    .A2(_02474_),
    .B1(_02439_),
    .Y(_02482_));
 sky130_fd_sc_hd__a21o_2 _13120_ (.A1(_02472_),
    .A2(_02474_),
    .B1(_02439_),
    .X(_02483_));
 sky130_fd_sc_hd__a32oi_2 _13121_ (.A1(_02427_),
    .A2(_02428_),
    .A3(_02432_),
    .B1(_02476_),
    .B2(_02478_),
    .Y(_02484_));
 sky130_fd_sc_hd__nand4_4 _13122_ (.A(_02434_),
    .B(_02437_),
    .C(_02481_),
    .D(_02483_),
    .Y(_02485_));
 sky130_fd_sc_hd__o2bb2ai_4 _13123_ (.A1_N(_02434_),
    .A2_N(_02437_),
    .B1(_02479_),
    .B2(_02482_),
    .Y(_02486_));
 sky130_fd_sc_hd__nand4_1 _13124_ (.A(_02434_),
    .B(_02437_),
    .C(_02476_),
    .D(_02478_),
    .Y(_02487_));
 sky130_fd_sc_hd__o2bb2ai_1 _13125_ (.A1_N(_02434_),
    .A2_N(_02437_),
    .B1(_02475_),
    .B2(_02477_),
    .Y(_02488_));
 sky130_fd_sc_hd__o211ai_4 _13126_ (.A1(_02276_),
    .A2(_02279_),
    .B1(_02485_),
    .C1(_02486_),
    .Y(_02489_));
 sky130_fd_sc_hd__and3_1 _13127_ (.A(_02488_),
    .B(_02286_),
    .C(_02487_),
    .X(_02490_));
 sky130_fd_sc_hd__nand3_2 _13128_ (.A(_02488_),
    .B(_02286_),
    .C(_02487_),
    .Y(_02492_));
 sky130_fd_sc_hd__nand2_1 _13129_ (.A(net12),
    .B(net42),
    .Y(_02493_));
 sky130_fd_sc_hd__and4_2 _13130_ (.A(net12),
    .B(net1),
    .C(net42),
    .D(net43),
    .X(_02494_));
 sky130_fd_sc_hd__a22oi_4 _13131_ (.A1(net12),
    .A2(net42),
    .B1(net43),
    .B2(net1),
    .Y(_02495_));
 sky130_fd_sc_hd__nor2_1 _13132_ (.A(_02494_),
    .B(_02495_),
    .Y(_02496_));
 sky130_fd_sc_hd__or2_1 _13133_ (.A(_02494_),
    .B(_02495_),
    .X(_02497_));
 sky130_fd_sc_hd__nand2_1 _13134_ (.A(_02307_),
    .B(_02313_),
    .Y(_02498_));
 sky130_fd_sc_hd__a22oi_1 _13135_ (.A1(_02295_),
    .A2(_02297_),
    .B1(_02298_),
    .B2(_02095_),
    .Y(_02499_));
 sky130_fd_sc_hd__a22o_1 _13136_ (.A1(_02295_),
    .A2(_02297_),
    .B1(_02298_),
    .B2(_02095_),
    .X(_02500_));
 sky130_fd_sc_hd__nand2_1 _13137_ (.A(_02176_),
    .B(_02180_),
    .Y(_02501_));
 sky130_fd_sc_hd__nor2_1 _13138_ (.A(_02176_),
    .B(_02177_),
    .Y(_02503_));
 sky130_fd_sc_hd__nand2_1 _13139_ (.A(net27),
    .B(net40),
    .Y(_02504_));
 sky130_fd_sc_hd__nand2_2 _13140_ (.A(net27),
    .B(net39),
    .Y(_02505_));
 sky130_fd_sc_hd__and4_1 _13141_ (.A(net27),
    .B(net26),
    .C(net39),
    .D(net40),
    .X(_02506_));
 sky130_fd_sc_hd__nand4_1 _13142_ (.A(net27),
    .B(net26),
    .C(net39),
    .D(net40),
    .Y(_02507_));
 sky130_fd_sc_hd__a22o_2 _13143_ (.A1(net27),
    .A2(net39),
    .B1(net40),
    .B2(net26),
    .X(_02508_));
 sky130_fd_sc_hd__o2111ai_4 _13144_ (.A1(_02298_),
    .A2(_02504_),
    .B1(net23),
    .C1(net41),
    .D1(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__o2bb2ai_2 _13145_ (.A1_N(_02507_),
    .A2_N(_02508_),
    .B1(_01802_),
    .B2(_02010_),
    .Y(_02510_));
 sky130_fd_sc_hd__o211a_1 _13146_ (.A1(_02179_),
    .A2(_02503_),
    .B1(_02509_),
    .C1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__o211ai_2 _13147_ (.A1(_02179_),
    .A2(_02503_),
    .B1(_02509_),
    .C1(_02510_),
    .Y(_02512_));
 sky130_fd_sc_hd__a22oi_4 _13148_ (.A1(_02178_),
    .A2(_02501_),
    .B1(_02509_),
    .B2(_02510_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand3b_2 _13149_ (.A_N(_02514_),
    .B(_02499_),
    .C(_02512_),
    .Y(_02515_));
 sky130_fd_sc_hd__o21ai_4 _13150_ (.A1(_02511_),
    .A2(_02514_),
    .B1(_02500_),
    .Y(_02516_));
 sky130_fd_sc_hd__o211a_1 _13151_ (.A1(_02308_),
    .A2(_02311_),
    .B1(_02515_),
    .C1(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__o211ai_4 _13152_ (.A1(_02308_),
    .A2(_02311_),
    .B1(_02515_),
    .C1(_02516_),
    .Y(_02518_));
 sky130_fd_sc_hd__a21oi_2 _13153_ (.A1(_02515_),
    .A2(_02516_),
    .B1(_02498_),
    .Y(_02519_));
 sky130_fd_sc_hd__a21o_1 _13154_ (.A1(_02515_),
    .A2(_02516_),
    .B1(_02498_),
    .X(_02520_));
 sky130_fd_sc_hd__o21ai_2 _13155_ (.A1(_02517_),
    .A2(_02519_),
    .B1(_02497_),
    .Y(_02521_));
 sky130_fd_sc_hd__nand3_2 _13156_ (.A(_02520_),
    .B(_02496_),
    .C(_02518_),
    .Y(_02522_));
 sky130_fd_sc_hd__o21ai_2 _13157_ (.A1(_02517_),
    .A2(_02519_),
    .B1(_02496_),
    .Y(_02523_));
 sky130_fd_sc_hd__o211ai_4 _13158_ (.A1(_02494_),
    .A2(_02495_),
    .B1(_02518_),
    .C1(_02520_),
    .Y(_02525_));
 sky130_fd_sc_hd__a21bo_1 _13159_ (.A1(_02193_),
    .A2(_02195_),
    .B1_N(_02194_),
    .X(_02526_));
 sky130_fd_sc_hd__a21boi_2 _13160_ (.A1(_02193_),
    .A2(_02195_),
    .B1_N(_02194_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand3_2 _13161_ (.A(_02523_),
    .B(_02525_),
    .C(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand3_4 _13162_ (.A(_02521_),
    .B(_02522_),
    .C(_02526_),
    .Y(_02529_));
 sky130_fd_sc_hd__inv_2 _13163_ (.A(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__a32oi_4 _13164_ (.A1(_02310_),
    .A2(_02313_),
    .A3(_02314_),
    .B1(net42),
    .B2(net1),
    .Y(_02531_));
 sky130_fd_sc_hd__o21a_1 _13165_ (.A1(_02319_),
    .A2(_02315_),
    .B1(_02318_),
    .X(_02532_));
 sky130_fd_sc_hd__a311oi_4 _13166_ (.A1(_02523_),
    .A2(_02525_),
    .A3(_02527_),
    .B1(_02531_),
    .C1(_02315_),
    .Y(_02533_));
 sky130_fd_sc_hd__and3b_1 _13167_ (.A_N(_02532_),
    .B(_02529_),
    .C(_02528_),
    .X(_02534_));
 sky130_fd_sc_hd__nand3b_2 _13168_ (.A_N(_02532_),
    .B(_02529_),
    .C(_02528_),
    .Y(_02536_));
 sky130_fd_sc_hd__o2bb2a_1 _13169_ (.A1_N(_02528_),
    .A2_N(_02529_),
    .B1(_02531_),
    .B2(_02315_),
    .X(_02537_));
 sky130_fd_sc_hd__o2bb2ai_2 _13170_ (.A1_N(_02528_),
    .A2_N(_02529_),
    .B1(_02531_),
    .B2(_02315_),
    .Y(_02538_));
 sky130_fd_sc_hd__a21oi_1 _13171_ (.A1(_02528_),
    .A2(_02529_),
    .B1(_02532_),
    .Y(_02539_));
 sky130_fd_sc_hd__and3_1 _13172_ (.A(_02528_),
    .B(_02529_),
    .C(_02532_),
    .X(_02540_));
 sky130_fd_sc_hd__nand2_1 _13173_ (.A(_02536_),
    .B(_02538_),
    .Y(_02541_));
 sky130_fd_sc_hd__o2bb2ai_2 _13174_ (.A1_N(_02489_),
    .A2_N(_02492_),
    .B1(_02534_),
    .B2(_02537_),
    .Y(_02542_));
 sky130_fd_sc_hd__o21ai_2 _13175_ (.A1(_02539_),
    .A2(_02540_),
    .B1(_02492_),
    .Y(_02543_));
 sky130_fd_sc_hd__nand4_2 _13176_ (.A(_02489_),
    .B(_02492_),
    .C(_02536_),
    .D(_02538_),
    .Y(_02544_));
 sky130_fd_sc_hd__nand3_1 _13177_ (.A(_02489_),
    .B(_02492_),
    .C(_02541_),
    .Y(_02545_));
 sky130_fd_sc_hd__o2bb2ai_1 _13178_ (.A1_N(_02489_),
    .A2_N(_02492_),
    .B1(_02539_),
    .B2(_02540_),
    .Y(_02547_));
 sky130_fd_sc_hd__a32oi_4 _13179_ (.A1(_02285_),
    .A2(_02159_),
    .A3(_02282_),
    .B1(_02331_),
    .B2(_02332_),
    .Y(_02548_));
 sky130_fd_sc_hd__o21ai_2 _13180_ (.A1(_02334_),
    .A2(_02290_),
    .B1(_02289_),
    .Y(_02549_));
 sky130_fd_sc_hd__and3_1 _13181_ (.A(_02549_),
    .B(_02544_),
    .C(_02542_),
    .X(_02550_));
 sky130_fd_sc_hd__nand3_4 _13182_ (.A(_02549_),
    .B(_02544_),
    .C(_02542_),
    .Y(_02551_));
 sky130_fd_sc_hd__o211ai_4 _13183_ (.A1(_02290_),
    .A2(_02548_),
    .B1(_02547_),
    .C1(_02545_),
    .Y(_02552_));
 sky130_fd_sc_hd__o211a_2 _13184_ (.A1(_02329_),
    .A2(_02333_),
    .B1(_02551_),
    .C1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__o211ai_4 _13185_ (.A1(_02329_),
    .A2(_02333_),
    .B1(_02551_),
    .C1(_02552_),
    .Y(_02554_));
 sky130_fd_sc_hd__a21oi_1 _13186_ (.A1(_02551_),
    .A2(_02552_),
    .B1(_02367_),
    .Y(_02555_));
 sky130_fd_sc_hd__a21o_1 _13187_ (.A1(_02551_),
    .A2(_02552_),
    .B1(_02367_),
    .X(_02556_));
 sky130_fd_sc_hd__nand2_1 _13188_ (.A(_02556_),
    .B(_02366_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand3_2 _13189_ (.A(_02556_),
    .B(_02366_),
    .C(_02554_),
    .Y(_02559_));
 sky130_fd_sc_hd__o22ai_4 _13190_ (.A1(_02341_),
    .A2(_02365_),
    .B1(_02553_),
    .B2(_02555_),
    .Y(_02560_));
 sky130_fd_sc_hd__o21ai_2 _13191_ (.A1(_02553_),
    .A2(_02558_),
    .B1(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__o2bb2ai_1 _13192_ (.A1_N(_02559_),
    .A2_N(_02560_),
    .B1(_02156_),
    .B2(_02351_),
    .Y(_02562_));
 sky130_fd_sc_hd__and2_1 _13193_ (.A(_02560_),
    .B(_02354_),
    .X(_02563_));
 sky130_fd_sc_hd__o211ai_1 _13194_ (.A1(_02553_),
    .A2(_02558_),
    .B1(_02560_),
    .C1(_02354_),
    .Y(_02564_));
 sky130_fd_sc_hd__nand2_1 _13195_ (.A(_02562_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__o2bb2ai_1 _13196_ (.A1_N(_02562_),
    .A2_N(_02564_),
    .B1(_02143_),
    .B2(_02356_),
    .Y(_02566_));
 sky130_fd_sc_hd__nor2_1 _13197_ (.A(_02359_),
    .B(_02561_),
    .Y(_02567_));
 sky130_fd_sc_hd__a21oi_1 _13198_ (.A1(_02359_),
    .A2(_02565_),
    .B1(_02567_),
    .Y(_02569_));
 sky130_fd_sc_hd__o21ai_1 _13199_ (.A1(_02359_),
    .A2(_02561_),
    .B1(_02566_),
    .Y(_02570_));
 sky130_fd_sc_hd__o32ai_2 _13200_ (.A1(_01952_),
    .A2(_02144_),
    .A3(_02357_),
    .B1(_02364_),
    .B2(_02154_),
    .Y(_02571_));
 sky130_fd_sc_hd__xor2_1 _13201_ (.A(_02569_),
    .B(_02571_),
    .X(net75));
 sky130_fd_sc_hd__a31o_1 _13202_ (.A1(_02521_),
    .A2(_02522_),
    .A3(_02526_),
    .B1(_02533_),
    .X(_02572_));
 sky130_fd_sc_hd__o21ai_2 _13203_ (.A1(_02500_),
    .A2(_02514_),
    .B1(_02512_),
    .Y(_02573_));
 sky130_fd_sc_hd__and3_1 _13204_ (.A(_02508_),
    .B(net41),
    .C(net23),
    .X(_02574_));
 sky130_fd_sc_hd__a31o_1 _13205_ (.A1(_02508_),
    .A2(net41),
    .A3(net23),
    .B1(_02506_),
    .X(_02575_));
 sky130_fd_sc_hd__a31oi_4 _13206_ (.A1(_02508_),
    .A2(net41),
    .A3(net23),
    .B1(_02506_),
    .Y(_02576_));
 sky130_fd_sc_hd__o21ai_1 _13207_ (.A1(_02442_),
    .A2(_02445_),
    .B1(_02444_),
    .Y(_02577_));
 sky130_fd_sc_hd__a21oi_1 _13208_ (.A1(_02446_),
    .A2(_02441_),
    .B1(_02443_),
    .Y(_02579_));
 sky130_fd_sc_hd__nor2_1 _13209_ (.A(_01791_),
    .B(_02010_),
    .Y(_02580_));
 sky130_fd_sc_hd__nand2_2 _13210_ (.A(net28),
    .B(net40),
    .Y(_02581_));
 sky130_fd_sc_hd__nand2_1 _13211_ (.A(net28),
    .B(net39),
    .Y(_02582_));
 sky130_fd_sc_hd__a22oi_1 _13212_ (.A1(net28),
    .A2(net39),
    .B1(net40),
    .B2(net27),
    .Y(_02583_));
 sky130_fd_sc_hd__a22o_2 _13213_ (.A1(net28),
    .A2(net39),
    .B1(net40),
    .B2(net27),
    .X(_02584_));
 sky130_fd_sc_hd__o2bb2ai_1 _13214_ (.A1_N(_02504_),
    .A2_N(_02582_),
    .B1(_02581_),
    .B2(_02505_),
    .Y(_02585_));
 sky130_fd_sc_hd__o221ai_4 _13215_ (.A1(_01791_),
    .A2(_02010_),
    .B1(_02505_),
    .B2(_02581_),
    .C1(_02584_),
    .Y(_02586_));
 sky130_fd_sc_hd__nand2_1 _13216_ (.A(_02580_),
    .B(_02585_),
    .Y(_02587_));
 sky130_fd_sc_hd__o2111ai_4 _13217_ (.A1(_02505_),
    .A2(_02581_),
    .B1(net26),
    .C1(net41),
    .D1(_02584_),
    .Y(_02588_));
 sky130_fd_sc_hd__o21ai_1 _13218_ (.A1(_01791_),
    .A2(_02010_),
    .B1(_02585_),
    .Y(_02590_));
 sky130_fd_sc_hd__and3_2 _13219_ (.A(_02590_),
    .B(_02577_),
    .C(_02588_),
    .X(_02591_));
 sky130_fd_sc_hd__nand3_2 _13220_ (.A(_02590_),
    .B(_02577_),
    .C(_02588_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21oi_1 _13221_ (.A1(_02588_),
    .A2(_02590_),
    .B1(_02577_),
    .Y(_02593_));
 sky130_fd_sc_hd__nand3_1 _13222_ (.A(_02579_),
    .B(_02586_),
    .C(_02587_),
    .Y(_02594_));
 sky130_fd_sc_hd__a31oi_2 _13223_ (.A1(_02579_),
    .A2(_02586_),
    .A3(_02587_),
    .B1(_02576_),
    .Y(_02595_));
 sky130_fd_sc_hd__a31o_1 _13224_ (.A1(_02579_),
    .A2(_02586_),
    .A3(_02587_),
    .B1(_02576_),
    .X(_02596_));
 sky130_fd_sc_hd__o211a_1 _13225_ (.A1(_02506_),
    .A2(_02574_),
    .B1(_02592_),
    .C1(_02594_),
    .X(_02597_));
 sky130_fd_sc_hd__a21oi_1 _13226_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02575_),
    .Y(_02598_));
 sky130_fd_sc_hd__a21o_1 _13227_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02575_),
    .X(_02599_));
 sky130_fd_sc_hd__o21bai_4 _13228_ (.A1(_02597_),
    .A2(_02598_),
    .B1_N(_02573_),
    .Y(_02601_));
 sky130_fd_sc_hd__o211ai_4 _13229_ (.A1(_02596_),
    .A2(_02591_),
    .B1(_02573_),
    .C1(_02599_),
    .Y(_02602_));
 sky130_fd_sc_hd__and2_1 _13230_ (.A(net1),
    .B(net45),
    .X(_02603_));
 sky130_fd_sc_hd__nand2_1 _13231_ (.A(net23),
    .B(net43),
    .Y(_02604_));
 sky130_fd_sc_hd__nand4_1 _13232_ (.A(net23),
    .B(net12),
    .C(net42),
    .D(net43),
    .Y(_02605_));
 sky130_fd_sc_hd__a22o_1 _13233_ (.A1(net23),
    .A2(net42),
    .B1(net43),
    .B2(net12),
    .X(_02606_));
 sky130_fd_sc_hd__a22o_1 _13234_ (.A1(net1),
    .A2(net45),
    .B1(_02605_),
    .B2(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__o2111ai_1 _13235_ (.A1(_02493_),
    .A2(_02604_),
    .B1(net1),
    .C1(net45),
    .D1(_02606_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_2 _13236_ (.A(_02607_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__or4bb_2 _13237_ (.A(_02609_),
    .B(_02319_),
    .C_N(net43),
    .D_N(net12),
    .X(_02610_));
 sky130_fd_sc_hd__and2_1 _13238_ (.A(_02494_),
    .B(_02609_),
    .X(_02612_));
 sky130_fd_sc_hd__nor2_1 _13239_ (.A(_02494_),
    .B(_02609_),
    .Y(_02613_));
 sky130_fd_sc_hd__xor2_1 _13240_ (.A(_02494_),
    .B(_02609_),
    .X(_02614_));
 sky130_fd_sc_hd__a21bo_1 _13241_ (.A1(_02601_),
    .A2(_02602_),
    .B1_N(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__o211ai_1 _13242_ (.A1(_02612_),
    .A2(_02613_),
    .B1(_02601_),
    .C1(_02602_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand3_1 _13243_ (.A(_02601_),
    .B(_02602_),
    .C(_02614_),
    .Y(_02617_));
 sky130_fd_sc_hd__o2bb2ai_1 _13244_ (.A1_N(_02601_),
    .A2_N(_02602_),
    .B1(_02612_),
    .B2(_02613_),
    .Y(_02618_));
 sky130_fd_sc_hd__nor2_1 _13245_ (.A(_02439_),
    .B(_02471_),
    .Y(_02619_));
 sky130_fd_sc_hd__a21o_1 _13246_ (.A1(_02439_),
    .A2(_02474_),
    .B1(_02471_),
    .X(_02620_));
 sky130_fd_sc_hd__o211ai_4 _13247_ (.A1(_02473_),
    .A2(_02619_),
    .B1(_02618_),
    .C1(_02617_),
    .Y(_02621_));
 sky130_fd_sc_hd__nand3_2 _13248_ (.A(_02615_),
    .B(_02616_),
    .C(_02620_),
    .Y(_02623_));
 sky130_fd_sc_hd__o21a_1 _13249_ (.A1(_02494_),
    .A2(_02495_),
    .B1(_02518_),
    .X(_02624_));
 sky130_fd_sc_hd__o21ai_2 _13250_ (.A1(_02497_),
    .A2(_02519_),
    .B1(_02518_),
    .Y(_02625_));
 sky130_fd_sc_hd__o2bb2ai_2 _13251_ (.A1_N(_02621_),
    .A2_N(_02623_),
    .B1(_02624_),
    .B2(_02519_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand3_2 _13252_ (.A(_02621_),
    .B(_02623_),
    .C(_02625_),
    .Y(_02627_));
 sky130_fd_sc_hd__nand2_1 _13253_ (.A(_02626_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__a32oi_4 _13254_ (.A1(_02419_),
    .A2(_02420_),
    .A3(_02422_),
    .B1(_02384_),
    .B2(_02383_),
    .Y(_02629_));
 sky130_fd_sc_hd__o21ai_2 _13255_ (.A1(_02385_),
    .A2(_02423_),
    .B1(_02426_),
    .Y(_02630_));
 sky130_fd_sc_hd__o21a_1 _13256_ (.A1(_01835_),
    .A2(_01966_),
    .B1(_02407_),
    .X(_02631_));
 sky130_fd_sc_hd__o21ai_2 _13257_ (.A1(_02408_),
    .A2(_02405_),
    .B1(_02407_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand2_1 _13258_ (.A(net63),
    .B(net4),
    .Y(_02634_));
 sky130_fd_sc_hd__nand2_1 _13259_ (.A(net61),
    .B(net6),
    .Y(_02635_));
 sky130_fd_sc_hd__and4_1 _13260_ (.A(net61),
    .B(net62),
    .C(net5),
    .D(net6),
    .X(_02636_));
 sky130_fd_sc_hd__nand4_4 _13261_ (.A(net61),
    .B(net62),
    .C(net5),
    .D(net6),
    .Y(_02637_));
 sky130_fd_sc_hd__a22oi_4 _13262_ (.A1(net62),
    .A2(net5),
    .B1(net6),
    .B2(net61),
    .Y(_02638_));
 sky130_fd_sc_hd__a22o_2 _13263_ (.A1(net62),
    .A2(net5),
    .B1(net6),
    .B2(net61),
    .X(_02639_));
 sky130_fd_sc_hd__o211a_1 _13264_ (.A1(_01890_),
    .A2(_01945_),
    .B1(_02637_),
    .C1(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__a21oi_1 _13265_ (.A1(_02637_),
    .A2(_02639_),
    .B1(_02634_),
    .Y(_02641_));
 sky130_fd_sc_hd__a2bb2oi_4 _13266_ (.A1_N(_01890_),
    .A2_N(_01945_),
    .B1(_02637_),
    .B2(_02639_),
    .Y(_02642_));
 sky130_fd_sc_hd__o21ai_1 _13267_ (.A1(_02636_),
    .A2(_02638_),
    .B1(_02634_),
    .Y(_02643_));
 sky130_fd_sc_hd__nor3_1 _13268_ (.A(_02638_),
    .B(_02634_),
    .C(_02636_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand4_1 _13269_ (.A(_02639_),
    .B(net4),
    .C(net63),
    .D(_02637_),
    .Y(_02646_));
 sky130_fd_sc_hd__o22ai_4 _13270_ (.A1(_02405_),
    .A2(_02631_),
    .B1(_02642_),
    .B2(_02645_),
    .Y(_02647_));
 sky130_fd_sc_hd__nand2_1 _13271_ (.A(_02632_),
    .B(_02646_),
    .Y(_02648_));
 sky130_fd_sc_hd__nand3_2 _13272_ (.A(_02643_),
    .B(_02646_),
    .C(_02632_),
    .Y(_02649_));
 sky130_fd_sc_hd__a31o_4 _13273_ (.A1(_02371_),
    .A2(net3),
    .A3(net63),
    .B1(_02373_),
    .X(_02650_));
 sky130_fd_sc_hd__a21oi_4 _13274_ (.A1(_02647_),
    .A2(_02649_),
    .B1(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__a21o_1 _13275_ (.A1(_02647_),
    .A2(_02649_),
    .B1(_02650_),
    .X(_02652_));
 sky130_fd_sc_hd__o31a_1 _13276_ (.A1(_02632_),
    .A2(_02640_),
    .A3(_02641_),
    .B1(_02650_),
    .X(_02653_));
 sky130_fd_sc_hd__and3_2 _13277_ (.A(_02647_),
    .B(_02649_),
    .C(_02650_),
    .X(_02654_));
 sky130_fd_sc_hd__o211ai_4 _13278_ (.A1(_02642_),
    .A2(_02648_),
    .B1(_02650_),
    .C1(_02647_),
    .Y(_02656_));
 sky130_fd_sc_hd__a21oi_2 _13279_ (.A1(_02653_),
    .A2(_02649_),
    .B1(_02651_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand2_1 _13280_ (.A(_02652_),
    .B(_02656_),
    .Y(_02658_));
 sky130_fd_sc_hd__o21ai_1 _13281_ (.A1(_01780_),
    .A2(_01999_),
    .B1(_02394_),
    .Y(_02659_));
 sky130_fd_sc_hd__o21ai_2 _13282_ (.A1(_02388_),
    .A2(_02389_),
    .B1(_02394_),
    .Y(_02660_));
 sky130_fd_sc_hd__o21a_1 _13283_ (.A1(_02388_),
    .A2(_02389_),
    .B1(_02394_),
    .X(_02661_));
 sky130_fd_sc_hd__nand2_1 _13284_ (.A(net55),
    .B(net10),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_1 _13285_ (.A(net33),
    .B(net13),
    .Y(_02663_));
 sky130_fd_sc_hd__a22oi_4 _13286_ (.A1(net44),
    .A2(net11),
    .B1(net13),
    .B2(net33),
    .Y(_02664_));
 sky130_fd_sc_hd__a22o_2 _13287_ (.A1(net44),
    .A2(net11),
    .B1(net13),
    .B2(net33),
    .X(_02665_));
 sky130_fd_sc_hd__and4_4 _13288_ (.A(net33),
    .B(net44),
    .C(net11),
    .D(net13),
    .X(_02667_));
 sky130_fd_sc_hd__nand4_2 _13289_ (.A(net33),
    .B(net44),
    .C(net11),
    .D(net13),
    .Y(_02668_));
 sky130_fd_sc_hd__o211ai_2 _13290_ (.A1(_01780_),
    .A2(_02021_),
    .B1(_02665_),
    .C1(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__o21bai_1 _13291_ (.A1(_02664_),
    .A2(_02667_),
    .B1_N(_02662_),
    .Y(_02670_));
 sky130_fd_sc_hd__o22a_4 _13292_ (.A1(_01780_),
    .A2(_02021_),
    .B1(_02664_),
    .B2(_02667_),
    .X(_02671_));
 sky130_fd_sc_hd__o22ai_4 _13293_ (.A1(_01780_),
    .A2(_02021_),
    .B1(_02664_),
    .B2(_02667_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand4_4 _13294_ (.A(_02665_),
    .B(_02668_),
    .C(net55),
    .D(net10),
    .Y(_02673_));
 sky130_fd_sc_hd__a22oi_2 _13295_ (.A1(_02390_),
    .A2(_02659_),
    .B1(_02672_),
    .B2(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__nand3_4 _13296_ (.A(_02661_),
    .B(_02669_),
    .C(_02670_),
    .Y(_02675_));
 sky130_fd_sc_hd__nand2_2 _13297_ (.A(_02660_),
    .B(_02673_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand3_1 _13298_ (.A(_02672_),
    .B(_02673_),
    .C(_02660_),
    .Y(_02678_));
 sky130_fd_sc_hd__nand2_1 _13299_ (.A(net60),
    .B(net7),
    .Y(_02679_));
 sky130_fd_sc_hd__a22oi_4 _13300_ (.A1(net59),
    .A2(net8),
    .B1(net9),
    .B2(net58),
    .Y(_02680_));
 sky130_fd_sc_hd__a22o_1 _13301_ (.A1(net59),
    .A2(net8),
    .B1(net9),
    .B2(net58),
    .X(_02681_));
 sky130_fd_sc_hd__and4_1 _13302_ (.A(net58),
    .B(net59),
    .C(net8),
    .D(net9),
    .X(_02682_));
 sky130_fd_sc_hd__nand4_2 _13303_ (.A(net58),
    .B(net59),
    .C(net8),
    .D(net9),
    .Y(_02683_));
 sky130_fd_sc_hd__and3_1 _13304_ (.A(_02679_),
    .B(_02681_),
    .C(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__o211ai_1 _13305_ (.A1(_01835_),
    .A2(_01977_),
    .B1(_02681_),
    .C1(_02683_),
    .Y(_02685_));
 sky130_fd_sc_hd__o211a_1 _13306_ (.A1(_02680_),
    .A2(_02682_),
    .B1(net60),
    .C1(net7),
    .X(_02686_));
 sky130_fd_sc_hd__o21bai_1 _13307_ (.A1(_02680_),
    .A2(_02682_),
    .B1_N(_02679_),
    .Y(_02687_));
 sky130_fd_sc_hd__o22a_1 _13308_ (.A1(_01835_),
    .A2(_01977_),
    .B1(_02680_),
    .B2(_02682_),
    .X(_02689_));
 sky130_fd_sc_hd__o21ai_1 _13309_ (.A1(_02680_),
    .A2(_02682_),
    .B1(_02679_),
    .Y(_02690_));
 sky130_fd_sc_hd__a41o_1 _13310_ (.A1(net58),
    .A2(net59),
    .A3(net8),
    .A4(net9),
    .B1(_02679_),
    .X(_02691_));
 sky130_fd_sc_hd__and4_1 _13311_ (.A(_02681_),
    .B(_02683_),
    .C(net60),
    .D(net7),
    .X(_02692_));
 sky130_fd_sc_hd__o21ai_2 _13312_ (.A1(_02680_),
    .A2(_02691_),
    .B1(_02690_),
    .Y(_02693_));
 sky130_fd_sc_hd__nand2_1 _13313_ (.A(_02685_),
    .B(_02687_),
    .Y(_02694_));
 sky130_fd_sc_hd__a21o_1 _13314_ (.A1(_02675_),
    .A2(_02678_),
    .B1(_02693_),
    .X(_02695_));
 sky130_fd_sc_hd__o221ai_4 _13315_ (.A1(_02689_),
    .A2(_02692_),
    .B1(_02671_),
    .B2(_02676_),
    .C1(_02675_),
    .Y(_02696_));
 sky130_fd_sc_hd__o2bb2ai_2 _13316_ (.A1_N(_02675_),
    .A2_N(_02678_),
    .B1(_02689_),
    .B2(_02692_),
    .Y(_02697_));
 sky130_fd_sc_hd__o221a_4 _13317_ (.A1(_02671_),
    .A2(_02676_),
    .B1(_02684_),
    .B2(_02686_),
    .C1(_02675_),
    .X(_02698_));
 sky130_fd_sc_hd__o221ai_2 _13318_ (.A1(_02671_),
    .A2(_02676_),
    .B1(_02684_),
    .B2(_02686_),
    .C1(_02675_),
    .Y(_02700_));
 sky130_fd_sc_hd__a2bb2oi_2 _13319_ (.A1_N(_02397_),
    .A2_N(_02402_),
    .B1(_02415_),
    .B2(_02401_),
    .Y(_02701_));
 sky130_fd_sc_hd__o22ai_4 _13320_ (.A1(_02397_),
    .A2(_02402_),
    .B1(_02416_),
    .B2(_02400_),
    .Y(_02702_));
 sky130_fd_sc_hd__nand3_4 _13321_ (.A(_02695_),
    .B(_02701_),
    .C(_02696_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand2_2 _13322_ (.A(_02697_),
    .B(_02702_),
    .Y(_02704_));
 sky130_fd_sc_hd__and3_2 _13323_ (.A(_02697_),
    .B(_02700_),
    .C(_02702_),
    .X(_02705_));
 sky130_fd_sc_hd__nand3_2 _13324_ (.A(_02697_),
    .B(_02700_),
    .C(_02702_),
    .Y(_02706_));
 sky130_fd_sc_hd__o221ai_4 _13325_ (.A1(_02651_),
    .A2(_02654_),
    .B1(_02698_),
    .B2(_02704_),
    .C1(_02703_),
    .Y(_02707_));
 sky130_fd_sc_hd__a21o_1 _13326_ (.A1(_02703_),
    .A2(_02706_),
    .B1(_02658_),
    .X(_02708_));
 sky130_fd_sc_hd__a22o_2 _13327_ (.A1(_02652_),
    .A2(_02656_),
    .B1(_02703_),
    .B2(_02706_),
    .X(_02709_));
 sky130_fd_sc_hd__a311oi_4 _13328_ (.A1(_02695_),
    .A2(_02701_),
    .A3(_02696_),
    .B1(_02651_),
    .C1(_02654_),
    .Y(_02711_));
 sky130_fd_sc_hd__nand2_2 _13329_ (.A(_02657_),
    .B(_02703_),
    .Y(_02712_));
 sky130_fd_sc_hd__o2111ai_4 _13330_ (.A1(_02698_),
    .A2(_02704_),
    .B1(_02703_),
    .C1(_02652_),
    .D1(_02656_),
    .Y(_02713_));
 sky130_fd_sc_hd__o211a_2 _13331_ (.A1(_02423_),
    .A2(_02629_),
    .B1(_02707_),
    .C1(_02708_),
    .X(_02714_));
 sky130_fd_sc_hd__o211ai_4 _13332_ (.A1(_02423_),
    .A2(_02629_),
    .B1(_02707_),
    .C1(_02708_),
    .Y(_02715_));
 sky130_fd_sc_hd__o211ai_4 _13333_ (.A1(_02705_),
    .A2(_02712_),
    .B1(_02709_),
    .C1(_02630_),
    .Y(_02716_));
 sky130_fd_sc_hd__a21boi_2 _13334_ (.A1(_02379_),
    .A2(_02382_),
    .B1_N(_02380_),
    .Y(_02717_));
 sky130_fd_sc_hd__nand2_1 _13335_ (.A(net29),
    .B(net38),
    .Y(_02718_));
 sky130_fd_sc_hd__nand4_4 _13336_ (.A(net30),
    .B(net31),
    .C(net36),
    .D(net37),
    .Y(_02719_));
 sky130_fd_sc_hd__a22oi_1 _13337_ (.A1(net31),
    .A2(net36),
    .B1(net37),
    .B2(net30),
    .Y(_02720_));
 sky130_fd_sc_hd__a22o_1 _13338_ (.A1(net31),
    .A2(net36),
    .B1(net37),
    .B2(net30),
    .X(_02722_));
 sky130_fd_sc_hd__and3_1 _13339_ (.A(_02718_),
    .B(_02719_),
    .C(_02722_),
    .X(_02723_));
 sky130_fd_sc_hd__a21oi_1 _13340_ (.A1(_02719_),
    .A2(_02722_),
    .B1(_02718_),
    .Y(_02724_));
 sky130_fd_sc_hd__a22oi_2 _13341_ (.A1(net29),
    .A2(net38),
    .B1(_02719_),
    .B2(_02722_),
    .Y(_02725_));
 sky130_fd_sc_hd__and4_1 _13342_ (.A(_02722_),
    .B(net38),
    .C(net29),
    .D(_02719_),
    .X(_02726_));
 sky130_fd_sc_hd__o21ai_1 _13343_ (.A1(_02454_),
    .A2(_02455_),
    .B1(_02457_),
    .Y(_02727_));
 sky130_fd_sc_hd__o31a_1 _13344_ (.A1(_01879_),
    .A2(_01934_),
    .A3(_02455_),
    .B1(_02457_),
    .X(_02728_));
 sky130_fd_sc_hd__nand2_1 _13345_ (.A(net32),
    .B(net35),
    .Y(_02729_));
 sky130_fd_sc_hd__a22oi_4 _13346_ (.A1(net2),
    .A2(net34),
    .B1(net3),
    .B2(net64),
    .Y(_02730_));
 sky130_fd_sc_hd__a22o_2 _13347_ (.A1(net2),
    .A2(net34),
    .B1(net3),
    .B2(net64),
    .X(_02731_));
 sky130_fd_sc_hd__nand4_4 _13348_ (.A(net2),
    .B(net64),
    .C(net34),
    .D(net3),
    .Y(_02733_));
 sky130_fd_sc_hd__o211ai_2 _13349_ (.A1(_01912_),
    .A2(_01934_),
    .B1(_02731_),
    .C1(_02733_),
    .Y(_02734_));
 sky130_fd_sc_hd__a21o_1 _13350_ (.A1(_02731_),
    .A2(_02733_),
    .B1(_02729_),
    .X(_02735_));
 sky130_fd_sc_hd__a41o_1 _13351_ (.A1(net2),
    .A2(net64),
    .A3(net34),
    .A4(net3),
    .B1(_02729_),
    .X(_02736_));
 sky130_fd_sc_hd__a22o_1 _13352_ (.A1(net32),
    .A2(net35),
    .B1(_02731_),
    .B2(_02733_),
    .X(_02737_));
 sky130_fd_sc_hd__o211ai_4 _13353_ (.A1(_02730_),
    .A2(_02736_),
    .B1(_02727_),
    .C1(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__and3_1 _13354_ (.A(_02728_),
    .B(_02734_),
    .C(_02735_),
    .X(_02739_));
 sky130_fd_sc_hd__nand3_1 _13355_ (.A(_02728_),
    .B(_02734_),
    .C(_02735_),
    .Y(_02740_));
 sky130_fd_sc_hd__a2bb2o_1 _13356_ (.A1_N(_02723_),
    .A2_N(_02724_),
    .B1(_02738_),
    .B2(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__o211ai_1 _13357_ (.A1(_02725_),
    .A2(_02726_),
    .B1(_02738_),
    .C1(_02740_),
    .Y(_02742_));
 sky130_fd_sc_hd__a311o_2 _13358_ (.A1(_02728_),
    .A2(_02734_),
    .A3(_02735_),
    .B1(_02726_),
    .C1(_02725_),
    .X(_02744_));
 sky130_fd_sc_hd__o211ai_2 _13359_ (.A1(_02723_),
    .A2(_02724_),
    .B1(_02738_),
    .C1(_02740_),
    .Y(_02745_));
 sky130_fd_sc_hd__a2bb2o_1 _13360_ (.A1_N(_02725_),
    .A2_N(_02726_),
    .B1(_02738_),
    .B2(_02740_),
    .X(_02746_));
 sky130_fd_sc_hd__nand3_2 _13361_ (.A(_02741_),
    .B(_02742_),
    .C(_02717_),
    .Y(_02747_));
 sky130_fd_sc_hd__nand3b_4 _13362_ (.A_N(_02717_),
    .B(_02745_),
    .C(_02746_),
    .Y(_02748_));
 sky130_fd_sc_hd__o31a_1 _13363_ (.A1(_02450_),
    .A2(_02451_),
    .A3(_02464_),
    .B1(_02463_),
    .X(_02749_));
 sky130_fd_sc_hd__o21ai_2 _13364_ (.A1(_02452_),
    .A2(_02464_),
    .B1(_02463_),
    .Y(_02750_));
 sky130_fd_sc_hd__a21oi_1 _13365_ (.A1(_02747_),
    .A2(_02748_),
    .B1(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__a21o_1 _13366_ (.A1(_02747_),
    .A2(_02748_),
    .B1(_02750_),
    .X(_02752_));
 sky130_fd_sc_hd__and3_1 _13367_ (.A(_02747_),
    .B(_02748_),
    .C(_02750_),
    .X(_02753_));
 sky130_fd_sc_hd__nand3_2 _13368_ (.A(_02747_),
    .B(_02748_),
    .C(_02750_),
    .Y(_02755_));
 sky130_fd_sc_hd__and3_1 _13369_ (.A(_02747_),
    .B(_02748_),
    .C(_02749_),
    .X(_02756_));
 sky130_fd_sc_hd__a21oi_1 _13370_ (.A1(_02747_),
    .A2(_02748_),
    .B1(_02749_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand3_1 _13371_ (.A(_02715_),
    .B(_02752_),
    .C(_02755_),
    .Y(_02758_));
 sky130_fd_sc_hd__nand4_4 _13372_ (.A(_02715_),
    .B(_02716_),
    .C(_02752_),
    .D(_02755_),
    .Y(_02759_));
 sky130_fd_sc_hd__o2bb2ai_2 _13373_ (.A1_N(_02715_),
    .A2_N(_02716_),
    .B1(_02751_),
    .B2(_02753_),
    .Y(_02760_));
 sky130_fd_sc_hd__o211ai_2 _13374_ (.A1(_02751_),
    .A2(_02753_),
    .B1(_02715_),
    .C1(_02716_),
    .Y(_02761_));
 sky130_fd_sc_hd__o2bb2ai_1 _13375_ (.A1_N(_02715_),
    .A2_N(_02716_),
    .B1(_02756_),
    .B2(_02757_),
    .Y(_02762_));
 sky130_fd_sc_hd__a32oi_4 _13376_ (.A1(_02429_),
    .A2(_02431_),
    .A3(_02430_),
    .B1(_02483_),
    .B2(_02481_),
    .Y(_02763_));
 sky130_fd_sc_hd__a31o_1 _13377_ (.A1(_02434_),
    .A2(_02481_),
    .A3(_02483_),
    .B1(_02435_),
    .X(_02764_));
 sky130_fd_sc_hd__o211a_1 _13378_ (.A1(_02433_),
    .A2(_02763_),
    .B1(_02762_),
    .C1(_02761_),
    .X(_02766_));
 sky130_fd_sc_hd__o211ai_2 _13379_ (.A1(_02433_),
    .A2(_02763_),
    .B1(_02762_),
    .C1(_02761_),
    .Y(_02767_));
 sky130_fd_sc_hd__o211ai_2 _13380_ (.A1(_02435_),
    .A2(_02484_),
    .B1(_02759_),
    .C1(_02760_),
    .Y(_02768_));
 sky130_fd_sc_hd__a21o_1 _13381_ (.A1(_02767_),
    .A2(_02768_),
    .B1(_02628_),
    .X(_02769_));
 sky130_fd_sc_hd__nand3_2 _13382_ (.A(_02628_),
    .B(_02767_),
    .C(_02768_),
    .Y(_02770_));
 sky130_fd_sc_hd__a32oi_4 _13383_ (.A1(_02287_),
    .A2(_02485_),
    .A3(_02486_),
    .B1(_02536_),
    .B2(_02538_),
    .Y(_02771_));
 sky130_fd_sc_hd__a22oi_4 _13384_ (.A1(_02489_),
    .A2(_02543_),
    .B1(_02769_),
    .B2(_02770_),
    .Y(_02772_));
 sky130_fd_sc_hd__a22o_1 _13385_ (.A1(_02489_),
    .A2(_02543_),
    .B1(_02769_),
    .B2(_02770_),
    .X(_02773_));
 sky130_fd_sc_hd__o211a_1 _13386_ (.A1(_02490_),
    .A2(_02771_),
    .B1(_02770_),
    .C1(_02769_),
    .X(_02774_));
 sky130_fd_sc_hd__o211ai_2 _13387_ (.A1(_02490_),
    .A2(_02771_),
    .B1(_02770_),
    .C1(_02769_),
    .Y(_02775_));
 sky130_fd_sc_hd__o22ai_2 _13388_ (.A1(_02530_),
    .A2(_02533_),
    .B1(_02772_),
    .B2(_02774_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand3b_1 _13389_ (.A_N(_02572_),
    .B(_02773_),
    .C(_02775_),
    .Y(_02778_));
 sky130_fd_sc_hd__o21ai_1 _13390_ (.A1(_02530_),
    .A2(_02533_),
    .B1(_02775_),
    .Y(_02779_));
 sky130_fd_sc_hd__o21bai_1 _13391_ (.A1(_02772_),
    .A2(_02774_),
    .B1_N(_02572_),
    .Y(_02780_));
 sky130_fd_sc_hd__o221ai_4 _13392_ (.A1(_02772_),
    .A2(_02779_),
    .B1(_02550_),
    .B2(_02553_),
    .C1(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand4_4 _13393_ (.A(_02551_),
    .B(_02554_),
    .C(_02777_),
    .D(_02778_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand3b_2 _13394_ (.A_N(_02559_),
    .B(_02781_),
    .C(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__o2bb2ai_1 _13395_ (.A1_N(_02781_),
    .A2_N(_02782_),
    .B1(_02553_),
    .B2(_02558_),
    .Y(_02784_));
 sky130_fd_sc_hd__o2bb2ai_1 _13396_ (.A1_N(_02783_),
    .A2_N(_02784_),
    .B1(_02355_),
    .B2(_02561_),
    .Y(_02785_));
 sky130_fd_sc_hd__and4_1 _13397_ (.A(_02563_),
    .B(_02781_),
    .C(_02782_),
    .D(_02559_),
    .X(_02786_));
 sky130_fd_sc_hd__nand4_2 _13398_ (.A(_02563_),
    .B(_02781_),
    .C(_02782_),
    .D(_02559_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _13399_ (.A(_02785_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__o211ai_2 _13400_ (.A1(_02359_),
    .A2(_02561_),
    .B1(_02566_),
    .C1(_02150_),
    .Y(_02790_));
 sky130_fd_sc_hd__a21oi_1 _13401_ (.A1(_02566_),
    .A2(_02362_),
    .B1(_02567_),
    .Y(_02791_));
 sky130_fd_sc_hd__o21ai_4 _13402_ (.A1(_02364_),
    .A2(_02790_),
    .B1(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__nor3_2 _13403_ (.A(_02153_),
    .B(_02364_),
    .C(_02570_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand3_2 _13404_ (.A(_02151_),
    .B(_02363_),
    .C(_02569_),
    .Y(_02794_));
 sky130_fd_sc_hd__a21oi_1 _13405_ (.A1(_01763_),
    .A2(_02793_),
    .B1(_02792_),
    .Y(_02795_));
 sky130_fd_sc_hd__nor2_1 _13406_ (.A(_02789_),
    .B(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__a221oi_1 _13407_ (.A1(_02785_),
    .A2(_02788_),
    .B1(_01763_),
    .B2(_02793_),
    .C1(_02792_),
    .Y(_02797_));
 sky130_fd_sc_hd__nor2_1 _13408_ (.A(_02796_),
    .B(_02797_),
    .Y(net77));
 sky130_fd_sc_hd__a32oi_4 _13409_ (.A1(_02764_),
    .A2(_02760_),
    .A3(_02759_),
    .B1(_02626_),
    .B2(_02627_),
    .Y(_02799_));
 sky130_fd_sc_hd__o21ai_1 _13410_ (.A1(_02628_),
    .A2(_02766_),
    .B1(_02768_),
    .Y(_02800_));
 sky130_fd_sc_hd__a32oi_4 _13411_ (.A1(_02630_),
    .A2(_02709_),
    .A3(_02713_),
    .B1(_02752_),
    .B2(_02755_),
    .Y(_02801_));
 sky130_fd_sc_hd__nand2_1 _13412_ (.A(_02716_),
    .B(_02758_),
    .Y(_02802_));
 sky130_fd_sc_hd__a21boi_2 _13413_ (.A1(_02647_),
    .A2(_02650_),
    .B1_N(_02649_),
    .Y(_02803_));
 sky130_fd_sc_hd__o2bb2ai_2 _13414_ (.A1_N(_02650_),
    .A2_N(_02647_),
    .B1(_02642_),
    .B2(_02648_),
    .Y(_02804_));
 sky130_fd_sc_hd__o21ai_1 _13415_ (.A1(_01912_),
    .A2(_01934_),
    .B1(_02733_),
    .Y(_02805_));
 sky130_fd_sc_hd__o21ai_2 _13416_ (.A1(_02729_),
    .A2(_02730_),
    .B1(_02733_),
    .Y(_02806_));
 sky130_fd_sc_hd__nand2_2 _13417_ (.A(net2),
    .B(net35),
    .Y(_02807_));
 sky130_fd_sc_hd__and4_1 _13418_ (.A(net64),
    .B(net34),
    .C(net3),
    .D(net4),
    .X(_02809_));
 sky130_fd_sc_hd__nand4_4 _13419_ (.A(net64),
    .B(net34),
    .C(net3),
    .D(net4),
    .Y(_02810_));
 sky130_fd_sc_hd__a22oi_4 _13420_ (.A1(net34),
    .A2(net3),
    .B1(net4),
    .B2(net64),
    .Y(_02811_));
 sky130_fd_sc_hd__a22o_1 _13421_ (.A1(net34),
    .A2(net3),
    .B1(net4),
    .B2(net64),
    .X(_02812_));
 sky130_fd_sc_hd__a2bb2oi_2 _13422_ (.A1_N(_01901_),
    .A2_N(_01934_),
    .B1(_02810_),
    .B2(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__o21ai_2 _13423_ (.A1(_02809_),
    .A2(_02811_),
    .B1(_02807_),
    .Y(_02814_));
 sky130_fd_sc_hd__nor3_2 _13424_ (.A(_02811_),
    .B(_02807_),
    .C(_02809_),
    .Y(_02815_));
 sky130_fd_sc_hd__nand4_4 _13425_ (.A(_02812_),
    .B(net35),
    .C(net2),
    .D(_02810_),
    .Y(_02816_));
 sky130_fd_sc_hd__o221a_1 _13426_ (.A1(_02729_),
    .A2(_02730_),
    .B1(_02813_),
    .B2(_02815_),
    .C1(_02733_),
    .X(_02817_));
 sky130_fd_sc_hd__o2bb2ai_4 _13427_ (.A1_N(_02731_),
    .A2_N(_02805_),
    .B1(_02813_),
    .B2(_02815_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand3_2 _13428_ (.A(_02814_),
    .B(_02816_),
    .C(_02806_),
    .Y(_02820_));
 sky130_fd_sc_hd__nand2_1 _13429_ (.A(net30),
    .B(net38),
    .Y(_02821_));
 sky130_fd_sc_hd__a22oi_4 _13430_ (.A1(net32),
    .A2(net36),
    .B1(net37),
    .B2(net31),
    .Y(_02822_));
 sky130_fd_sc_hd__and4_1 _13431_ (.A(net31),
    .B(net32),
    .C(net36),
    .D(net37),
    .X(_02823_));
 sky130_fd_sc_hd__nand4_1 _13432_ (.A(net31),
    .B(net32),
    .C(net36),
    .D(net37),
    .Y(_02824_));
 sky130_fd_sc_hd__a211oi_2 _13433_ (.A1(net30),
    .A2(net38),
    .B1(_02822_),
    .C1(_02823_),
    .Y(_02825_));
 sky130_fd_sc_hd__a211o_1 _13434_ (.A1(net30),
    .A2(net38),
    .B1(_02822_),
    .C1(_02823_),
    .X(_02826_));
 sky130_fd_sc_hd__o211a_1 _13435_ (.A1(_02822_),
    .A2(_02823_),
    .B1(net30),
    .C1(net38),
    .X(_02827_));
 sky130_fd_sc_hd__o211ai_2 _13436_ (.A1(_02822_),
    .A2(_02823_),
    .B1(net30),
    .C1(net38),
    .Y(_02828_));
 sky130_fd_sc_hd__o2bb2a_1 _13437_ (.A1_N(net30),
    .A2_N(net38),
    .B1(_02822_),
    .B2(_02823_),
    .X(_02829_));
 sky130_fd_sc_hd__and4b_1 _13438_ (.A_N(_02822_),
    .B(_02824_),
    .C(net30),
    .D(net38),
    .X(_02831_));
 sky130_fd_sc_hd__nand2_1 _13439_ (.A(_02826_),
    .B(_02828_),
    .Y(_02832_));
 sky130_fd_sc_hd__o21ai_2 _13440_ (.A1(_02825_),
    .A2(_02827_),
    .B1(_02820_),
    .Y(_02833_));
 sky130_fd_sc_hd__o2bb2ai_2 _13441_ (.A1_N(_02818_),
    .A2_N(_02820_),
    .B1(_02829_),
    .B2(_02831_),
    .Y(_02834_));
 sky130_fd_sc_hd__nand4_2 _13442_ (.A(_02818_),
    .B(_02820_),
    .C(_02826_),
    .D(_02828_),
    .Y(_02835_));
 sky130_fd_sc_hd__o2bb2ai_2 _13443_ (.A1_N(_02818_),
    .A2_N(_02820_),
    .B1(_02825_),
    .B2(_02827_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand3_4 _13444_ (.A(_02836_),
    .B(_02803_),
    .C(_02835_),
    .Y(_02837_));
 sky130_fd_sc_hd__o211a_2 _13445_ (.A1(_02833_),
    .A2(_02817_),
    .B1(_02804_),
    .C1(_02834_),
    .X(_02838_));
 sky130_fd_sc_hd__o211ai_4 _13446_ (.A1(_02833_),
    .A2(_02817_),
    .B1(_02804_),
    .C1(_02834_),
    .Y(_02839_));
 sky130_fd_sc_hd__o31a_1 _13447_ (.A1(_02725_),
    .A2(_02726_),
    .A3(_02739_),
    .B1(_02738_),
    .X(_02840_));
 sky130_fd_sc_hd__nand2_2 _13448_ (.A(_02738_),
    .B(_02744_),
    .Y(_02842_));
 sky130_fd_sc_hd__a21oi_1 _13449_ (.A1(_02837_),
    .A2(_02839_),
    .B1(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__a21o_1 _13450_ (.A1(_02837_),
    .A2(_02839_),
    .B1(_02842_),
    .X(_02844_));
 sky130_fd_sc_hd__a32o_1 _13451_ (.A1(_02836_),
    .A2(_02803_),
    .A3(_02835_),
    .B1(_02744_),
    .B2(_02738_),
    .X(_02845_));
 sky130_fd_sc_hd__and3_1 _13452_ (.A(_02837_),
    .B(_02839_),
    .C(_02842_),
    .X(_02846_));
 sky130_fd_sc_hd__a21oi_1 _13453_ (.A1(_02837_),
    .A2(_02839_),
    .B1(_02840_),
    .Y(_02847_));
 sky130_fd_sc_hd__a22o_1 _13454_ (.A1(_02738_),
    .A2(_02744_),
    .B1(_02837_),
    .B2(_02839_),
    .X(_02848_));
 sky130_fd_sc_hd__and3_1 _13455_ (.A(_02840_),
    .B(_02839_),
    .C(_02837_),
    .X(_02849_));
 sky130_fd_sc_hd__nand4_2 _13456_ (.A(_02738_),
    .B(_02744_),
    .C(_02837_),
    .D(_02839_),
    .Y(_02850_));
 sky130_fd_sc_hd__o21ai_1 _13457_ (.A1(_02838_),
    .A2(_02845_),
    .B1(_02844_),
    .Y(_02851_));
 sky130_fd_sc_hd__o21a_1 _13458_ (.A1(_01835_),
    .A2(_01977_),
    .B1(_02683_),
    .X(_02853_));
 sky130_fd_sc_hd__o21ai_1 _13459_ (.A1(_02679_),
    .A2(_02680_),
    .B1(_02683_),
    .Y(_02854_));
 sky130_fd_sc_hd__o31a_1 _13460_ (.A1(_01835_),
    .A2(_01977_),
    .A3(_02680_),
    .B1(_02683_),
    .X(_02855_));
 sky130_fd_sc_hd__nand2_1 _13461_ (.A(net62),
    .B(net7),
    .Y(_02856_));
 sky130_fd_sc_hd__nand2_2 _13462_ (.A(net61),
    .B(net7),
    .Y(_02857_));
 sky130_fd_sc_hd__and4_1 _13463_ (.A(net61),
    .B(net62),
    .C(net6),
    .D(net7),
    .X(_02858_));
 sky130_fd_sc_hd__nand4_1 _13464_ (.A(net61),
    .B(net62),
    .C(net6),
    .D(net7),
    .Y(_02859_));
 sky130_fd_sc_hd__a22o_1 _13465_ (.A1(net62),
    .A2(net6),
    .B1(net7),
    .B2(net61),
    .X(_02860_));
 sky130_fd_sc_hd__a2bb2oi_1 _13466_ (.A1_N(_01890_),
    .A2_N(_01956_),
    .B1(_02859_),
    .B2(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__o2bb2ai_1 _13467_ (.A1_N(_02859_),
    .A2_N(_02860_),
    .B1(_01890_),
    .B2(_01956_),
    .Y(_02862_));
 sky130_fd_sc_hd__o2111a_1 _13468_ (.A1(_02635_),
    .A2(_02856_),
    .B1(net63),
    .C1(net5),
    .D1(_02860_),
    .X(_02864_));
 sky130_fd_sc_hd__o2111ai_2 _13469_ (.A1(_02635_),
    .A2(_02856_),
    .B1(net63),
    .C1(net5),
    .D1(_02860_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _13470_ (.A(_02862_),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__o22ai_4 _13471_ (.A1(_02680_),
    .A2(_02853_),
    .B1(_02861_),
    .B2(_02864_),
    .Y(_02867_));
 sky130_fd_sc_hd__and3_4 _13472_ (.A(_02862_),
    .B(_02865_),
    .C(_02854_),
    .X(_02868_));
 sky130_fd_sc_hd__nand3_1 _13473_ (.A(_02862_),
    .B(_02865_),
    .C(_02854_),
    .Y(_02869_));
 sky130_fd_sc_hd__o22a_1 _13474_ (.A1(_01890_),
    .A2(_01945_),
    .B1(_02372_),
    .B2(_02635_),
    .X(_02870_));
 sky130_fd_sc_hd__a211o_1 _13475_ (.A1(_02372_),
    .A2(_02635_),
    .B1(_01890_),
    .C1(_01945_),
    .X(_02871_));
 sky130_fd_sc_hd__a31o_1 _13476_ (.A1(_02639_),
    .A2(net4),
    .A3(net63),
    .B1(_02636_),
    .X(_02872_));
 sky130_fd_sc_hd__o2bb2ai_4 _13477_ (.A1_N(_02867_),
    .A2_N(_02869_),
    .B1(_02870_),
    .B2(_02638_),
    .Y(_02873_));
 sky130_fd_sc_hd__a22oi_4 _13478_ (.A1(_02637_),
    .A2(_02871_),
    .B1(_02866_),
    .B2(_02855_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_2 _13479_ (.A(_02867_),
    .B(_02872_),
    .Y(_02876_));
 sky130_fd_sc_hd__o21ai_1 _13480_ (.A1(_02855_),
    .A2(_02866_),
    .B1(_02875_),
    .Y(_02877_));
 sky130_fd_sc_hd__o21ai_4 _13481_ (.A1(_02868_),
    .A2(_02876_),
    .B1(_02873_),
    .Y(_02878_));
 sky130_fd_sc_hd__o21ai_1 _13482_ (.A1(_02391_),
    .A2(_02663_),
    .B1(_02662_),
    .Y(_02879_));
 sky130_fd_sc_hd__a21oi_2 _13483_ (.A1(_02391_),
    .A2(_02663_),
    .B1(_02662_),
    .Y(_02880_));
 sky130_fd_sc_hd__o21a_1 _13484_ (.A1(_02662_),
    .A2(_02664_),
    .B1(_02668_),
    .X(_02881_));
 sky130_fd_sc_hd__nand2_1 _13485_ (.A(net55),
    .B(net11),
    .Y(_02882_));
 sky130_fd_sc_hd__a22oi_4 _13486_ (.A1(net44),
    .A2(net13),
    .B1(net14),
    .B2(net33),
    .Y(_02883_));
 sky130_fd_sc_hd__a22o_2 _13487_ (.A1(net44),
    .A2(net13),
    .B1(net14),
    .B2(net33),
    .X(_02884_));
 sky130_fd_sc_hd__and4_1 _13488_ (.A(net33),
    .B(net44),
    .C(net13),
    .D(net14),
    .X(_02886_));
 sky130_fd_sc_hd__nand4_4 _13489_ (.A(net33),
    .B(net44),
    .C(net13),
    .D(net14),
    .Y(_02887_));
 sky130_fd_sc_hd__o211ai_2 _13490_ (.A1(_01780_),
    .A2(_02032_),
    .B1(_02884_),
    .C1(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__o21bai_2 _13491_ (.A1(_02883_),
    .A2(_02886_),
    .B1_N(_02882_),
    .Y(_02889_));
 sky130_fd_sc_hd__and4_2 _13492_ (.A(_02884_),
    .B(_02887_),
    .C(net55),
    .D(net11),
    .X(_02890_));
 sky130_fd_sc_hd__nand4_2 _13493_ (.A(_02884_),
    .B(_02887_),
    .C(net55),
    .D(net11),
    .Y(_02891_));
 sky130_fd_sc_hd__o22ai_4 _13494_ (.A1(_01780_),
    .A2(_02032_),
    .B1(_02883_),
    .B2(_02886_),
    .Y(_02892_));
 sky130_fd_sc_hd__o21ai_4 _13495_ (.A1(_02667_),
    .A2(_02880_),
    .B1(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__o211ai_4 _13496_ (.A1(_02667_),
    .A2(_02880_),
    .B1(_02891_),
    .C1(_02892_),
    .Y(_02894_));
 sky130_fd_sc_hd__a22oi_2 _13497_ (.A1(_02665_),
    .A2(_02879_),
    .B1(_02891_),
    .B2(_02892_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand3_4 _13498_ (.A(_02881_),
    .B(_02888_),
    .C(_02889_),
    .Y(_02897_));
 sky130_fd_sc_hd__nand2_1 _13499_ (.A(net60),
    .B(net8),
    .Y(_02898_));
 sky130_fd_sc_hd__a22oi_4 _13500_ (.A1(net59),
    .A2(net9),
    .B1(net10),
    .B2(net58),
    .Y(_02899_));
 sky130_fd_sc_hd__a22o_2 _13501_ (.A1(net59),
    .A2(net9),
    .B1(net10),
    .B2(net58),
    .X(_02900_));
 sky130_fd_sc_hd__and4_1 _13502_ (.A(net58),
    .B(net59),
    .C(net9),
    .D(net10),
    .X(_02901_));
 sky130_fd_sc_hd__nand4_4 _13503_ (.A(net58),
    .B(net59),
    .C(net9),
    .D(net10),
    .Y(_02902_));
 sky130_fd_sc_hd__and3_1 _13504_ (.A(_02898_),
    .B(_02900_),
    .C(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__o211a_1 _13505_ (.A1(_02899_),
    .A2(_02901_),
    .B1(net60),
    .C1(net8),
    .X(_02904_));
 sky130_fd_sc_hd__a22oi_4 _13506_ (.A1(net60),
    .A2(net8),
    .B1(_02900_),
    .B2(_02902_),
    .Y(_02905_));
 sky130_fd_sc_hd__a22o_1 _13507_ (.A1(net60),
    .A2(net8),
    .B1(_02900_),
    .B2(_02902_),
    .X(_02906_));
 sky130_fd_sc_hd__a41oi_1 _13508_ (.A1(net58),
    .A2(net59),
    .A3(net9),
    .A4(net10),
    .B1(_02898_),
    .Y(_02908_));
 sky130_fd_sc_hd__a41o_1 _13509_ (.A1(net58),
    .A2(net59),
    .A3(net9),
    .A4(net10),
    .B1(_02898_),
    .X(_02909_));
 sky130_fd_sc_hd__and4_1 _13510_ (.A(_02900_),
    .B(_02902_),
    .C(net60),
    .D(net8),
    .X(_02910_));
 sky130_fd_sc_hd__o21ai_2 _13511_ (.A1(_02899_),
    .A2(_02909_),
    .B1(_02906_),
    .Y(_02911_));
 sky130_fd_sc_hd__a21oi_1 _13512_ (.A1(_02900_),
    .A2(_02908_),
    .B1(_02905_),
    .Y(_02912_));
 sky130_fd_sc_hd__o2bb2ai_2 _13513_ (.A1_N(_02894_),
    .A2_N(_02897_),
    .B1(_02903_),
    .B2(_02904_),
    .Y(_02913_));
 sky130_fd_sc_hd__o221ai_4 _13514_ (.A1(_02905_),
    .A2(_02910_),
    .B1(_02890_),
    .B2(_02893_),
    .C1(_02897_),
    .Y(_02914_));
 sky130_fd_sc_hd__o2bb2ai_2 _13515_ (.A1_N(_02894_),
    .A2_N(_02897_),
    .B1(_02905_),
    .B2(_02910_),
    .Y(_02915_));
 sky130_fd_sc_hd__o2111ai_4 _13516_ (.A1(_02899_),
    .A2(_02909_),
    .B1(_02906_),
    .C1(_02894_),
    .D1(_02897_),
    .Y(_02916_));
 sky130_fd_sc_hd__a32oi_4 _13517_ (.A1(_02660_),
    .A2(_02672_),
    .A3(_02673_),
    .B1(_02675_),
    .B2(_02694_),
    .Y(_02917_));
 sky130_fd_sc_hd__o22ai_4 _13518_ (.A1(_02671_),
    .A2(_02676_),
    .B1(_02693_),
    .B2(_02674_),
    .Y(_02919_));
 sky130_fd_sc_hd__and3_1 _13519_ (.A(_02913_),
    .B(_02917_),
    .C(_02914_),
    .X(_02920_));
 sky130_fd_sc_hd__nand3_2 _13520_ (.A(_02913_),
    .B(_02917_),
    .C(_02914_),
    .Y(_02921_));
 sky130_fd_sc_hd__and3_1 _13521_ (.A(_02915_),
    .B(_02916_),
    .C(_02919_),
    .X(_02922_));
 sky130_fd_sc_hd__nand3_4 _13522_ (.A(_02915_),
    .B(_02916_),
    .C(_02919_),
    .Y(_02923_));
 sky130_fd_sc_hd__a21o_2 _13523_ (.A1(_02921_),
    .A2(_02923_),
    .B1(_02878_),
    .X(_02924_));
 sky130_fd_sc_hd__nand3_4 _13524_ (.A(_02878_),
    .B(_02921_),
    .C(_02923_),
    .Y(_02925_));
 sky130_fd_sc_hd__a22o_1 _13525_ (.A1(_02873_),
    .A2(_02877_),
    .B1(_02921_),
    .B2(_02923_),
    .X(_02926_));
 sky130_fd_sc_hd__o211ai_2 _13526_ (.A1(_02876_),
    .A2(_02868_),
    .B1(_02873_),
    .C1(_02921_),
    .Y(_02927_));
 sky130_fd_sc_hd__o2111ai_1 _13527_ (.A1(_02876_),
    .A2(_02868_),
    .B1(_02873_),
    .C1(_02921_),
    .D1(_02923_),
    .Y(_02928_));
 sky130_fd_sc_hd__a2bb2oi_4 _13528_ (.A1_N(_02698_),
    .A2_N(_02704_),
    .B1(_02703_),
    .B2(_02657_),
    .Y(_02930_));
 sky130_fd_sc_hd__a22oi_4 _13529_ (.A1(_02706_),
    .A2(_02712_),
    .B1(_02924_),
    .B2(_02925_),
    .Y(_02931_));
 sky130_fd_sc_hd__o221ai_4 _13530_ (.A1(_02922_),
    .A2(_02927_),
    .B1(_02705_),
    .B2(_02711_),
    .C1(_02926_),
    .Y(_02932_));
 sky130_fd_sc_hd__a21boi_2 _13531_ (.A1(_02926_),
    .A2(_02928_),
    .B1_N(_02930_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand3_4 _13532_ (.A(_02924_),
    .B(_02930_),
    .C(_02925_),
    .Y(_02934_));
 sky130_fd_sc_hd__a32oi_4 _13533_ (.A1(_02924_),
    .A2(_02930_),
    .A3(_02925_),
    .B1(_02848_),
    .B2(_02850_),
    .Y(_02935_));
 sky130_fd_sc_hd__o211a_2 _13534_ (.A1(_02847_),
    .A2(_02849_),
    .B1(_02932_),
    .C1(_02934_),
    .X(_02936_));
 sky130_fd_sc_hd__o2111ai_4 _13535_ (.A1(_02845_),
    .A2(_02838_),
    .B1(_02844_),
    .C1(_02932_),
    .D1(_02934_),
    .Y(_02937_));
 sky130_fd_sc_hd__a21boi_1 _13536_ (.A1(_02932_),
    .A2(_02934_),
    .B1_N(_02851_),
    .Y(_02938_));
 sky130_fd_sc_hd__o22ai_4 _13537_ (.A1(_02843_),
    .A2(_02846_),
    .B1(_02931_),
    .B2(_02933_),
    .Y(_02939_));
 sky130_fd_sc_hd__nand2_1 _13538_ (.A(_02802_),
    .B(_02939_),
    .Y(_02941_));
 sky130_fd_sc_hd__nand3_2 _13539_ (.A(_02802_),
    .B(_02937_),
    .C(_02939_),
    .Y(_02942_));
 sky130_fd_sc_hd__a2bb2oi_2 _13540_ (.A1_N(_02714_),
    .A2_N(_02801_),
    .B1(_02937_),
    .B2(_02939_),
    .Y(_02943_));
 sky130_fd_sc_hd__o22ai_4 _13541_ (.A1(_02714_),
    .A2(_02801_),
    .B1(_02936_),
    .B2(_02938_),
    .Y(_02944_));
 sky130_fd_sc_hd__o21ai_1 _13542_ (.A1(_02718_),
    .A2(_02720_),
    .B1(_02719_),
    .Y(_02945_));
 sky130_fd_sc_hd__o21a_1 _13543_ (.A1(_02718_),
    .A2(_02720_),
    .B1(_02719_),
    .X(_02946_));
 sky130_fd_sc_hd__nor2_1 _13544_ (.A(_01769_),
    .B(_02010_),
    .Y(_02947_));
 sky130_fd_sc_hd__a22oi_2 _13545_ (.A1(net29),
    .A2(net39),
    .B1(net40),
    .B2(net28),
    .Y(_02948_));
 sky130_fd_sc_hd__a22o_1 _13546_ (.A1(net29),
    .A2(net39),
    .B1(net40),
    .B2(net28),
    .X(_02949_));
 sky130_fd_sc_hd__and4_1 _13547_ (.A(net28),
    .B(net29),
    .C(net39),
    .D(net40),
    .X(_02950_));
 sky130_fd_sc_hd__nand4_2 _13548_ (.A(net28),
    .B(net29),
    .C(net39),
    .D(net40),
    .Y(_02952_));
 sky130_fd_sc_hd__o211ai_1 _13549_ (.A1(_01769_),
    .A2(_02010_),
    .B1(_02949_),
    .C1(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__o21ai_1 _13550_ (.A1(_02948_),
    .A2(_02950_),
    .B1(_02947_),
    .Y(_02954_));
 sky130_fd_sc_hd__a22o_1 _13551_ (.A1(net27),
    .A2(net41),
    .B1(_02949_),
    .B2(_02952_),
    .X(_02955_));
 sky130_fd_sc_hd__and3_1 _13552_ (.A(_02947_),
    .B(_02949_),
    .C(_02952_),
    .X(_02956_));
 sky130_fd_sc_hd__nand4_1 _13553_ (.A(_02949_),
    .B(_02952_),
    .C(net27),
    .D(net41),
    .Y(_02957_));
 sky130_fd_sc_hd__nand3_2 _13554_ (.A(_02946_),
    .B(_02953_),
    .C(_02954_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand2_1 _13555_ (.A(_02955_),
    .B(_02945_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand3_1 _13556_ (.A(_02955_),
    .B(_02957_),
    .C(_02945_),
    .Y(_02960_));
 sky130_fd_sc_hd__o22a_1 _13557_ (.A1(_01791_),
    .A2(_02010_),
    .B1(_02505_),
    .B2(_02581_),
    .X(_02961_));
 sky130_fd_sc_hd__a2bb2o_1 _13558_ (.A1_N(_02505_),
    .A2_N(_02581_),
    .B1(_02584_),
    .B2(_02580_),
    .X(_02963_));
 sky130_fd_sc_hd__o2bb2ai_2 _13559_ (.A1_N(_02958_),
    .A2_N(_02960_),
    .B1(_02961_),
    .B2(_02583_),
    .Y(_02964_));
 sky130_fd_sc_hd__nand3_2 _13560_ (.A(_02958_),
    .B(_02960_),
    .C(_02963_),
    .Y(_02965_));
 sky130_fd_sc_hd__o21ai_2 _13561_ (.A1(_02576_),
    .A2(_02593_),
    .B1(_02592_),
    .Y(_02966_));
 sky130_fd_sc_hd__a21oi_4 _13562_ (.A1(_02964_),
    .A2(_02965_),
    .B1(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__a21o_1 _13563_ (.A1(_02964_),
    .A2(_02965_),
    .B1(_02966_),
    .X(_02968_));
 sky130_fd_sc_hd__o211a_2 _13564_ (.A1(_02591_),
    .A2(_02595_),
    .B1(_02964_),
    .C1(_02965_),
    .X(_02969_));
 sky130_fd_sc_hd__o211ai_2 _13565_ (.A1(_02591_),
    .A2(_02595_),
    .B1(_02964_),
    .C1(_02965_),
    .Y(_02970_));
 sky130_fd_sc_hd__o2bb2ai_1 _13566_ (.A1_N(_02603_),
    .A2_N(_02606_),
    .B1(_02604_),
    .B2(_02493_),
    .Y(_02971_));
 sky130_fd_sc_hd__a21boi_1 _13567_ (.A1(_02606_),
    .A2(_02603_),
    .B1_N(_02605_),
    .Y(_02972_));
 sky130_fd_sc_hd__nand2_1 _13568_ (.A(net12),
    .B(net45),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_1 _13569_ (.A(net26),
    .B(net42),
    .Y(_02975_));
 sky130_fd_sc_hd__a22oi_2 _13570_ (.A1(net26),
    .A2(net42),
    .B1(net43),
    .B2(net23),
    .Y(_02976_));
 sky130_fd_sc_hd__a22o_1 _13571_ (.A1(net26),
    .A2(net42),
    .B1(net43),
    .B2(net23),
    .X(_02977_));
 sky130_fd_sc_hd__nand2_1 _13572_ (.A(net26),
    .B(net43),
    .Y(_02978_));
 sky130_fd_sc_hd__and4_1 _13573_ (.A(net26),
    .B(net23),
    .C(net42),
    .D(net43),
    .X(_02979_));
 sky130_fd_sc_hd__nand4_2 _13574_ (.A(net26),
    .B(net23),
    .C(net42),
    .D(net43),
    .Y(_02980_));
 sky130_fd_sc_hd__o211ai_1 _13575_ (.A1(_01824_),
    .A2(_02054_),
    .B1(_02977_),
    .C1(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__o21bai_1 _13576_ (.A1(_02976_),
    .A2(_02979_),
    .B1_N(_02974_),
    .Y(_02982_));
 sky130_fd_sc_hd__o21ai_1 _13577_ (.A1(_02976_),
    .A2(_02979_),
    .B1(_02974_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand4_1 _13578_ (.A(_02977_),
    .B(_02980_),
    .C(net12),
    .D(net45),
    .Y(_02985_));
 sky130_fd_sc_hd__nand3_1 _13579_ (.A(_02972_),
    .B(_02981_),
    .C(_02982_),
    .Y(_02986_));
 sky130_fd_sc_hd__nand3_1 _13580_ (.A(_02983_),
    .B(_02985_),
    .C(_02971_),
    .Y(_02987_));
 sky130_fd_sc_hd__and2_1 _13581_ (.A(net1),
    .B(net46),
    .X(_02988_));
 sky130_fd_sc_hd__nand2_2 _13582_ (.A(net1),
    .B(net46),
    .Y(_02989_));
 sky130_fd_sc_hd__a21oi_1 _13583_ (.A1(_02986_),
    .A2(_02987_),
    .B1(_02988_),
    .Y(_02990_));
 sky130_fd_sc_hd__and3_1 _13584_ (.A(_02986_),
    .B(_02987_),
    .C(_02988_),
    .X(_02991_));
 sky130_fd_sc_hd__nor2_1 _13585_ (.A(_02990_),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__o21bai_4 _13586_ (.A1(_02967_),
    .A2(_02969_),
    .B1_N(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__nand2_1 _13587_ (.A(_02992_),
    .B(_02970_),
    .Y(_02994_));
 sky130_fd_sc_hd__and3_1 _13588_ (.A(_02968_),
    .B(_02992_),
    .C(_02970_),
    .X(_02996_));
 sky130_fd_sc_hd__nand3_1 _13589_ (.A(_02968_),
    .B(_02970_),
    .C(_02992_),
    .Y(_02997_));
 sky130_fd_sc_hd__a21boi_4 _13590_ (.A1(_02748_),
    .A2(_02749_),
    .B1_N(_02747_),
    .Y(_02998_));
 sky130_fd_sc_hd__a21oi_2 _13591_ (.A1(_02993_),
    .A2(_02997_),
    .B1(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21o_2 _13592_ (.A1(_02993_),
    .A2(_02997_),
    .B1(_02998_),
    .X(_03000_));
 sky130_fd_sc_hd__o211a_1 _13593_ (.A1(_02994_),
    .A2(_02967_),
    .B1(_02993_),
    .C1(_02998_),
    .X(_03001_));
 sky130_fd_sc_hd__o211ai_4 _13594_ (.A1(_02994_),
    .A2(_02967_),
    .B1(_02993_),
    .C1(_02998_),
    .Y(_03002_));
 sky130_fd_sc_hd__nand2_2 _13595_ (.A(_02602_),
    .B(_02614_),
    .Y(_03003_));
 sky130_fd_sc_hd__and2_1 _13596_ (.A(_02601_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__nand2_1 _13597_ (.A(_02601_),
    .B(_03003_),
    .Y(_03005_));
 sky130_fd_sc_hd__a21oi_1 _13598_ (.A1(_03000_),
    .A2(_03002_),
    .B1(_03004_),
    .Y(_03007_));
 sky130_fd_sc_hd__o21ai_1 _13599_ (.A1(_02999_),
    .A2(_03001_),
    .B1(_03005_),
    .Y(_03008_));
 sky130_fd_sc_hd__and3_1 _13600_ (.A(_03000_),
    .B(_03002_),
    .C(_03004_),
    .X(_03009_));
 sky130_fd_sc_hd__nand4_4 _13601_ (.A(_02601_),
    .B(_03000_),
    .C(_03002_),
    .D(_03003_),
    .Y(_03010_));
 sky130_fd_sc_hd__and3_1 _13602_ (.A(_03000_),
    .B(_03002_),
    .C(_03005_),
    .X(_03011_));
 sky130_fd_sc_hd__nand3_1 _13603_ (.A(_03000_),
    .B(_03002_),
    .C(_03005_),
    .Y(_03012_));
 sky130_fd_sc_hd__o211a_1 _13604_ (.A1(_02999_),
    .A2(_03001_),
    .B1(_03003_),
    .C1(_02601_),
    .X(_03013_));
 sky130_fd_sc_hd__o21ai_1 _13605_ (.A1(_02999_),
    .A2(_03001_),
    .B1(_03004_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_1 _13606_ (.A(_03012_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand2_1 _13607_ (.A(_03008_),
    .B(_03010_),
    .Y(_03016_));
 sky130_fd_sc_hd__nand4_2 _13608_ (.A(_02942_),
    .B(_02944_),
    .C(_03012_),
    .D(_03014_),
    .Y(_03018_));
 sky130_fd_sc_hd__o2bb2ai_1 _13609_ (.A1_N(_02942_),
    .A2_N(_02944_),
    .B1(_03011_),
    .B2(_03013_),
    .Y(_03019_));
 sky130_fd_sc_hd__o2bb2a_1 _13610_ (.A1_N(_02942_),
    .A2_N(_02944_),
    .B1(_03007_),
    .B2(_03009_),
    .X(_03020_));
 sky130_fd_sc_hd__o2bb2ai_1 _13611_ (.A1_N(_02942_),
    .A2_N(_02944_),
    .B1(_03007_),
    .B2(_03009_),
    .Y(_03021_));
 sky130_fd_sc_hd__nand4_1 _13612_ (.A(_02942_),
    .B(_02944_),
    .C(_03008_),
    .D(_03010_),
    .Y(_03022_));
 sky130_fd_sc_hd__o211ai_4 _13613_ (.A1(_02766_),
    .A2(_02799_),
    .B1(_03018_),
    .C1(_03019_),
    .Y(_03023_));
 sky130_fd_sc_hd__nand2_1 _13614_ (.A(_02800_),
    .B(_03022_),
    .Y(_03024_));
 sky130_fd_sc_hd__and3_1 _13615_ (.A(_02800_),
    .B(_03021_),
    .C(_03022_),
    .X(_03025_));
 sky130_fd_sc_hd__nand3_1 _13616_ (.A(_02800_),
    .B(_03021_),
    .C(_03022_),
    .Y(_03026_));
 sky130_fd_sc_hd__a21boi_2 _13617_ (.A1(_02621_),
    .A2(_02625_),
    .B1_N(_02623_),
    .Y(_03027_));
 sky130_fd_sc_hd__a21o_2 _13618_ (.A1(_02623_),
    .A2(_02627_),
    .B1(_02610_),
    .X(_03029_));
 sky130_fd_sc_hd__inv_2 _13619_ (.A(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand2_1 _13620_ (.A(_03027_),
    .B(_02610_),
    .Y(_03031_));
 sky130_fd_sc_hd__and2_2 _13621_ (.A(_03029_),
    .B(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__a21o_1 _13622_ (.A1(_03023_),
    .A2(_03026_),
    .B1(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__nand2_1 _13623_ (.A(_03023_),
    .B(_03032_),
    .Y(_03034_));
 sky130_fd_sc_hd__o211ai_1 _13624_ (.A1(_03020_),
    .A2(_03024_),
    .B1(_03032_),
    .C1(_03023_),
    .Y(_03035_));
 sky130_fd_sc_hd__a21o_1 _13625_ (.A1(_02775_),
    .A2(_02572_),
    .B1(_02772_),
    .X(_03036_));
 sky130_fd_sc_hd__a21oi_1 _13626_ (.A1(_03033_),
    .A2(_03035_),
    .B1(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__a21o_1 _13627_ (.A1(_03033_),
    .A2(_03035_),
    .B1(_03036_),
    .X(_03038_));
 sky130_fd_sc_hd__o211a_2 _13628_ (.A1(_03025_),
    .A2(_03034_),
    .B1(_03036_),
    .C1(_03033_),
    .X(_03040_));
 sky130_fd_sc_hd__o211ai_2 _13629_ (.A1(_03025_),
    .A2(_03034_),
    .B1(_03036_),
    .C1(_03033_),
    .Y(_03041_));
 sky130_fd_sc_hd__nand2_1 _13630_ (.A(_03038_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__o21ai_1 _13631_ (.A1(_03037_),
    .A2(_03040_),
    .B1(_02781_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand3b_2 _13632_ (.A_N(_02781_),
    .B(_03038_),
    .C(_03041_),
    .Y(_03044_));
 sky130_fd_sc_hd__nand2_1 _13633_ (.A(_03043_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand3_2 _13634_ (.A(_02783_),
    .B(_03043_),
    .C(_03044_),
    .Y(_03046_));
 sky130_fd_sc_hd__nand4b_2 _13635_ (.A_N(_02559_),
    .B(_02781_),
    .C(_02782_),
    .D(_03042_),
    .Y(_03047_));
 sky130_fd_sc_hd__nand2_1 _13636_ (.A(_03046_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__o211ai_1 _13637_ (.A1(_02786_),
    .A2(_02796_),
    .B1(_03046_),
    .C1(_03047_),
    .Y(_03049_));
 sky130_fd_sc_hd__a211o_1 _13638_ (.A1(_03046_),
    .A2(_03047_),
    .B1(_02786_),
    .C1(_02796_),
    .X(_03051_));
 sky130_fd_sc_hd__nand2_1 _13639_ (.A(_03049_),
    .B(_03051_),
    .Y(net78));
 sky130_fd_sc_hd__a21oi_2 _13640_ (.A1(_03046_),
    .A2(_03047_),
    .B1(_02789_),
    .Y(_03052_));
 sky130_fd_sc_hd__nand3_1 _13641_ (.A(_02785_),
    .B(_02788_),
    .C(_03048_),
    .Y(_03053_));
 sky130_fd_sc_hd__a21oi_2 _13642_ (.A1(_02783_),
    .A2(_02788_),
    .B1(_03045_),
    .Y(_03054_));
 sky130_fd_sc_hd__a21o_1 _13643_ (.A1(_02796_),
    .A2(_03048_),
    .B1(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__o2bb2ai_1 _13644_ (.A1_N(_03032_),
    .A2_N(_03023_),
    .B1(_03020_),
    .B2(_03024_),
    .Y(_03056_));
 sky130_fd_sc_hd__a21boi_4 _13645_ (.A1(_03023_),
    .A2(_03032_),
    .B1_N(_03026_),
    .Y(_03057_));
 sky130_fd_sc_hd__a21boi_4 _13646_ (.A1(_03015_),
    .A2(_02944_),
    .B1_N(_02942_),
    .Y(_03058_));
 sky130_fd_sc_hd__o22ai_4 _13647_ (.A1(_02936_),
    .A2(_02941_),
    .B1(_02943_),
    .B2(_03016_),
    .Y(_03059_));
 sky130_fd_sc_hd__o31a_1 _13648_ (.A1(_02967_),
    .A2(_02990_),
    .A3(_02991_),
    .B1(_02970_),
    .X(_03061_));
 sky130_fd_sc_hd__nand2_1 _13649_ (.A(net12),
    .B(net47),
    .Y(_03062_));
 sky130_fd_sc_hd__or3_2 _13650_ (.A(_01824_),
    .B(_02087_),
    .C(_02989_),
    .X(_03063_));
 sky130_fd_sc_hd__a22o_1 _13651_ (.A1(net12),
    .A2(net46),
    .B1(net47),
    .B2(net1),
    .X(_03064_));
 sky130_fd_sc_hd__o21ai_2 _13652_ (.A1(_02974_),
    .A2(_02976_),
    .B1(_02980_),
    .Y(_03065_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(net23),
    .B(net45),
    .Y(_03066_));
 sky130_fd_sc_hd__nand2_1 _13654_ (.A(net27),
    .B(net43),
    .Y(_03067_));
 sky130_fd_sc_hd__and4_1 _13655_ (.A(net27),
    .B(net26),
    .C(net42),
    .D(net43),
    .X(_03068_));
 sky130_fd_sc_hd__nand2_1 _13656_ (.A(net27),
    .B(net42),
    .Y(_03069_));
 sky130_fd_sc_hd__a22o_1 _13657_ (.A1(net27),
    .A2(net42),
    .B1(net43),
    .B2(net26),
    .X(_03070_));
 sky130_fd_sc_hd__o2bb2ai_1 _13658_ (.A1_N(_02978_),
    .A2_N(_03069_),
    .B1(_03067_),
    .B2(_02975_),
    .Y(_03071_));
 sky130_fd_sc_hd__o221ai_2 _13659_ (.A1(_01802_),
    .A2(_02054_),
    .B1(_02975_),
    .B2(_03067_),
    .C1(_03070_),
    .Y(_03072_));
 sky130_fd_sc_hd__nand3_1 _13660_ (.A(_03071_),
    .B(net45),
    .C(net23),
    .Y(_03073_));
 sky130_fd_sc_hd__a211o_1 _13661_ (.A1(_02978_),
    .A2(_03069_),
    .B1(_03066_),
    .C1(_03068_),
    .X(_03074_));
 sky130_fd_sc_hd__o21ai_2 _13662_ (.A1(_01802_),
    .A2(_02054_),
    .B1(_03071_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand3_4 _13663_ (.A(_03074_),
    .B(_03075_),
    .C(_03065_),
    .Y(_03076_));
 sky130_fd_sc_hd__nand3b_2 _13664_ (.A_N(_03065_),
    .B(_03072_),
    .C(_03073_),
    .Y(_03077_));
 sky130_fd_sc_hd__o311a_1 _13665_ (.A1(_01824_),
    .A2(_02087_),
    .A3(_02989_),
    .B1(_03064_),
    .C1(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__and4_1 _13666_ (.A(_03063_),
    .B(_03064_),
    .C(_03076_),
    .D(_03077_),
    .X(_03079_));
 sky130_fd_sc_hd__nand2_1 _13667_ (.A(_03078_),
    .B(_03076_),
    .Y(_03080_));
 sky130_fd_sc_hd__a22oi_2 _13668_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_03076_),
    .B2(_03077_),
    .Y(_03082_));
 sky130_fd_sc_hd__a21oi_1 _13669_ (.A1(_03078_),
    .A2(_03076_),
    .B1(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__o2bb2ai_2 _13670_ (.A1_N(_02963_),
    .A2_N(_02958_),
    .B1(_02956_),
    .B2(_02959_),
    .Y(_03084_));
 sky130_fd_sc_hd__o21ai_1 _13671_ (.A1(_02821_),
    .A2(_02822_),
    .B1(_02824_),
    .Y(_03085_));
 sky130_fd_sc_hd__o21a_1 _13672_ (.A1(_02821_),
    .A2(_02822_),
    .B1(_02824_),
    .X(_03086_));
 sky130_fd_sc_hd__nand2_1 _13673_ (.A(net28),
    .B(net41),
    .Y(_03087_));
 sky130_fd_sc_hd__nand2_1 _13674_ (.A(net30),
    .B(net39),
    .Y(_03088_));
 sky130_fd_sc_hd__a22oi_2 _13675_ (.A1(net30),
    .A2(net39),
    .B1(net40),
    .B2(net29),
    .Y(_03089_));
 sky130_fd_sc_hd__a22o_1 _13676_ (.A1(net30),
    .A2(net39),
    .B1(net40),
    .B2(net29),
    .X(_03090_));
 sky130_fd_sc_hd__and4_1 _13677_ (.A(net29),
    .B(net30),
    .C(net39),
    .D(net40),
    .X(_03091_));
 sky130_fd_sc_hd__nand4_2 _13678_ (.A(net29),
    .B(net30),
    .C(net39),
    .D(net40),
    .Y(_03093_));
 sky130_fd_sc_hd__o211ai_1 _13679_ (.A1(_01748_),
    .A2(_02010_),
    .B1(_03090_),
    .C1(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__o21bai_1 _13680_ (.A1(_03089_),
    .A2(_03091_),
    .B1_N(_03087_),
    .Y(_03095_));
 sky130_fd_sc_hd__o21ai_1 _13681_ (.A1(_03089_),
    .A2(_03091_),
    .B1(_03087_),
    .Y(_03096_));
 sky130_fd_sc_hd__and4_1 _13682_ (.A(_03090_),
    .B(_03093_),
    .C(net28),
    .D(net41),
    .X(_03097_));
 sky130_fd_sc_hd__nand4_1 _13683_ (.A(_03090_),
    .B(_03093_),
    .C(net28),
    .D(net41),
    .Y(_03098_));
 sky130_fd_sc_hd__nand3_2 _13684_ (.A(_03086_),
    .B(_03094_),
    .C(_03095_),
    .Y(_03099_));
 sky130_fd_sc_hd__nand2_1 _13685_ (.A(_03096_),
    .B(_03085_),
    .Y(_03100_));
 sky130_fd_sc_hd__nand3_2 _13686_ (.A(_03096_),
    .B(_03098_),
    .C(_03085_),
    .Y(_03101_));
 sky130_fd_sc_hd__inv_2 _13687_ (.A(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__o21a_1 _13688_ (.A1(_01769_),
    .A2(_02010_),
    .B1(_02952_),
    .X(_03104_));
 sky130_fd_sc_hd__a31o_1 _13689_ (.A1(_02949_),
    .A2(net41),
    .A3(net27),
    .B1(_02950_),
    .X(_03105_));
 sky130_fd_sc_hd__o2bb2ai_2 _13690_ (.A1_N(_03099_),
    .A2_N(_03101_),
    .B1(_03104_),
    .B2(_02948_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2_2 _13691_ (.A(_03099_),
    .B(_03105_),
    .Y(_03107_));
 sky130_fd_sc_hd__nand3_1 _13692_ (.A(_03099_),
    .B(_03101_),
    .C(_03105_),
    .Y(_03108_));
 sky130_fd_sc_hd__a21oi_1 _13693_ (.A1(_03106_),
    .A2(_03108_),
    .B1(_03084_),
    .Y(_03109_));
 sky130_fd_sc_hd__a21o_1 _13694_ (.A1(_03106_),
    .A2(_03108_),
    .B1(_03084_),
    .X(_03110_));
 sky130_fd_sc_hd__o211a_1 _13695_ (.A1(_03107_),
    .A2(_03102_),
    .B1(_03084_),
    .C1(_03106_),
    .X(_03111_));
 sky130_fd_sc_hd__o211ai_4 _13696_ (.A1(_03107_),
    .A2(_03102_),
    .B1(_03084_),
    .C1(_03106_),
    .Y(_03112_));
 sky130_fd_sc_hd__o22ai_2 _13697_ (.A1(_03079_),
    .A2(_03082_),
    .B1(_03109_),
    .B2(_03111_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand3_2 _13698_ (.A(_03110_),
    .B(_03112_),
    .C(_03083_),
    .Y(_03115_));
 sky130_fd_sc_hd__nand2_2 _13699_ (.A(_03113_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__o21ai_2 _13700_ (.A1(_02842_),
    .A2(_02838_),
    .B1(_02837_),
    .Y(_03117_));
 sky130_fd_sc_hd__a21boi_1 _13701_ (.A1(_02840_),
    .A2(_02839_),
    .B1_N(_02837_),
    .Y(_03118_));
 sky130_fd_sc_hd__a21oi_1 _13702_ (.A1(_03113_),
    .A2(_03115_),
    .B1(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__o2111a_2 _13703_ (.A1(_02842_),
    .A2(_02838_),
    .B1(_02837_),
    .C1(_03115_),
    .D1(_03113_),
    .X(_03120_));
 sky130_fd_sc_hd__o21a_2 _13704_ (.A1(_03119_),
    .A2(_03120_),
    .B1(_03061_),
    .X(_03121_));
 sky130_fd_sc_hd__o21ai_2 _13705_ (.A1(_03119_),
    .A2(_03120_),
    .B1(_03061_),
    .Y(_03122_));
 sky130_fd_sc_hd__o2bb2ai_4 _13706_ (.A1_N(_03117_),
    .A2_N(_03116_),
    .B1(_02996_),
    .B2(_02969_),
    .Y(_03123_));
 sky130_fd_sc_hd__nor2_2 _13707_ (.A(_03120_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__o21ai_4 _13708_ (.A1(_03120_),
    .A2(_03123_),
    .B1(_03122_),
    .Y(_03126_));
 sky130_fd_sc_hd__nand2_1 _13709_ (.A(_02851_),
    .B(_02932_),
    .Y(_03127_));
 sky130_fd_sc_hd__a32oi_1 _13710_ (.A1(_02915_),
    .A2(_02916_),
    .A3(_02919_),
    .B1(_02877_),
    .B2(_02873_),
    .Y(_03128_));
 sky130_fd_sc_hd__a32oi_4 _13711_ (.A1(_02913_),
    .A2(_02917_),
    .A3(_02914_),
    .B1(_02878_),
    .B2(_02923_),
    .Y(_03129_));
 sky130_fd_sc_hd__a32o_1 _13712_ (.A1(_02913_),
    .A2(_02917_),
    .A3(_02914_),
    .B1(_02878_),
    .B2(_02923_),
    .X(_03130_));
 sky130_fd_sc_hd__o21ai_1 _13713_ (.A1(_01780_),
    .A2(_02032_),
    .B1(_02887_),
    .Y(_03131_));
 sky130_fd_sc_hd__o21ai_4 _13714_ (.A1(_02882_),
    .A2(_02883_),
    .B1(_02887_),
    .Y(_03132_));
 sky130_fd_sc_hd__o21a_1 _13715_ (.A1(_02882_),
    .A2(_02883_),
    .B1(_02887_),
    .X(_03133_));
 sky130_fd_sc_hd__nand2_1 _13716_ (.A(net55),
    .B(net13),
    .Y(_03134_));
 sky130_fd_sc_hd__a22oi_4 _13717_ (.A1(net44),
    .A2(net14),
    .B1(net15),
    .B2(net33),
    .Y(_03135_));
 sky130_fd_sc_hd__a22o_2 _13718_ (.A1(net44),
    .A2(net14),
    .B1(net15),
    .B2(net33),
    .X(_03137_));
 sky130_fd_sc_hd__and4_1 _13719_ (.A(net33),
    .B(net44),
    .C(net14),
    .D(net15),
    .X(_03138_));
 sky130_fd_sc_hd__nand4_4 _13720_ (.A(net33),
    .B(net44),
    .C(net14),
    .D(net15),
    .Y(_03139_));
 sky130_fd_sc_hd__o211ai_2 _13721_ (.A1(_01780_),
    .A2(_02043_),
    .B1(_03137_),
    .C1(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__o21bai_1 _13722_ (.A1(_03135_),
    .A2(_03138_),
    .B1_N(_03134_),
    .Y(_03141_));
 sky130_fd_sc_hd__o22ai_4 _13723_ (.A1(_01780_),
    .A2(_02043_),
    .B1(_03135_),
    .B2(_03138_),
    .Y(_03142_));
 sky130_fd_sc_hd__a41o_1 _13724_ (.A1(net33),
    .A2(net44),
    .A3(net14),
    .A4(net15),
    .B1(_03134_),
    .X(_03143_));
 sky130_fd_sc_hd__and4_1 _13725_ (.A(_03137_),
    .B(_03139_),
    .C(net55),
    .D(net13),
    .X(_03144_));
 sky130_fd_sc_hd__nand4_4 _13726_ (.A(_03137_),
    .B(_03139_),
    .C(net55),
    .D(net13),
    .Y(_03145_));
 sky130_fd_sc_hd__a22oi_4 _13727_ (.A1(_02884_),
    .A2(_03131_),
    .B1(_03142_),
    .B2(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand3_4 _13728_ (.A(_03133_),
    .B(_03140_),
    .C(_03141_),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2_1 _13729_ (.A(_03142_),
    .B(_03132_),
    .Y(_03149_));
 sky130_fd_sc_hd__o211a_1 _13730_ (.A1(_03135_),
    .A2(_03143_),
    .B1(_03132_),
    .C1(_03142_),
    .X(_03150_));
 sky130_fd_sc_hd__o211ai_4 _13731_ (.A1(_03135_),
    .A2(_03143_),
    .B1(_03132_),
    .C1(_03142_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand2_1 _13732_ (.A(net60),
    .B(net9),
    .Y(_03152_));
 sky130_fd_sc_hd__a22oi_4 _13733_ (.A1(net59),
    .A2(net10),
    .B1(net11),
    .B2(net58),
    .Y(_03153_));
 sky130_fd_sc_hd__a22o_1 _13734_ (.A1(net59),
    .A2(net10),
    .B1(net11),
    .B2(net58),
    .X(_03154_));
 sky130_fd_sc_hd__and4_2 _13735_ (.A(net58),
    .B(net59),
    .C(net10),
    .D(net11),
    .X(_03155_));
 sky130_fd_sc_hd__nand4_1 _13736_ (.A(net58),
    .B(net59),
    .C(net10),
    .D(net11),
    .Y(_03156_));
 sky130_fd_sc_hd__and3_1 _13737_ (.A(_03152_),
    .B(_03154_),
    .C(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__o211ai_1 _13738_ (.A1(_01835_),
    .A2(_01999_),
    .B1(_03154_),
    .C1(_03156_),
    .Y(_03159_));
 sky130_fd_sc_hd__o211a_1 _13739_ (.A1(_03153_),
    .A2(_03155_),
    .B1(net60),
    .C1(net9),
    .X(_03160_));
 sky130_fd_sc_hd__o21bai_1 _13740_ (.A1(_03153_),
    .A2(_03155_),
    .B1_N(_03152_),
    .Y(_03161_));
 sky130_fd_sc_hd__o21ai_1 _13741_ (.A1(_03153_),
    .A2(_03155_),
    .B1(_03152_),
    .Y(_03162_));
 sky130_fd_sc_hd__a41o_1 _13742_ (.A1(net58),
    .A2(net59),
    .A3(net10),
    .A4(net11),
    .B1(_03152_),
    .X(_03163_));
 sky130_fd_sc_hd__o21ai_4 _13743_ (.A1(_03153_),
    .A2(_03163_),
    .B1(_03162_),
    .Y(_03164_));
 sky130_fd_sc_hd__nand2_2 _13744_ (.A(_03159_),
    .B(_03161_),
    .Y(_03165_));
 sky130_fd_sc_hd__o21ai_1 _13745_ (.A1(_03146_),
    .A2(_03150_),
    .B1(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__o211ai_2 _13746_ (.A1(_03144_),
    .A2(_03149_),
    .B1(_03164_),
    .C1(_03148_),
    .Y(_03167_));
 sky130_fd_sc_hd__a21oi_1 _13747_ (.A1(_03148_),
    .A2(_03151_),
    .B1(_03165_),
    .Y(_03168_));
 sky130_fd_sc_hd__o21ai_4 _13748_ (.A1(_03146_),
    .A2(_03150_),
    .B1(_03164_),
    .Y(_03170_));
 sky130_fd_sc_hd__and3_1 _13749_ (.A(_03148_),
    .B(_03151_),
    .C(_03165_),
    .X(_03171_));
 sky130_fd_sc_hd__o211ai_4 _13750_ (.A1(_03157_),
    .A2(_03160_),
    .B1(_03148_),
    .C1(_03151_),
    .Y(_03172_));
 sky130_fd_sc_hd__a21boi_2 _13751_ (.A1(_02897_),
    .A2(_02912_),
    .B1_N(_02894_),
    .Y(_03173_));
 sky130_fd_sc_hd__o22ai_4 _13752_ (.A1(_02893_),
    .A2(_02890_),
    .B1(_02911_),
    .B2(_02895_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand3_4 _13753_ (.A(_03170_),
    .B(_03172_),
    .C(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__a21oi_4 _13754_ (.A1(_03170_),
    .A2(_03172_),
    .B1(_03174_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand3_4 _13755_ (.A(_03166_),
    .B(_03173_),
    .C(_03167_),
    .Y(_03177_));
 sky130_fd_sc_hd__and3_1 _13756_ (.A(_02860_),
    .B(net5),
    .C(net63),
    .X(_03178_));
 sky130_fd_sc_hd__a31o_2 _13757_ (.A1(_02860_),
    .A2(net5),
    .A3(net63),
    .B1(_02858_),
    .X(_03179_));
 sky130_fd_sc_hd__a31o_1 _13758_ (.A1(_02900_),
    .A2(net8),
    .A3(net60),
    .B1(_02901_),
    .X(_03181_));
 sky130_fd_sc_hd__o21a_1 _13759_ (.A1(_02898_),
    .A2(_02899_),
    .B1(_02902_),
    .X(_03182_));
 sky130_fd_sc_hd__nand2_1 _13760_ (.A(net63),
    .B(net6),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2_2 _13761_ (.A(net62),
    .B(net8),
    .Y(_03184_));
 sky130_fd_sc_hd__nand4_1 _13762_ (.A(net61),
    .B(net62),
    .C(net7),
    .D(net8),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_2 _13763_ (.A(net61),
    .B(net8),
    .Y(_03186_));
 sky130_fd_sc_hd__a22o_2 _13764_ (.A1(net62),
    .A2(net7),
    .B1(net8),
    .B2(net61),
    .X(_03187_));
 sky130_fd_sc_hd__o2bb2ai_1 _13765_ (.A1_N(_02856_),
    .A2_N(_03186_),
    .B1(_03184_),
    .B2(_02857_),
    .Y(_03188_));
 sky130_fd_sc_hd__o221ai_4 _13766_ (.A1(_01890_),
    .A2(_01966_),
    .B1(_02857_),
    .B2(_03184_),
    .C1(_03187_),
    .Y(_03189_));
 sky130_fd_sc_hd__nand3_2 _13767_ (.A(_03188_),
    .B(net6),
    .C(net63),
    .Y(_03190_));
 sky130_fd_sc_hd__o2111ai_2 _13768_ (.A1(_02857_),
    .A2(_03184_),
    .B1(net63),
    .C1(net6),
    .D1(_03187_),
    .Y(_03192_));
 sky130_fd_sc_hd__a22o_1 _13769_ (.A1(net63),
    .A2(net6),
    .B1(_03185_),
    .B2(_03187_),
    .X(_03193_));
 sky130_fd_sc_hd__a21oi_4 _13770_ (.A1(_03189_),
    .A2(_03190_),
    .B1(_03182_),
    .Y(_03194_));
 sky130_fd_sc_hd__nand3_1 _13771_ (.A(_03193_),
    .B(_03181_),
    .C(_03192_),
    .Y(_03195_));
 sky130_fd_sc_hd__nand3_4 _13772_ (.A(_03182_),
    .B(_03189_),
    .C(_03190_),
    .Y(_03196_));
 sky130_fd_sc_hd__o21a_1 _13773_ (.A1(_02858_),
    .A2(_03178_),
    .B1(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__o21ai_1 _13774_ (.A1(_02858_),
    .A2(_03178_),
    .B1(_03196_),
    .Y(_03198_));
 sky130_fd_sc_hd__and3_1 _13775_ (.A(_03195_),
    .B(_03196_),
    .C(_03179_),
    .X(_03199_));
 sky130_fd_sc_hd__a21oi_2 _13776_ (.A1(_03195_),
    .A2(_03196_),
    .B1(_03179_),
    .Y(_03200_));
 sky130_fd_sc_hd__a21o_1 _13777_ (.A1(_03195_),
    .A2(_03196_),
    .B1(_03179_),
    .X(_03201_));
 sky130_fd_sc_hd__a21oi_1 _13778_ (.A1(_03195_),
    .A2(_03197_),
    .B1(_03200_),
    .Y(_03203_));
 sky130_fd_sc_hd__o21ai_4 _13779_ (.A1(_03194_),
    .A2(_03198_),
    .B1(_03201_),
    .Y(_03204_));
 sky130_fd_sc_hd__a21oi_1 _13780_ (.A1(_03175_),
    .A2(_03177_),
    .B1(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__a21o_1 _13781_ (.A1(_03175_),
    .A2(_03177_),
    .B1(_03204_),
    .X(_03206_));
 sky130_fd_sc_hd__and3_1 _13782_ (.A(_03175_),
    .B(_03177_),
    .C(_03204_),
    .X(_03207_));
 sky130_fd_sc_hd__o211ai_2 _13783_ (.A1(_03199_),
    .A2(_03200_),
    .B1(_03175_),
    .C1(_03177_),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(_03203_),
    .B(_03177_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand3_2 _13785_ (.A(_03203_),
    .B(_03177_),
    .C(_03175_),
    .Y(_03210_));
 sky130_fd_sc_hd__inv_2 _13786_ (.A(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__o2bb2ai_2 _13787_ (.A1_N(_03175_),
    .A2_N(_03177_),
    .B1(_03199_),
    .B2(_03200_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _13788_ (.A(_03212_),
    .B(_03129_),
    .Y(_03214_));
 sky130_fd_sc_hd__and3_1 _13789_ (.A(_03212_),
    .B(_03129_),
    .C(_03210_),
    .X(_03215_));
 sky130_fd_sc_hd__nand3_2 _13790_ (.A(_03212_),
    .B(_03129_),
    .C(_03210_),
    .Y(_03216_));
 sky130_fd_sc_hd__a2bb2oi_1 _13791_ (.A1_N(_02920_),
    .A2_N(_03128_),
    .B1(_03210_),
    .B2(_03212_),
    .Y(_03217_));
 sky130_fd_sc_hd__nand3_4 _13792_ (.A(_03130_),
    .B(_03206_),
    .C(_03208_),
    .Y(_03218_));
 sky130_fd_sc_hd__a21oi_2 _13793_ (.A1(_02867_),
    .A2(_02872_),
    .B1(_02868_),
    .Y(_03219_));
 sky130_fd_sc_hd__o21ai_4 _13794_ (.A1(_02807_),
    .A2(_02811_),
    .B1(_02810_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_2 _13795_ (.A(net3),
    .B(net35),
    .Y(_03221_));
 sky130_fd_sc_hd__and4_1 _13796_ (.A(net64),
    .B(net34),
    .C(net4),
    .D(net5),
    .X(_03222_));
 sky130_fd_sc_hd__nand4_4 _13797_ (.A(net64),
    .B(net34),
    .C(net4),
    .D(net5),
    .Y(_03223_));
 sky130_fd_sc_hd__a22oi_4 _13798_ (.A1(net34),
    .A2(net4),
    .B1(net5),
    .B2(net64),
    .Y(_03225_));
 sky130_fd_sc_hd__a22o_1 _13799_ (.A1(net34),
    .A2(net4),
    .B1(net5),
    .B2(net64),
    .X(_03226_));
 sky130_fd_sc_hd__o211ai_1 _13800_ (.A1(_01923_),
    .A2(_01934_),
    .B1(_03223_),
    .C1(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__o21bai_1 _13801_ (.A1(_03222_),
    .A2(_03225_),
    .B1_N(_03221_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand4_4 _13802_ (.A(_03226_),
    .B(net35),
    .C(net3),
    .D(_03223_),
    .Y(_03229_));
 sky130_fd_sc_hd__o21ai_4 _13803_ (.A1(_03222_),
    .A2(_03225_),
    .B1(_03221_),
    .Y(_03230_));
 sky130_fd_sc_hd__nand3_4 _13804_ (.A(_03230_),
    .B(_03220_),
    .C(_03229_),
    .Y(_03231_));
 sky130_fd_sc_hd__a21oi_4 _13805_ (.A1(_03229_),
    .A2(_03230_),
    .B1(_03220_),
    .Y(_03232_));
 sky130_fd_sc_hd__nand3b_2 _13806_ (.A_N(_03220_),
    .B(_03227_),
    .C(_03228_),
    .Y(_03233_));
 sky130_fd_sc_hd__a22oi_4 _13807_ (.A1(net2),
    .A2(net36),
    .B1(net37),
    .B2(net32),
    .Y(_03234_));
 sky130_fd_sc_hd__a22o_1 _13808_ (.A1(net2),
    .A2(net36),
    .B1(net37),
    .B2(net32),
    .X(_03236_));
 sky130_fd_sc_hd__nand4_4 _13809_ (.A(net2),
    .B(net32),
    .C(net36),
    .D(net37),
    .Y(_03237_));
 sky130_fd_sc_hd__nand2_1 _13810_ (.A(net31),
    .B(net38),
    .Y(_03238_));
 sky130_fd_sc_hd__a22oi_4 _13811_ (.A1(net31),
    .A2(net38),
    .B1(_03236_),
    .B2(_03237_),
    .Y(_03239_));
 sky130_fd_sc_hd__and4_1 _13812_ (.A(_03236_),
    .B(_03237_),
    .C(net31),
    .D(net38),
    .X(_03240_));
 sky130_fd_sc_hd__a21oi_2 _13813_ (.A1(_03236_),
    .A2(_03237_),
    .B1(_03238_),
    .Y(_03241_));
 sky130_fd_sc_hd__and3_1 _13814_ (.A(_03236_),
    .B(_03237_),
    .C(_03238_),
    .X(_03242_));
 sky130_fd_sc_hd__nor2_1 _13815_ (.A(_03241_),
    .B(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__o211ai_4 _13816_ (.A1(_03239_),
    .A2(_03240_),
    .B1(_03231_),
    .C1(_03233_),
    .Y(_03244_));
 sky130_fd_sc_hd__o2bb2ai_2 _13817_ (.A1_N(_03231_),
    .A2_N(_03233_),
    .B1(_03241_),
    .B2(_03242_),
    .Y(_03245_));
 sky130_fd_sc_hd__o2bb2ai_2 _13818_ (.A1_N(_03231_),
    .A2_N(_03233_),
    .B1(_03239_),
    .B2(_03240_),
    .Y(_03247_));
 sky130_fd_sc_hd__o21ai_2 _13819_ (.A1(_03241_),
    .A2(_03242_),
    .B1(_03231_),
    .Y(_03248_));
 sky130_fd_sc_hd__nand3_2 _13820_ (.A(_03219_),
    .B(_03244_),
    .C(_03245_),
    .Y(_03249_));
 sky130_fd_sc_hd__o221a_4 _13821_ (.A1(_03232_),
    .A2(_03248_),
    .B1(_02868_),
    .B2(_02875_),
    .C1(_03247_),
    .X(_03250_));
 sky130_fd_sc_hd__o221ai_4 _13822_ (.A1(_03232_),
    .A2(_03248_),
    .B1(_02868_),
    .B2(_02875_),
    .C1(_03247_),
    .Y(_03251_));
 sky130_fd_sc_hd__a32oi_4 _13823_ (.A1(_02806_),
    .A2(_02814_),
    .A3(_02816_),
    .B1(_02818_),
    .B2(_02832_),
    .Y(_03252_));
 sky130_fd_sc_hd__a32o_1 _13824_ (.A1(_02806_),
    .A2(_02814_),
    .A3(_02816_),
    .B1(_02818_),
    .B2(_02832_),
    .X(_03253_));
 sky130_fd_sc_hd__a21oi_2 _13825_ (.A1(_03249_),
    .A2(_03251_),
    .B1(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__a21o_1 _13826_ (.A1(_03249_),
    .A2(_03251_),
    .B1(_03253_),
    .X(_03255_));
 sky130_fd_sc_hd__a31oi_4 _13827_ (.A1(_03245_),
    .A2(_03219_),
    .A3(_03244_),
    .B1(_03252_),
    .Y(_03256_));
 sky130_fd_sc_hd__a31o_1 _13828_ (.A1(_03245_),
    .A2(_03219_),
    .A3(_03244_),
    .B1(_03252_),
    .X(_03258_));
 sky130_fd_sc_hd__and3_1 _13829_ (.A(_03249_),
    .B(_03251_),
    .C(_03253_),
    .X(_03259_));
 sky130_fd_sc_hd__a21oi_1 _13830_ (.A1(_03251_),
    .A2(_03256_),
    .B1(_03254_),
    .Y(_03260_));
 sky130_fd_sc_hd__o21ai_1 _13831_ (.A1(_03250_),
    .A2(_03258_),
    .B1(_03255_),
    .Y(_03261_));
 sky130_fd_sc_hd__o2bb2ai_4 _13832_ (.A1_N(_03216_),
    .A2_N(_03218_),
    .B1(_03254_),
    .B2(_03259_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _13833_ (.A(_03218_),
    .B(_03260_),
    .Y(_03263_));
 sky130_fd_sc_hd__o2111ai_4 _13834_ (.A1(_03250_),
    .A2(_03258_),
    .B1(_03255_),
    .C1(_03216_),
    .D1(_03218_),
    .Y(_03264_));
 sky130_fd_sc_hd__inv_2 _13835_ (.A(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__a22oi_4 _13836_ (.A1(_02934_),
    .A2(_03127_),
    .B1(_03262_),
    .B2(_03264_),
    .Y(_03266_));
 sky130_fd_sc_hd__a22o_1 _13837_ (.A1(_02934_),
    .A2(_03127_),
    .B1(_03262_),
    .B2(_03264_),
    .X(_03267_));
 sky130_fd_sc_hd__o21ai_4 _13838_ (.A1(_02931_),
    .A2(_02935_),
    .B1(_03262_),
    .Y(_03269_));
 sky130_fd_sc_hd__o221a_2 _13839_ (.A1(_02931_),
    .A2(_02935_),
    .B1(_03215_),
    .B2(_03263_),
    .C1(_03262_),
    .X(_03270_));
 sky130_fd_sc_hd__o221ai_4 _13840_ (.A1(_02931_),
    .A2(_02935_),
    .B1(_03215_),
    .B2(_03263_),
    .C1(_03262_),
    .Y(_03271_));
 sky130_fd_sc_hd__o211ai_2 _13841_ (.A1(_03123_),
    .A2(_03120_),
    .B1(_03122_),
    .C1(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__nand3b_1 _13842_ (.A_N(_03126_),
    .B(_03267_),
    .C(_03271_),
    .Y(_03273_));
 sky130_fd_sc_hd__o22ai_4 _13843_ (.A1(_03121_),
    .A2(_03124_),
    .B1(_03266_),
    .B2(_03270_),
    .Y(_03274_));
 sky130_fd_sc_hd__o221ai_4 _13844_ (.A1(_03121_),
    .A2(_03124_),
    .B1(_03269_),
    .B2(_03265_),
    .C1(_03267_),
    .Y(_03275_));
 sky130_fd_sc_hd__o21bai_4 _13845_ (.A1(_03266_),
    .A2(_03270_),
    .B1_N(_03126_),
    .Y(_03276_));
 sky130_fd_sc_hd__o211ai_4 _13846_ (.A1(_03266_),
    .A2(_03272_),
    .B1(_03274_),
    .C1(_03059_),
    .Y(_03277_));
 sky130_fd_sc_hd__o2111a_1 _13847_ (.A1(_02943_),
    .A2(_03016_),
    .B1(_03275_),
    .C1(_03276_),
    .D1(_02942_),
    .X(_03278_));
 sky130_fd_sc_hd__nand3_4 _13848_ (.A(_03058_),
    .B(_03275_),
    .C(_03276_),
    .Y(_03280_));
 sky130_fd_sc_hd__a21oi_2 _13849_ (.A1(_03000_),
    .A2(_03004_),
    .B1(_03001_),
    .Y(_03281_));
 sky130_fd_sc_hd__a21bo_1 _13850_ (.A1(_02986_),
    .A2(_02988_),
    .B1_N(_02987_),
    .X(_03282_));
 sky130_fd_sc_hd__a32o_2 _13851_ (.A1(_02972_),
    .A2(_02981_),
    .A3(_02982_),
    .B1(_02987_),
    .B2(_02989_),
    .X(_03283_));
 sky130_fd_sc_hd__a21oi_2 _13852_ (.A1(_03002_),
    .A2(_03010_),
    .B1(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__a21o_1 _13853_ (.A1(_03002_),
    .A2(_03010_),
    .B1(_03283_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_1 _13854_ (.A1(_03005_),
    .A2(_02999_),
    .B1(_03002_),
    .C1(_03283_),
    .X(_03286_));
 sky130_fd_sc_hd__a21oi_2 _13855_ (.A1(_03002_),
    .A2(_03010_),
    .B1(_03282_),
    .Y(_03287_));
 sky130_fd_sc_hd__and3_1 _13856_ (.A(_03002_),
    .B(_03010_),
    .C(_03282_),
    .X(_03288_));
 sky130_fd_sc_hd__nor2_1 _13857_ (.A(_03284_),
    .B(_03286_),
    .Y(_03289_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(_03287_),
    .B(_03288_),
    .Y(_03291_));
 sky130_fd_sc_hd__o2bb2ai_4 _13859_ (.A1_N(_03277_),
    .A2_N(_03280_),
    .B1(_03287_),
    .B2(_03288_),
    .Y(_03292_));
 sky130_fd_sc_hd__o211ai_4 _13860_ (.A1(_03284_),
    .A2(_03286_),
    .B1(_03277_),
    .C1(_03280_),
    .Y(_03293_));
 sky130_fd_sc_hd__o2bb2ai_1 _13861_ (.A1_N(_03277_),
    .A2_N(_03280_),
    .B1(_03284_),
    .B2(_03286_),
    .Y(_03294_));
 sky130_fd_sc_hd__o211ai_1 _13862_ (.A1(_03287_),
    .A2(_03288_),
    .B1(_03277_),
    .C1(_03280_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand3_4 _13863_ (.A(_03057_),
    .B(_03292_),
    .C(_03293_),
    .Y(_03296_));
 sky130_fd_sc_hd__a21oi_4 _13864_ (.A1(_03292_),
    .A2(_03293_),
    .B1(_03057_),
    .Y(_03297_));
 sky130_fd_sc_hd__nand3_2 _13865_ (.A(_03294_),
    .B(_03295_),
    .C(_03056_),
    .Y(_03298_));
 sky130_fd_sc_hd__o2bb2ai_2 _13866_ (.A1_N(_03296_),
    .A2_N(_03298_),
    .B1(_02610_),
    .B2(_03027_),
    .Y(_03299_));
 sky130_fd_sc_hd__a21o_1 _13867_ (.A1(_03296_),
    .A2(_03298_),
    .B1(_03029_),
    .X(_03300_));
 sky130_fd_sc_hd__o211ai_2 _13868_ (.A1(_03027_),
    .A2(_02610_),
    .B1(_03298_),
    .C1(_03296_),
    .Y(_03302_));
 sky130_fd_sc_hd__a31oi_4 _13869_ (.A1(_03057_),
    .A2(_03292_),
    .A3(_03293_),
    .B1(_03029_),
    .Y(_03303_));
 sky130_fd_sc_hd__nand2_2 _13870_ (.A(_03303_),
    .B(_03298_),
    .Y(_03304_));
 sky130_fd_sc_hd__nand3_1 _13871_ (.A(_03041_),
    .B(_03300_),
    .C(_03302_),
    .Y(_03305_));
 sky130_fd_sc_hd__and3_1 _13872_ (.A(_03299_),
    .B(_03304_),
    .C(_03040_),
    .X(_03306_));
 sky130_fd_sc_hd__nand3_1 _13873_ (.A(_03304_),
    .B(_03040_),
    .C(_03299_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand2_1 _13874_ (.A(_03305_),
    .B(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__a2bb2o_2 _13875_ (.A1_N(_02781_),
    .A2_N(_03042_),
    .B1(_03305_),
    .B2(_03307_),
    .X(_03309_));
 sky130_fd_sc_hd__a21oi_1 _13876_ (.A1(_03300_),
    .A2(_03302_),
    .B1(_03044_),
    .Y(_03310_));
 sky130_fd_sc_hd__a21o_2 _13877_ (.A1(_03300_),
    .A2(_03302_),
    .B1(_03044_),
    .X(_03311_));
 sky130_fd_sc_hd__a21oi_2 _13878_ (.A1(_03044_),
    .A2(_03308_),
    .B1(_03310_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _13879_ (.A(_03055_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__a21oi_1 _13880_ (.A1(_03309_),
    .A2(_03311_),
    .B1(_03055_),
    .Y(_03315_));
 sky130_fd_sc_hd__a21oi_1 _13881_ (.A1(_03055_),
    .A2(_03309_),
    .B1(_03315_),
    .Y(net79));
 sky130_fd_sc_hd__o2bb2a_1 _13882_ (.A1_N(_03105_),
    .A2_N(_03099_),
    .B1(_03097_),
    .B2(_03100_),
    .X(_03316_));
 sky130_fd_sc_hd__o21ai_2 _13883_ (.A1(_03097_),
    .A2(_03100_),
    .B1(_03107_),
    .Y(_03317_));
 sky130_fd_sc_hd__and2_1 _13884_ (.A(_03237_),
    .B(_03238_),
    .X(_03318_));
 sky130_fd_sc_hd__o21ai_1 _13885_ (.A1(_03238_),
    .A2(_03234_),
    .B1(_03237_),
    .Y(_03319_));
 sky130_fd_sc_hd__o21a_1 _13886_ (.A1(_03238_),
    .A2(_03234_),
    .B1(_03237_),
    .X(_03320_));
 sky130_fd_sc_hd__nand2_2 _13887_ (.A(net31),
    .B(net40),
    .Y(_03321_));
 sky130_fd_sc_hd__nand2_1 _13888_ (.A(net31),
    .B(net39),
    .Y(_03323_));
 sky130_fd_sc_hd__and4_1 _13889_ (.A(net30),
    .B(net31),
    .C(net39),
    .D(net40),
    .X(_03324_));
 sky130_fd_sc_hd__nand4_1 _13890_ (.A(net30),
    .B(net31),
    .C(net39),
    .D(net40),
    .Y(_03325_));
 sky130_fd_sc_hd__a22oi_2 _13891_ (.A1(net31),
    .A2(net39),
    .B1(net40),
    .B2(net30),
    .Y(_03326_));
 sky130_fd_sc_hd__a22o_1 _13892_ (.A1(net31),
    .A2(net39),
    .B1(net40),
    .B2(net30),
    .X(_03327_));
 sky130_fd_sc_hd__a2bb2oi_1 _13893_ (.A1_N(_01857_),
    .A2_N(_02010_),
    .B1(_03325_),
    .B2(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__o22ai_2 _13894_ (.A1(_01857_),
    .A2(_02010_),
    .B1(_03324_),
    .B2(_03326_),
    .Y(_03329_));
 sky130_fd_sc_hd__o2111a_1 _13895_ (.A1(_03088_),
    .A2(_03321_),
    .B1(net29),
    .C1(net41),
    .D1(_03327_),
    .X(_03330_));
 sky130_fd_sc_hd__o2111ai_2 _13896_ (.A1(_03088_),
    .A2(_03321_),
    .B1(net29),
    .C1(net41),
    .D1(_03327_),
    .Y(_03331_));
 sky130_fd_sc_hd__nand2_1 _13897_ (.A(_03329_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__o22ai_4 _13898_ (.A1(_03234_),
    .A2(_03318_),
    .B1(_03328_),
    .B2(_03330_),
    .Y(_03334_));
 sky130_fd_sc_hd__nand2_1 _13899_ (.A(_03329_),
    .B(_03319_),
    .Y(_03335_));
 sky130_fd_sc_hd__and3_2 _13900_ (.A(_03329_),
    .B(_03331_),
    .C(_03319_),
    .X(_03336_));
 sky130_fd_sc_hd__nand3_1 _13901_ (.A(_03329_),
    .B(_03331_),
    .C(_03319_),
    .Y(_03337_));
 sky130_fd_sc_hd__o21a_1 _13902_ (.A1(_01748_),
    .A2(_02010_),
    .B1(_03093_),
    .X(_03338_));
 sky130_fd_sc_hd__and3_1 _13903_ (.A(_03090_),
    .B(net41),
    .C(net28),
    .X(_03339_));
 sky130_fd_sc_hd__a31o_1 _13904_ (.A1(_03090_),
    .A2(net41),
    .A3(net28),
    .B1(_03091_),
    .X(_03340_));
 sky130_fd_sc_hd__a21oi_1 _13905_ (.A1(_03334_),
    .A2(_03337_),
    .B1(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__o2bb2ai_2 _13906_ (.A1_N(_03334_),
    .A2_N(_03337_),
    .B1(_03338_),
    .B2(_03089_),
    .Y(_03342_));
 sky130_fd_sc_hd__a21boi_2 _13907_ (.A1(_03332_),
    .A2(_03320_),
    .B1_N(_03340_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21ai_1 _13908_ (.A1(_03091_),
    .A2(_03339_),
    .B1(_03334_),
    .Y(_03345_));
 sky130_fd_sc_hd__o211a_1 _13909_ (.A1(_03091_),
    .A2(_03339_),
    .B1(_03337_),
    .C1(_03334_),
    .X(_03346_));
 sky130_fd_sc_hd__o21ai_2 _13910_ (.A1(_03341_),
    .A2(_03346_),
    .B1(_03316_),
    .Y(_03347_));
 sky130_fd_sc_hd__nand2_1 _13911_ (.A(_03317_),
    .B(_03342_),
    .Y(_03348_));
 sky130_fd_sc_hd__o211ai_4 _13912_ (.A1(_03336_),
    .A2(_03345_),
    .B1(_03342_),
    .C1(_03317_),
    .Y(_03349_));
 sky130_fd_sc_hd__a21oi_1 _13913_ (.A1(_02978_),
    .A2(_03069_),
    .B1(_03066_),
    .Y(_03350_));
 sky130_fd_sc_hd__a31o_1 _13914_ (.A1(_03070_),
    .A2(net45),
    .A3(net23),
    .B1(_03068_),
    .X(_03351_));
 sky130_fd_sc_hd__nand2_1 _13915_ (.A(net26),
    .B(net45),
    .Y(_03352_));
 sky130_fd_sc_hd__a22oi_1 _13916_ (.A1(net28),
    .A2(net42),
    .B1(net43),
    .B2(net27),
    .Y(_03353_));
 sky130_fd_sc_hd__a22o_2 _13917_ (.A1(net28),
    .A2(net42),
    .B1(net43),
    .B2(net27),
    .X(_03354_));
 sky130_fd_sc_hd__nand4_2 _13918_ (.A(net28),
    .B(net27),
    .C(net42),
    .D(net43),
    .Y(_03356_));
 sky130_fd_sc_hd__nand4_2 _13919_ (.A(_03354_),
    .B(_03356_),
    .C(net26),
    .D(net45),
    .Y(_03357_));
 sky130_fd_sc_hd__o2bb2ai_2 _13920_ (.A1_N(_03354_),
    .A2_N(_03356_),
    .B1(_01791_),
    .B2(_02054_),
    .Y(_03358_));
 sky130_fd_sc_hd__o211a_1 _13921_ (.A1(_03068_),
    .A2(_03350_),
    .B1(_03357_),
    .C1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__a21oi_4 _13922_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03351_),
    .Y(_03360_));
 sky130_fd_sc_hd__a22o_1 _13923_ (.A1(net23),
    .A2(net46),
    .B1(net47),
    .B2(net12),
    .X(_03361_));
 sky130_fd_sc_hd__and4_1 _13924_ (.A(net23),
    .B(net12),
    .C(net46),
    .D(net47),
    .X(_03362_));
 sky130_fd_sc_hd__nand4_2 _13925_ (.A(net23),
    .B(net12),
    .C(net46),
    .D(net47),
    .Y(_03363_));
 sky130_fd_sc_hd__and4_1 _13926_ (.A(_03361_),
    .B(_03363_),
    .C(net1),
    .D(net48),
    .X(_03364_));
 sky130_fd_sc_hd__nand4_1 _13927_ (.A(_03361_),
    .B(_03363_),
    .C(net1),
    .D(net48),
    .Y(_03365_));
 sky130_fd_sc_hd__o2bb2ai_1 _13928_ (.A1_N(_03361_),
    .A2_N(_03363_),
    .B1(_01846_),
    .B2(_02109_),
    .Y(_03367_));
 sky130_fd_sc_hd__nand2_1 _13929_ (.A(_03365_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__o21ai_2 _13930_ (.A1(_03359_),
    .A2(_03360_),
    .B1(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__a31o_1 _13931_ (.A1(_03351_),
    .A2(_03357_),
    .A3(_03358_),
    .B1(_03368_),
    .X(_03370_));
 sky130_fd_sc_hd__o21a_1 _13932_ (.A1(_03360_),
    .A2(_03370_),
    .B1(_03369_),
    .X(_03371_));
 sky130_fd_sc_hd__a21oi_1 _13933_ (.A1(_03347_),
    .A2(_03349_),
    .B1(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__a21o_1 _13934_ (.A1(_03347_),
    .A2(_03349_),
    .B1(_03371_),
    .X(_03373_));
 sky130_fd_sc_hd__o211a_1 _13935_ (.A1(_03346_),
    .A2(_03348_),
    .B1(_03347_),
    .C1(_03371_),
    .X(_03374_));
 sky130_fd_sc_hd__o2111ai_4 _13936_ (.A1(_03360_),
    .A2(_03370_),
    .B1(_03369_),
    .C1(_03347_),
    .D1(_03349_),
    .Y(_03375_));
 sky130_fd_sc_hd__nand2_1 _13937_ (.A(_03373_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__a21oi_2 _13938_ (.A1(_03249_),
    .A2(_03253_),
    .B1(_03250_),
    .Y(_03378_));
 sky130_fd_sc_hd__o21ai_2 _13939_ (.A1(_03372_),
    .A2(_03374_),
    .B1(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__o211ai_4 _13940_ (.A1(_03250_),
    .A2(_03256_),
    .B1(_03373_),
    .C1(_03375_),
    .Y(_03380_));
 sky130_fd_sc_hd__inv_2 _13941_ (.A(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__a21o_1 _13942_ (.A1(_03110_),
    .A2(_03083_),
    .B1(_03111_),
    .X(_03382_));
 sky130_fd_sc_hd__a21oi_1 _13943_ (.A1(_03379_),
    .A2(_03380_),
    .B1(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__a21o_2 _13944_ (.A1(_03379_),
    .A2(_03380_),
    .B1(_03382_),
    .X(_03384_));
 sky130_fd_sc_hd__a22oi_4 _13945_ (.A1(_03112_),
    .A2(_03115_),
    .B1(_03376_),
    .B2(_03378_),
    .Y(_03385_));
 sky130_fd_sc_hd__nand2_1 _13946_ (.A(_03379_),
    .B(_03382_),
    .Y(_03386_));
 sky130_fd_sc_hd__and3_1 _13947_ (.A(_03379_),
    .B(_03380_),
    .C(_03382_),
    .X(_03387_));
 sky130_fd_sc_hd__nand3_2 _13948_ (.A(_03379_),
    .B(_03380_),
    .C(_03382_),
    .Y(_03389_));
 sky130_fd_sc_hd__a21oi_1 _13949_ (.A1(_03380_),
    .A2(_03385_),
    .B1(_03383_),
    .Y(_03390_));
 sky130_fd_sc_hd__o21a_1 _13950_ (.A1(_03243_),
    .A2(_03232_),
    .B1(_03231_),
    .X(_03391_));
 sky130_fd_sc_hd__o21ai_2 _13951_ (.A1(_03243_),
    .A2(_03232_),
    .B1(_03231_),
    .Y(_03392_));
 sky130_fd_sc_hd__a21oi_4 _13952_ (.A1(_03179_),
    .A2(_03196_),
    .B1(_03194_),
    .Y(_03393_));
 sky130_fd_sc_hd__a32o_1 _13953_ (.A1(_03181_),
    .A2(_03192_),
    .A3(_03193_),
    .B1(_03196_),
    .B2(_03179_),
    .X(_03394_));
 sky130_fd_sc_hd__a22oi_4 _13954_ (.A1(net3),
    .A2(net36),
    .B1(net37),
    .B2(net2),
    .Y(_03395_));
 sky130_fd_sc_hd__and4_1 _13955_ (.A(net2),
    .B(net3),
    .C(net36),
    .D(net37),
    .X(_03396_));
 sky130_fd_sc_hd__nand4_1 _13956_ (.A(net2),
    .B(net3),
    .C(net36),
    .D(net37),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _13957_ (.A(net32),
    .B(net38),
    .Y(_03398_));
 sky130_fd_sc_hd__o2bb2a_1 _13958_ (.A1_N(net32),
    .A2_N(net38),
    .B1(_03395_),
    .B2(_03396_),
    .X(_03400_));
 sky130_fd_sc_hd__and4b_1 _13959_ (.A_N(_03395_),
    .B(_03397_),
    .C(net32),
    .D(net38),
    .X(_03401_));
 sky130_fd_sc_hd__o211a_1 _13960_ (.A1(_03395_),
    .A2(_03396_),
    .B1(net32),
    .C1(net38),
    .X(_03402_));
 sky130_fd_sc_hd__o211ai_1 _13961_ (.A1(_03395_),
    .A2(_03396_),
    .B1(net32),
    .C1(net38),
    .Y(_03403_));
 sky130_fd_sc_hd__a211oi_2 _13962_ (.A1(net32),
    .A2(net38),
    .B1(_03395_),
    .C1(_03396_),
    .Y(_03404_));
 sky130_fd_sc_hd__a211o_1 _13963_ (.A1(net32),
    .A2(net38),
    .B1(_03395_),
    .C1(_03396_),
    .X(_03405_));
 sky130_fd_sc_hd__o21ai_2 _13964_ (.A1(_03221_),
    .A2(_03225_),
    .B1(_03223_),
    .Y(_03406_));
 sky130_fd_sc_hd__nand2_1 _13965_ (.A(net35),
    .B(net4),
    .Y(_03407_));
 sky130_fd_sc_hd__and4_2 _13966_ (.A(net64),
    .B(net34),
    .C(net5),
    .D(net6),
    .X(_03408_));
 sky130_fd_sc_hd__nand4_2 _13967_ (.A(net64),
    .B(net34),
    .C(net5),
    .D(net6),
    .Y(_03409_));
 sky130_fd_sc_hd__a22oi_4 _13968_ (.A1(net34),
    .A2(net5),
    .B1(net6),
    .B2(net64),
    .Y(_03411_));
 sky130_fd_sc_hd__a22o_1 _13969_ (.A1(net34),
    .A2(net5),
    .B1(net6),
    .B2(net64),
    .X(_03412_));
 sky130_fd_sc_hd__o211ai_2 _13970_ (.A1(_01934_),
    .A2(_01945_),
    .B1(_03409_),
    .C1(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__o21bai_2 _13971_ (.A1(_03408_),
    .A2(_03411_),
    .B1_N(_03407_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand4_2 _13972_ (.A(_03412_),
    .B(net4),
    .C(net35),
    .D(_03409_),
    .Y(_03415_));
 sky130_fd_sc_hd__o22ai_4 _13973_ (.A1(_01934_),
    .A2(_01945_),
    .B1(_03408_),
    .B2(_03411_),
    .Y(_03416_));
 sky130_fd_sc_hd__and3_1 _13974_ (.A(_03416_),
    .B(_03406_),
    .C(_03415_),
    .X(_03417_));
 sky130_fd_sc_hd__nand3_4 _13975_ (.A(_03416_),
    .B(_03406_),
    .C(_03415_),
    .Y(_03418_));
 sky130_fd_sc_hd__a21oi_1 _13976_ (.A1(_03415_),
    .A2(_03416_),
    .B1(_03406_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand3b_4 _13977_ (.A_N(_03406_),
    .B(_03413_),
    .C(_03414_),
    .Y(_03420_));
 sky130_fd_sc_hd__o211ai_4 _13978_ (.A1(_03400_),
    .A2(_03401_),
    .B1(_03418_),
    .C1(_03420_),
    .Y(_03422_));
 sky130_fd_sc_hd__a22o_2 _13979_ (.A1(_03403_),
    .A2(_03405_),
    .B1(_03418_),
    .B2(_03420_),
    .X(_03423_));
 sky130_fd_sc_hd__o21ai_4 _13980_ (.A1(_03402_),
    .A2(_03404_),
    .B1(_03420_),
    .Y(_03424_));
 sky130_fd_sc_hd__o211ai_1 _13981_ (.A1(_03402_),
    .A2(_03404_),
    .B1(_03418_),
    .C1(_03420_),
    .Y(_03425_));
 sky130_fd_sc_hd__a2bb2o_1 _13982_ (.A1_N(_03400_),
    .A2_N(_03401_),
    .B1(_03418_),
    .B2(_03420_),
    .X(_03426_));
 sky130_fd_sc_hd__o221a_2 _13983_ (.A1(_03417_),
    .A2(_03424_),
    .B1(_03194_),
    .B2(_03197_),
    .C1(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__o221ai_4 _13984_ (.A1(_03417_),
    .A2(_03424_),
    .B1(_03194_),
    .B2(_03197_),
    .C1(_03426_),
    .Y(_03428_));
 sky130_fd_sc_hd__nand3_4 _13985_ (.A(_03423_),
    .B(_03393_),
    .C(_03422_),
    .Y(_03429_));
 sky130_fd_sc_hd__a31o_1 _13986_ (.A1(_03394_),
    .A2(_03425_),
    .A3(_03426_),
    .B1(_03392_),
    .X(_03430_));
 sky130_fd_sc_hd__a31oi_4 _13987_ (.A1(_03423_),
    .A2(_03393_),
    .A3(_03422_),
    .B1(_03391_),
    .Y(_03431_));
 sky130_fd_sc_hd__a31o_1 _13988_ (.A1(_03423_),
    .A2(_03393_),
    .A3(_03422_),
    .B1(_03391_),
    .X(_03433_));
 sky130_fd_sc_hd__and3_1 _13989_ (.A(_03428_),
    .B(_03429_),
    .C(_03391_),
    .X(_03434_));
 sky130_fd_sc_hd__a21oi_2 _13990_ (.A1(_03428_),
    .A2(_03429_),
    .B1(_03391_),
    .Y(_03435_));
 sky130_fd_sc_hd__a21oi_2 _13991_ (.A1(_03428_),
    .A2(_03429_),
    .B1(_03392_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21o_1 _13992_ (.A1(_03428_),
    .A2(_03429_),
    .B1(_03392_),
    .X(_03437_));
 sky130_fd_sc_hd__and3_1 _13993_ (.A(_03392_),
    .B(_03428_),
    .C(_03429_),
    .X(_03438_));
 sky130_fd_sc_hd__o21ai_2 _13994_ (.A1(_03427_),
    .A2(_03433_),
    .B1(_03437_),
    .Y(_03439_));
 sky130_fd_sc_hd__o21ai_1 _13995_ (.A1(_01780_),
    .A2(_02043_),
    .B1(_03139_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21ai_2 _13996_ (.A1(_03134_),
    .A2(_03135_),
    .B1(_03139_),
    .Y(_03441_));
 sky130_fd_sc_hd__o21a_1 _13997_ (.A1(_03134_),
    .A2(_03135_),
    .B1(_03139_),
    .X(_03442_));
 sky130_fd_sc_hd__nand2_1 _13998_ (.A(net55),
    .B(net14),
    .Y(_03444_));
 sky130_fd_sc_hd__a22oi_4 _13999_ (.A1(net44),
    .A2(net15),
    .B1(net16),
    .B2(net33),
    .Y(_03445_));
 sky130_fd_sc_hd__a22o_2 _14000_ (.A1(net44),
    .A2(net15),
    .B1(net16),
    .B2(net33),
    .X(_03446_));
 sky130_fd_sc_hd__and4_1 _14001_ (.A(net33),
    .B(net44),
    .C(net15),
    .D(net16),
    .X(_03447_));
 sky130_fd_sc_hd__nand4_4 _14002_ (.A(net33),
    .B(net44),
    .C(net15),
    .D(net16),
    .Y(_03448_));
 sky130_fd_sc_hd__o211ai_2 _14003_ (.A1(_01780_),
    .A2(_02065_),
    .B1(_03446_),
    .C1(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__o21bai_1 _14004_ (.A1(_03445_),
    .A2(_03447_),
    .B1_N(_03444_),
    .Y(_03450_));
 sky130_fd_sc_hd__o22ai_4 _14005_ (.A1(_01780_),
    .A2(_02065_),
    .B1(_03445_),
    .B2(_03447_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand4_4 _14006_ (.A(_03446_),
    .B(_03448_),
    .C(net55),
    .D(net14),
    .Y(_03452_));
 sky130_fd_sc_hd__a22oi_1 _14007_ (.A1(_03137_),
    .A2(_03440_),
    .B1(_03451_),
    .B2(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand3_4 _14008_ (.A(_03442_),
    .B(_03449_),
    .C(_03450_),
    .Y(_03455_));
 sky130_fd_sc_hd__o31a_1 _14009_ (.A1(_03444_),
    .A2(_03445_),
    .A3(_03447_),
    .B1(_03441_),
    .X(_03456_));
 sky130_fd_sc_hd__nand3_4 _14010_ (.A(_03451_),
    .B(_03452_),
    .C(_03441_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_1 _14011_ (.A(net60),
    .B(net10),
    .Y(_03458_));
 sky130_fd_sc_hd__nand2_2 _14012_ (.A(net58),
    .B(net13),
    .Y(_03459_));
 sky130_fd_sc_hd__a22oi_4 _14013_ (.A1(net59),
    .A2(net11),
    .B1(net13),
    .B2(net58),
    .Y(_03460_));
 sky130_fd_sc_hd__a22o_1 _14014_ (.A1(net59),
    .A2(net11),
    .B1(net13),
    .B2(net58),
    .X(_03461_));
 sky130_fd_sc_hd__and4_1 _14015_ (.A(net58),
    .B(net59),
    .C(net11),
    .D(net13),
    .X(_03462_));
 sky130_fd_sc_hd__nand4_2 _14016_ (.A(net58),
    .B(net59),
    .C(net11),
    .D(net13),
    .Y(_03463_));
 sky130_fd_sc_hd__and3_1 _14017_ (.A(_03458_),
    .B(_03461_),
    .C(_03463_),
    .X(_03464_));
 sky130_fd_sc_hd__o211ai_2 _14018_ (.A1(_01835_),
    .A2(_02021_),
    .B1(_03461_),
    .C1(_03463_),
    .Y(_03466_));
 sky130_fd_sc_hd__o211a_1 _14019_ (.A1(_03460_),
    .A2(_03462_),
    .B1(net60),
    .C1(net10),
    .X(_03467_));
 sky130_fd_sc_hd__o21bai_2 _14020_ (.A1(_03460_),
    .A2(_03462_),
    .B1_N(_03458_),
    .Y(_03468_));
 sky130_fd_sc_hd__o22a_1 _14021_ (.A1(_01835_),
    .A2(_02021_),
    .B1(_03460_),
    .B2(_03462_),
    .X(_03469_));
 sky130_fd_sc_hd__o21ai_2 _14022_ (.A1(_03460_),
    .A2(_03462_),
    .B1(_03458_),
    .Y(_03470_));
 sky130_fd_sc_hd__a41o_1 _14023_ (.A1(net58),
    .A2(net59),
    .A3(net11),
    .A4(net13),
    .B1(_03458_),
    .X(_03471_));
 sky130_fd_sc_hd__and4_1 _14024_ (.A(_03461_),
    .B(_03463_),
    .C(net60),
    .D(net10),
    .X(_03472_));
 sky130_fd_sc_hd__o21ai_1 _14025_ (.A1(_03460_),
    .A2(_03471_),
    .B1(_03470_),
    .Y(_03473_));
 sky130_fd_sc_hd__nand2_1 _14026_ (.A(_03466_),
    .B(_03468_),
    .Y(_03474_));
 sky130_fd_sc_hd__o2bb2ai_4 _14027_ (.A1_N(_03455_),
    .A2_N(_03457_),
    .B1(_03464_),
    .B2(_03467_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand4_4 _14028_ (.A(_03455_),
    .B(_03457_),
    .C(_03466_),
    .D(_03468_),
    .Y(_03477_));
 sky130_fd_sc_hd__o2bb2ai_1 _14029_ (.A1_N(_03455_),
    .A2_N(_03457_),
    .B1(_03469_),
    .B2(_03472_),
    .Y(_03478_));
 sky130_fd_sc_hd__o2111ai_4 _14030_ (.A1(_03460_),
    .A2(_03471_),
    .B1(_03470_),
    .C1(_03455_),
    .D1(_03457_),
    .Y(_03479_));
 sky130_fd_sc_hd__a32oi_4 _14031_ (.A1(_03132_),
    .A2(_03142_),
    .A3(_03145_),
    .B1(_03148_),
    .B2(_03165_),
    .Y(_03480_));
 sky130_fd_sc_hd__o22ai_2 _14032_ (.A1(_03144_),
    .A2(_03149_),
    .B1(_03164_),
    .B2(_03146_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand3_4 _14033_ (.A(_03475_),
    .B(_03480_),
    .C(_03477_),
    .Y(_03482_));
 sky130_fd_sc_hd__a21oi_4 _14034_ (.A1(_03475_),
    .A2(_03477_),
    .B1(_03480_),
    .Y(_03483_));
 sky130_fd_sc_hd__nand3_4 _14035_ (.A(_03478_),
    .B(_03479_),
    .C(_03481_),
    .Y(_03484_));
 sky130_fd_sc_hd__nand2_1 _14036_ (.A(_03482_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__o21ai_2 _14037_ (.A1(_02857_),
    .A2(_03184_),
    .B1(_03183_),
    .Y(_03486_));
 sky130_fd_sc_hd__a22o_1 _14038_ (.A1(_03183_),
    .A2(_03185_),
    .B1(_03186_),
    .B2(_02856_),
    .X(_03488_));
 sky130_fd_sc_hd__nor2_1 _14039_ (.A(_03152_),
    .B(_03153_),
    .Y(_03489_));
 sky130_fd_sc_hd__o21a_1 _14040_ (.A1(_03152_),
    .A2(_03153_),
    .B1(_03156_),
    .X(_03490_));
 sky130_fd_sc_hd__nand2_2 _14041_ (.A(net62),
    .B(net9),
    .Y(_03491_));
 sky130_fd_sc_hd__and4_1 _14042_ (.A(net61),
    .B(net62),
    .C(net8),
    .D(net9),
    .X(_03492_));
 sky130_fd_sc_hd__nand2_1 _14043_ (.A(net61),
    .B(net9),
    .Y(_03493_));
 sky130_fd_sc_hd__a22o_2 _14044_ (.A1(net62),
    .A2(net8),
    .B1(net9),
    .B2(net61),
    .X(_03494_));
 sky130_fd_sc_hd__o2bb2ai_1 _14045_ (.A1_N(_03184_),
    .A2_N(_03493_),
    .B1(_03491_),
    .B2(_03186_),
    .Y(_03495_));
 sky130_fd_sc_hd__o221ai_4 _14046_ (.A1(_01890_),
    .A2(_01977_),
    .B1(_03186_),
    .B2(_03491_),
    .C1(_03494_),
    .Y(_03496_));
 sky130_fd_sc_hd__nand3_2 _14047_ (.A(_03495_),
    .B(net7),
    .C(net63),
    .Y(_03497_));
 sky130_fd_sc_hd__o2111ai_4 _14048_ (.A1(_03186_),
    .A2(_03491_),
    .B1(net63),
    .C1(net7),
    .D1(_03494_),
    .Y(_03499_));
 sky130_fd_sc_hd__o21ai_2 _14049_ (.A1(_01890_),
    .A2(_01977_),
    .B1(_03495_),
    .Y(_03500_));
 sky130_fd_sc_hd__o211a_1 _14050_ (.A1(_03155_),
    .A2(_03489_),
    .B1(_03499_),
    .C1(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__o211ai_4 _14051_ (.A1(_03155_),
    .A2(_03489_),
    .B1(_03499_),
    .C1(_03500_),
    .Y(_03502_));
 sky130_fd_sc_hd__nand3_2 _14052_ (.A(_03490_),
    .B(_03496_),
    .C(_03497_),
    .Y(_03503_));
 sky130_fd_sc_hd__a31oi_4 _14053_ (.A1(_03490_),
    .A2(_03496_),
    .A3(_03497_),
    .B1(_03488_),
    .Y(_03504_));
 sky130_fd_sc_hd__and3b_2 _14054_ (.A_N(_03488_),
    .B(_03502_),
    .C(_03503_),
    .X(_03505_));
 sky130_fd_sc_hd__a22oi_4 _14055_ (.A1(_03187_),
    .A2(_03486_),
    .B1(_03502_),
    .B2(_03503_),
    .Y(_03506_));
 sky130_fd_sc_hd__a21oi_4 _14056_ (.A1(_03502_),
    .A2(_03504_),
    .B1(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__nand2_2 _14057_ (.A(_03485_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__o211ai_4 _14058_ (.A1(_03505_),
    .A2(_03506_),
    .B1(_03482_),
    .C1(_03484_),
    .Y(_03510_));
 sky130_fd_sc_hd__o2bb2ai_4 _14059_ (.A1_N(_03482_),
    .A2_N(_03484_),
    .B1(_03505_),
    .B2(_03506_),
    .Y(_03511_));
 sky130_fd_sc_hd__a311oi_2 _14060_ (.A1(_03475_),
    .A2(_03480_),
    .A3(_03477_),
    .B1(_03506_),
    .C1(_03505_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_2 _14061_ (.A(_03507_),
    .B(_03482_),
    .Y(_03513_));
 sky130_fd_sc_hd__and3_1 _14062_ (.A(_03482_),
    .B(_03507_),
    .C(_03484_),
    .X(_03514_));
 sky130_fd_sc_hd__nand3_1 _14063_ (.A(_03507_),
    .B(_03484_),
    .C(_03482_),
    .Y(_03515_));
 sky130_fd_sc_hd__o32ai_4 _14064_ (.A1(_03168_),
    .A2(_03171_),
    .A3(_03173_),
    .B1(_03204_),
    .B2(_03176_),
    .Y(_03516_));
 sky130_fd_sc_hd__a21oi_4 _14065_ (.A1(_03511_),
    .A2(_03515_),
    .B1(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__o2111ai_4 _14066_ (.A1(_03204_),
    .A2(_03176_),
    .B1(_03175_),
    .C1(_03510_),
    .D1(_03508_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2_1 _14067_ (.A(_03511_),
    .B(_03516_),
    .Y(_03519_));
 sky130_fd_sc_hd__a22oi_4 _14068_ (.A1(_03175_),
    .A2(_03209_),
    .B1(_03508_),
    .B2(_03510_),
    .Y(_03521_));
 sky130_fd_sc_hd__o211ai_4 _14069_ (.A1(_03513_),
    .A2(_03483_),
    .B1(_03511_),
    .C1(_03516_),
    .Y(_03522_));
 sky130_fd_sc_hd__o22ai_4 _14070_ (.A1(_03514_),
    .A2(_03519_),
    .B1(_03517_),
    .B2(_03439_),
    .Y(_03523_));
 sky130_fd_sc_hd__o211ai_2 _14071_ (.A1(_03436_),
    .A2(_03438_),
    .B1(_03518_),
    .C1(_03522_),
    .Y(_03524_));
 sky130_fd_sc_hd__o22ai_2 _14072_ (.A1(_03434_),
    .A2(_03435_),
    .B1(_03517_),
    .B2(_03521_),
    .Y(_03525_));
 sky130_fd_sc_hd__o22ai_4 _14073_ (.A1(_03436_),
    .A2(_03438_),
    .B1(_03517_),
    .B2(_03521_),
    .Y(_03526_));
 sky130_fd_sc_hd__o211ai_4 _14074_ (.A1(_03434_),
    .A2(_03435_),
    .B1(_03518_),
    .C1(_03522_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _14075_ (.A(_03526_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__o21ai_1 _14076_ (.A1(_03254_),
    .A2(_03259_),
    .B1(_03216_),
    .Y(_03529_));
 sky130_fd_sc_hd__o22ai_4 _14077_ (.A1(_03211_),
    .A2(_03214_),
    .B1(_03217_),
    .B2(_03261_),
    .Y(_03530_));
 sky130_fd_sc_hd__o31ai_4 _14078_ (.A1(_03129_),
    .A2(_03205_),
    .A3(_03207_),
    .B1(_03529_),
    .Y(_03532_));
 sky130_fd_sc_hd__and3_1 _14079_ (.A(_03524_),
    .B(_03525_),
    .C(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__nand3_4 _14080_ (.A(_03524_),
    .B(_03525_),
    .C(_03532_),
    .Y(_03534_));
 sky130_fd_sc_hd__and3_2 _14081_ (.A(_03526_),
    .B(_03530_),
    .C(_03527_),
    .X(_03535_));
 sky130_fd_sc_hd__nand3_4 _14082_ (.A(_03526_),
    .B(_03530_),
    .C(_03527_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _14083_ (.A(_03534_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__a22o_2 _14084_ (.A1(_03384_),
    .A2(_03389_),
    .B1(_03534_),
    .B2(_03536_),
    .X(_03538_));
 sky130_fd_sc_hd__o211a_1 _14085_ (.A1(_03386_),
    .A2(_03381_),
    .B1(_03384_),
    .C1(_03534_),
    .X(_03539_));
 sky130_fd_sc_hd__o211ai_4 _14086_ (.A1(_03386_),
    .A2(_03381_),
    .B1(_03384_),
    .C1(_03534_),
    .Y(_03540_));
 sky130_fd_sc_hd__nand4_2 _14087_ (.A(_03384_),
    .B(_03389_),
    .C(_03534_),
    .D(_03536_),
    .Y(_03541_));
 sky130_fd_sc_hd__o211ai_2 _14088_ (.A1(_03383_),
    .A2(_03387_),
    .B1(_03534_),
    .C1(_03536_),
    .Y(_03543_));
 sky130_fd_sc_hd__nand2_1 _14089_ (.A(_03537_),
    .B(_03390_),
    .Y(_03544_));
 sky130_fd_sc_hd__o22ai_4 _14090_ (.A1(_03265_),
    .A2(_03269_),
    .B1(_03266_),
    .B2(_03126_),
    .Y(_03545_));
 sky130_fd_sc_hd__o211ai_4 _14091_ (.A1(_03535_),
    .A2(_03540_),
    .B1(_03545_),
    .C1(_03538_),
    .Y(_03546_));
 sky130_fd_sc_hd__a21oi_1 _14092_ (.A1(_03538_),
    .A2(_03541_),
    .B1(_03545_),
    .Y(_03547_));
 sky130_fd_sc_hd__o2111ai_4 _14093_ (.A1(_03126_),
    .A2(_03266_),
    .B1(_03271_),
    .C1(_03543_),
    .D1(_03544_),
    .Y(_03548_));
 sky130_fd_sc_hd__and4b_2 _14094_ (.A_N(_03063_),
    .B(_03065_),
    .C(_03074_),
    .D(_03075_),
    .X(_03549_));
 sky130_fd_sc_hd__a31o_1 _14095_ (.A1(_03063_),
    .A2(_03076_),
    .A3(_03080_),
    .B1(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__o21ai_2 _14096_ (.A1(_03116_),
    .A2(_03117_),
    .B1(_03123_),
    .Y(_03551_));
 sky130_fd_sc_hd__inv_2 _14097_ (.A(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__and2b_2 _14098_ (.A_N(_03550_),
    .B(_03551_),
    .X(_03554_));
 sky130_fd_sc_hd__a311o_1 _14099_ (.A1(_03063_),
    .A2(_03076_),
    .A3(_03080_),
    .B1(_03549_),
    .C1(_03552_),
    .X(_03555_));
 sky130_fd_sc_hd__o211a_1 _14100_ (.A1(_03117_),
    .A2(_03116_),
    .B1(_03550_),
    .C1(_03123_),
    .X(_03556_));
 sky130_fd_sc_hd__and2_1 _14101_ (.A(_03550_),
    .B(_03551_),
    .X(_03557_));
 sky130_fd_sc_hd__nor2_1 _14102_ (.A(_03550_),
    .B(_03551_),
    .Y(_03558_));
 sky130_fd_sc_hd__nor2_2 _14103_ (.A(_03554_),
    .B(_03556_),
    .Y(_03559_));
 sky130_fd_sc_hd__nor2_1 _14104_ (.A(_03557_),
    .B(_03558_),
    .Y(_03560_));
 sky130_fd_sc_hd__a21oi_2 _14105_ (.A1(_03546_),
    .A2(_03548_),
    .B1(_03559_),
    .Y(_03561_));
 sky130_fd_sc_hd__o2bb2ai_2 _14106_ (.A1_N(_03546_),
    .A2_N(_03548_),
    .B1(_03554_),
    .B2(_03556_),
    .Y(_03562_));
 sky130_fd_sc_hd__and3_1 _14107_ (.A(_03546_),
    .B(_03548_),
    .C(_03559_),
    .X(_03563_));
 sky130_fd_sc_hd__o211ai_2 _14108_ (.A1(_03557_),
    .A2(_03558_),
    .B1(_03546_),
    .C1(_03548_),
    .Y(_03565_));
 sky130_fd_sc_hd__o2bb2ai_1 _14109_ (.A1_N(_03546_),
    .A2_N(_03548_),
    .B1(_03557_),
    .B2(_03558_),
    .Y(_03566_));
 sky130_fd_sc_hd__o211ai_2 _14110_ (.A1(_03554_),
    .A2(_03556_),
    .B1(_03546_),
    .C1(_03548_),
    .Y(_03567_));
 sky130_fd_sc_hd__a31oi_2 _14111_ (.A1(_03059_),
    .A2(_03273_),
    .A3(_03274_),
    .B1(_03289_),
    .Y(_03568_));
 sky130_fd_sc_hd__a32oi_4 _14112_ (.A1(_03058_),
    .A2(_03275_),
    .A3(_03276_),
    .B1(_03277_),
    .B2(_03291_),
    .Y(_03569_));
 sky130_fd_sc_hd__a32o_1 _14113_ (.A1(_03058_),
    .A2(_03275_),
    .A3(_03276_),
    .B1(_03277_),
    .B2(_03291_),
    .X(_03570_));
 sky130_fd_sc_hd__a21oi_2 _14114_ (.A1(_03562_),
    .A2(_03565_),
    .B1(_03569_),
    .Y(_03571_));
 sky130_fd_sc_hd__o211ai_4 _14115_ (.A1(_03278_),
    .A2(_03568_),
    .B1(_03567_),
    .C1(_03566_),
    .Y(_03572_));
 sky130_fd_sc_hd__and3_1 _14116_ (.A(_03562_),
    .B(_03569_),
    .C(_03565_),
    .X(_03573_));
 sky130_fd_sc_hd__nand3_2 _14117_ (.A(_03562_),
    .B(_03569_),
    .C(_03565_),
    .Y(_03574_));
 sky130_fd_sc_hd__a21o_1 _14118_ (.A1(_03572_),
    .A2(_03574_),
    .B1(_03285_),
    .X(_03576_));
 sky130_fd_sc_hd__o211ai_2 _14119_ (.A1(_03283_),
    .A2(_03281_),
    .B1(_03574_),
    .C1(_03572_),
    .Y(_03577_));
 sky130_fd_sc_hd__o2bb2ai_2 _14120_ (.A1_N(_03572_),
    .A2_N(_03574_),
    .B1(_03281_),
    .B2(_03283_),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_2 _14121_ (.A(_03572_),
    .B(_03284_),
    .Y(_03579_));
 sky130_fd_sc_hd__o21ai_2 _14122_ (.A1(_03573_),
    .A2(_03579_),
    .B1(_03578_),
    .Y(_03580_));
 sky130_fd_sc_hd__a21oi_4 _14123_ (.A1(_03296_),
    .A2(_03030_),
    .B1(_03297_),
    .Y(_03581_));
 sky130_fd_sc_hd__nand3_4 _14124_ (.A(_03576_),
    .B(_03577_),
    .C(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__o221a_1 _14125_ (.A1(_03297_),
    .A2(_03303_),
    .B1(_03573_),
    .B2(_03579_),
    .C1(_03578_),
    .X(_03583_));
 sky130_fd_sc_hd__o221ai_4 _14126_ (.A1(_03297_),
    .A2(_03303_),
    .B1(_03573_),
    .B2(_03579_),
    .C1(_03578_),
    .Y(_03584_));
 sky130_fd_sc_hd__a32oi_4 _14127_ (.A1(_03040_),
    .A2(_03299_),
    .A3(_03304_),
    .B1(_03582_),
    .B2(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__a32o_1 _14128_ (.A1(_03040_),
    .A2(_03299_),
    .A3(_03304_),
    .B1(_03582_),
    .B2(_03584_),
    .X(_03587_));
 sky130_fd_sc_hd__a21o_1 _14129_ (.A1(_03580_),
    .A2(_03581_),
    .B1(_03307_),
    .X(_03588_));
 sky130_fd_sc_hd__a21oi_4 _14130_ (.A1(_03306_),
    .A2(_03582_),
    .B1(_03585_),
    .Y(_03589_));
 sky130_fd_sc_hd__and3_1 _14131_ (.A(_03311_),
    .B(_03314_),
    .C(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__a21oi_1 _14132_ (.A1(_03311_),
    .A2(_03314_),
    .B1(_03589_),
    .Y(_03591_));
 sky130_fd_sc_hd__or2_1 _14133_ (.A(_03590_),
    .B(_03591_),
    .X(net80));
 sky130_fd_sc_hd__o31a_1 _14134_ (.A1(_03372_),
    .A2(_03374_),
    .A3(_03378_),
    .B1(_03386_),
    .X(_03592_));
 sky130_fd_sc_hd__o21bai_2 _14135_ (.A1(_03368_),
    .A2(_03360_),
    .B1_N(_03359_),
    .Y(_03593_));
 sky130_fd_sc_hd__nor2_2 _14136_ (.A(_01846_),
    .B(_02120_),
    .Y(_03594_));
 sky130_fd_sc_hd__a31o_1 _14137_ (.A1(_03361_),
    .A2(net48),
    .A3(net1),
    .B1(_03362_),
    .X(_03595_));
 sky130_fd_sc_hd__a211o_1 _14138_ (.A1(_03363_),
    .A2(_03365_),
    .B1(_01846_),
    .C1(_02120_),
    .X(_03596_));
 sky130_fd_sc_hd__a211o_1 _14139_ (.A1(net1),
    .A2(net49),
    .B1(_03362_),
    .C1(_03364_),
    .X(_03597_));
 sky130_fd_sc_hd__nand2_1 _14140_ (.A(_03596_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__and3_2 _14141_ (.A(_03593_),
    .B(_03596_),
    .C(_03597_),
    .X(_03599_));
 sky130_fd_sc_hd__xor2_2 _14142_ (.A(_03593_),
    .B(_03598_),
    .X(_03600_));
 sky130_fd_sc_hd__inv_2 _14143_ (.A(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__nor4_2 _14144_ (.A(_02989_),
    .B(_03062_),
    .C(_03076_),
    .D(_03600_),
    .Y(_03602_));
 sky130_fd_sc_hd__o31a_1 _14145_ (.A1(_02989_),
    .A2(_03062_),
    .A3(_03076_),
    .B1(_03600_),
    .X(_03603_));
 sky130_fd_sc_hd__nor2_1 _14146_ (.A(_03602_),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__or2_1 _14147_ (.A(_03602_),
    .B(_03603_),
    .X(_03605_));
 sky130_fd_sc_hd__o21ai_2 _14148_ (.A1(_03602_),
    .A2(_03603_),
    .B1(_03592_),
    .Y(_03607_));
 sky130_fd_sc_hd__inv_2 _14149_ (.A(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21a_2 _14150_ (.A1(_03381_),
    .A2(_03385_),
    .B1(_03604_),
    .X(_03609_));
 sky130_fd_sc_hd__o21ai_4 _14151_ (.A1(_03381_),
    .A2(_03385_),
    .B1(_03604_),
    .Y(_03610_));
 sky130_fd_sc_hd__and2_1 _14152_ (.A(_03607_),
    .B(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__nand2_1 _14153_ (.A(_03607_),
    .B(_03610_),
    .Y(_03612_));
 sky130_fd_sc_hd__a32oi_4 _14154_ (.A1(_03526_),
    .A2(_03530_),
    .A3(_03527_),
    .B1(_03384_),
    .B2(_03389_),
    .Y(_03613_));
 sky130_fd_sc_hd__o21ai_1 _14155_ (.A1(_03383_),
    .A2(_03387_),
    .B1(_03536_),
    .Y(_03614_));
 sky130_fd_sc_hd__o21ai_1 _14156_ (.A1(_03528_),
    .A2(_03532_),
    .B1(_03540_),
    .Y(_03615_));
 sky130_fd_sc_hd__o2bb2ai_1 _14157_ (.A1_N(_03340_),
    .A2_N(_03334_),
    .B1(_03330_),
    .B2(_03335_),
    .Y(_03616_));
 sky130_fd_sc_hd__and2_1 _14158_ (.A(_03397_),
    .B(_03398_),
    .X(_03618_));
 sky130_fd_sc_hd__o21ai_1 _14159_ (.A1(_03398_),
    .A2(_03395_),
    .B1(_03397_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand2_1 _14160_ (.A(net32),
    .B(net40),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_1 _14161_ (.A(net32),
    .B(net39),
    .Y(_03621_));
 sky130_fd_sc_hd__and4_2 _14162_ (.A(net31),
    .B(net32),
    .C(net39),
    .D(net40),
    .X(_03622_));
 sky130_fd_sc_hd__nand4_1 _14163_ (.A(net31),
    .B(net32),
    .C(net39),
    .D(net40),
    .Y(_03623_));
 sky130_fd_sc_hd__a22oi_2 _14164_ (.A1(net32),
    .A2(net39),
    .B1(net40),
    .B2(net31),
    .Y(_03624_));
 sky130_fd_sc_hd__nand2_1 _14165_ (.A(_03321_),
    .B(_03621_),
    .Y(_03625_));
 sky130_fd_sc_hd__a2bb2oi_1 _14166_ (.A1_N(_01868_),
    .A2_N(_02010_),
    .B1(_03623_),
    .B2(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__o22ai_1 _14167_ (.A1(_01868_),
    .A2(_02010_),
    .B1(_03622_),
    .B2(_03624_),
    .Y(_03627_));
 sky130_fd_sc_hd__o2111a_2 _14168_ (.A1(_03323_),
    .A2(_03620_),
    .B1(net30),
    .C1(net41),
    .D1(_03625_),
    .X(_03629_));
 sky130_fd_sc_hd__o2111ai_1 _14169_ (.A1(_03323_),
    .A2(_03620_),
    .B1(net30),
    .C1(net41),
    .D1(_03625_),
    .Y(_03630_));
 sky130_fd_sc_hd__o22ai_4 _14170_ (.A1(_03395_),
    .A2(_03618_),
    .B1(_03626_),
    .B2(_03629_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_1 _14171_ (.A(_03627_),
    .B(_03619_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand3_1 _14172_ (.A(_03627_),
    .B(_03630_),
    .C(_03619_),
    .Y(_03633_));
 sky130_fd_sc_hd__o22a_1 _14173_ (.A1(_01857_),
    .A2(_02010_),
    .B1(_03088_),
    .B2(_03321_),
    .X(_03634_));
 sky130_fd_sc_hd__a31o_2 _14174_ (.A1(_03327_),
    .A2(net41),
    .A3(net29),
    .B1(_03324_),
    .X(_03635_));
 sky130_fd_sc_hd__a21oi_1 _14175_ (.A1(_03631_),
    .A2(_03633_),
    .B1(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__o2bb2ai_2 _14176_ (.A1_N(_03631_),
    .A2_N(_03633_),
    .B1(_03634_),
    .B2(_03326_),
    .Y(_03637_));
 sky130_fd_sc_hd__and3_2 _14177_ (.A(_03631_),
    .B(_03633_),
    .C(_03635_),
    .X(_03638_));
 sky130_fd_sc_hd__o211ai_2 _14178_ (.A1(_03629_),
    .A2(_03632_),
    .B1(_03635_),
    .C1(_03631_),
    .Y(_03640_));
 sky130_fd_sc_hd__a21oi_1 _14179_ (.A1(_03637_),
    .A2(_03640_),
    .B1(_03616_),
    .Y(_03641_));
 sky130_fd_sc_hd__o21bai_4 _14180_ (.A1(_03636_),
    .A2(_03638_),
    .B1_N(_03616_),
    .Y(_03642_));
 sky130_fd_sc_hd__o21ai_2 _14181_ (.A1(_03336_),
    .A2(_03343_),
    .B1(_03637_),
    .Y(_03643_));
 sky130_fd_sc_hd__o211a_1 _14182_ (.A1(_03336_),
    .A2(_03343_),
    .B1(_03637_),
    .C1(_03640_),
    .X(_03644_));
 sky130_fd_sc_hd__o211ai_1 _14183_ (.A1(_03336_),
    .A2(_03343_),
    .B1(_03637_),
    .C1(_03640_),
    .Y(_03645_));
 sky130_fd_sc_hd__o21ai_1 _14184_ (.A1(_01791_),
    .A2(_02054_),
    .B1(_03356_),
    .Y(_03646_));
 sky130_fd_sc_hd__o21ai_1 _14185_ (.A1(_03352_),
    .A2(_03353_),
    .B1(_03356_),
    .Y(_03647_));
 sky130_fd_sc_hd__nand2_1 _14186_ (.A(net27),
    .B(net45),
    .Y(_03648_));
 sky130_fd_sc_hd__a22oi_4 _14187_ (.A1(net29),
    .A2(net42),
    .B1(net43),
    .B2(net28),
    .Y(_03649_));
 sky130_fd_sc_hd__a22o_1 _14188_ (.A1(net29),
    .A2(net42),
    .B1(net43),
    .B2(net28),
    .X(_03651_));
 sky130_fd_sc_hd__and4_1 _14189_ (.A(net28),
    .B(net29),
    .C(net42),
    .D(net43),
    .X(_03652_));
 sky130_fd_sc_hd__nand4_4 _14190_ (.A(net28),
    .B(net29),
    .C(net42),
    .D(net43),
    .Y(_03653_));
 sky130_fd_sc_hd__a22oi_1 _14191_ (.A1(net27),
    .A2(net45),
    .B1(_03651_),
    .B2(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__o22ai_4 _14192_ (.A1(_01769_),
    .A2(_02054_),
    .B1(_03649_),
    .B2(_03652_),
    .Y(_03655_));
 sky130_fd_sc_hd__nor3_1 _14193_ (.A(_03648_),
    .B(_03649_),
    .C(_03652_),
    .Y(_03656_));
 sky130_fd_sc_hd__nand4_2 _14194_ (.A(_03651_),
    .B(_03653_),
    .C(net27),
    .D(net45),
    .Y(_03657_));
 sky130_fd_sc_hd__a22oi_4 _14195_ (.A1(_03354_),
    .A2(_03646_),
    .B1(_03655_),
    .B2(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__o21bai_2 _14196_ (.A1(_03654_),
    .A2(_03656_),
    .B1_N(_03647_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_1 _14197_ (.A(_03655_),
    .B(_03647_),
    .Y(_03660_));
 sky130_fd_sc_hd__nand3_2 _14198_ (.A(_03655_),
    .B(_03657_),
    .C(_03647_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand2_1 _14199_ (.A(net12),
    .B(net48),
    .Y(_03663_));
 sky130_fd_sc_hd__a22oi_2 _14200_ (.A1(net26),
    .A2(net46),
    .B1(net47),
    .B2(net23),
    .Y(_03664_));
 sky130_fd_sc_hd__and4_1 _14201_ (.A(net26),
    .B(net23),
    .C(net46),
    .D(net47),
    .X(_03665_));
 sky130_fd_sc_hd__nand4_2 _14202_ (.A(net26),
    .B(net23),
    .C(net46),
    .D(net47),
    .Y(_03666_));
 sky130_fd_sc_hd__o21ai_1 _14203_ (.A1(_03664_),
    .A2(_03665_),
    .B1(_03663_),
    .Y(_03667_));
 sky130_fd_sc_hd__nand4b_2 _14204_ (.A_N(_03664_),
    .B(_03666_),
    .C(net12),
    .D(net48),
    .Y(_03668_));
 sky130_fd_sc_hd__nand2_1 _14205_ (.A(_03667_),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__a22oi_2 _14206_ (.A1(_03659_),
    .A2(_03662_),
    .B1(_03667_),
    .B2(_03668_),
    .Y(_03670_));
 sky130_fd_sc_hd__and3_1 _14207_ (.A(_03662_),
    .B(_03667_),
    .C(_03668_),
    .X(_03671_));
 sky130_fd_sc_hd__a21oi_4 _14208_ (.A1(_03659_),
    .A2(_03671_),
    .B1(_03670_),
    .Y(_03673_));
 sky130_fd_sc_hd__a21oi_1 _14209_ (.A1(_03642_),
    .A2(_03645_),
    .B1(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__o21bai_4 _14210_ (.A1(_03641_),
    .A2(_03644_),
    .B1_N(_03673_),
    .Y(_03675_));
 sky130_fd_sc_hd__o211a_1 _14211_ (.A1(_03638_),
    .A2(_03643_),
    .B1(_03673_),
    .C1(_03642_),
    .X(_03676_));
 sky130_fd_sc_hd__o211ai_4 _14212_ (.A1(_03638_),
    .A2(_03643_),
    .B1(_03673_),
    .C1(_03642_),
    .Y(_03677_));
 sky130_fd_sc_hd__a22oi_4 _14213_ (.A1(_03429_),
    .A2(_03430_),
    .B1(_03675_),
    .B2(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__o2bb2ai_2 _14214_ (.A1_N(_03429_),
    .A2_N(_03430_),
    .B1(_03674_),
    .B2(_03676_),
    .Y(_03679_));
 sky130_fd_sc_hd__o21ai_1 _14215_ (.A1(_03427_),
    .A2(_03431_),
    .B1(_03675_),
    .Y(_03680_));
 sky130_fd_sc_hd__o211a_1 _14216_ (.A1(_03427_),
    .A2(_03431_),
    .B1(_03675_),
    .C1(_03677_),
    .X(_03681_));
 sky130_fd_sc_hd__o211ai_4 _14217_ (.A1(_03427_),
    .A2(_03431_),
    .B1(_03675_),
    .C1(_03677_),
    .Y(_03682_));
 sky130_fd_sc_hd__o31a_2 _14218_ (.A1(_03316_),
    .A2(_03341_),
    .A3(_03346_),
    .B1(_03375_),
    .X(_03684_));
 sky130_fd_sc_hd__a2bb2o_1 _14219_ (.A1_N(_03346_),
    .A2_N(_03348_),
    .B1(_03347_),
    .B2(_03371_),
    .X(_03685_));
 sky130_fd_sc_hd__a21oi_4 _14220_ (.A1(_03679_),
    .A2(_03682_),
    .B1(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__o21ai_1 _14221_ (.A1(_03678_),
    .A2(_03681_),
    .B1(_03684_),
    .Y(_03687_));
 sky130_fd_sc_hd__a21oi_1 _14222_ (.A1(_03349_),
    .A2(_03375_),
    .B1(_03678_),
    .Y(_03688_));
 sky130_fd_sc_hd__nand2_1 _14223_ (.A(_03679_),
    .B(_03685_),
    .Y(_03689_));
 sky130_fd_sc_hd__and3_2 _14224_ (.A(_03679_),
    .B(_03682_),
    .C(_03685_),
    .X(_03690_));
 sky130_fd_sc_hd__a21oi_2 _14225_ (.A1(_03682_),
    .A2(_03688_),
    .B1(_03686_),
    .Y(_03691_));
 sky130_fd_sc_hd__o21ai_1 _14226_ (.A1(_03681_),
    .A2(_03689_),
    .B1(_03687_),
    .Y(_03692_));
 sky130_fd_sc_hd__o21a_1 _14227_ (.A1(_01835_),
    .A2(_02021_),
    .B1(_03463_),
    .X(_03693_));
 sky130_fd_sc_hd__o21ai_1 _14228_ (.A1(_03458_),
    .A2(_03460_),
    .B1(_03463_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_1 _14229_ (.A(net62),
    .B(net10),
    .Y(_03696_));
 sky130_fd_sc_hd__nand2_2 _14230_ (.A(net61),
    .B(net10),
    .Y(_03697_));
 sky130_fd_sc_hd__and4_1 _14231_ (.A(net61),
    .B(net62),
    .C(net9),
    .D(net10),
    .X(_03698_));
 sky130_fd_sc_hd__nand4_1 _14232_ (.A(net61),
    .B(net62),
    .C(net9),
    .D(net10),
    .Y(_03699_));
 sky130_fd_sc_hd__a22o_1 _14233_ (.A1(net62),
    .A2(net9),
    .B1(net10),
    .B2(net61),
    .X(_03700_));
 sky130_fd_sc_hd__a2bb2oi_1 _14234_ (.A1_N(_01890_),
    .A2_N(_01988_),
    .B1(_03699_),
    .B2(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__o2bb2ai_1 _14235_ (.A1_N(_03699_),
    .A2_N(_03700_),
    .B1(_01890_),
    .B2(_01988_),
    .Y(_03702_));
 sky130_fd_sc_hd__o2111a_1 _14236_ (.A1(_03493_),
    .A2(_03696_),
    .B1(net63),
    .C1(net8),
    .D1(_03700_),
    .X(_03703_));
 sky130_fd_sc_hd__o2111ai_1 _14237_ (.A1(_03493_),
    .A2(_03696_),
    .B1(net63),
    .C1(net8),
    .D1(_03700_),
    .Y(_03704_));
 sky130_fd_sc_hd__o22ai_4 _14238_ (.A1(_03460_),
    .A2(_03693_),
    .B1(_03701_),
    .B2(_03703_),
    .Y(_03706_));
 sky130_fd_sc_hd__nand2_1 _14239_ (.A(_03702_),
    .B(_03695_),
    .Y(_03707_));
 sky130_fd_sc_hd__nand3_2 _14240_ (.A(_03702_),
    .B(_03704_),
    .C(_03695_),
    .Y(_03708_));
 sky130_fd_sc_hd__a31o_1 _14241_ (.A1(_03494_),
    .A2(net7),
    .A3(net63),
    .B1(_03492_),
    .X(_03709_));
 sky130_fd_sc_hd__a21oi_2 _14242_ (.A1(_03706_),
    .A2(_03708_),
    .B1(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__a21o_1 _14243_ (.A1(_03706_),
    .A2(_03708_),
    .B1(_03709_),
    .X(_03711_));
 sky130_fd_sc_hd__and3_1 _14244_ (.A(_03706_),
    .B(_03708_),
    .C(_03709_),
    .X(_03712_));
 sky130_fd_sc_hd__nand3_1 _14245_ (.A(_03706_),
    .B(_03708_),
    .C(_03709_),
    .Y(_03713_));
 sky130_fd_sc_hd__nand2_1 _14246_ (.A(_03711_),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__o21ai_1 _14247_ (.A1(_01780_),
    .A2(_02065_),
    .B1(_03448_),
    .Y(_03715_));
 sky130_fd_sc_hd__o21ai_2 _14248_ (.A1(_03444_),
    .A2(_03445_),
    .B1(_03448_),
    .Y(_03717_));
 sky130_fd_sc_hd__o21a_1 _14249_ (.A1(_03444_),
    .A2(_03445_),
    .B1(_03448_),
    .X(_03718_));
 sky130_fd_sc_hd__nand2_1 _14250_ (.A(net55),
    .B(net15),
    .Y(_03719_));
 sky130_fd_sc_hd__a22oi_4 _14251_ (.A1(net44),
    .A2(net16),
    .B1(net17),
    .B2(net33),
    .Y(_03720_));
 sky130_fd_sc_hd__a22o_2 _14252_ (.A1(net44),
    .A2(net16),
    .B1(net17),
    .B2(net33),
    .X(_03721_));
 sky130_fd_sc_hd__and4_1 _14253_ (.A(net33),
    .B(net44),
    .C(net16),
    .D(net17),
    .X(_03722_));
 sky130_fd_sc_hd__nand4_2 _14254_ (.A(net33),
    .B(net44),
    .C(net16),
    .D(net17),
    .Y(_03723_));
 sky130_fd_sc_hd__o211ai_2 _14255_ (.A1(_01780_),
    .A2(_02076_),
    .B1(_03721_),
    .C1(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__o21bai_1 _14256_ (.A1(_03720_),
    .A2(_03722_),
    .B1_N(_03719_),
    .Y(_03725_));
 sky130_fd_sc_hd__o22a_2 _14257_ (.A1(_01780_),
    .A2(_02076_),
    .B1(_03720_),
    .B2(_03722_),
    .X(_03726_));
 sky130_fd_sc_hd__o22ai_4 _14258_ (.A1(_01780_),
    .A2(_02076_),
    .B1(_03720_),
    .B2(_03722_),
    .Y(_03728_));
 sky130_fd_sc_hd__a41o_1 _14259_ (.A1(net33),
    .A2(net44),
    .A3(net16),
    .A4(net17),
    .B1(_03719_),
    .X(_03729_));
 sky130_fd_sc_hd__nand4_1 _14260_ (.A(_03721_),
    .B(_03723_),
    .C(net55),
    .D(net15),
    .Y(_03730_));
 sky130_fd_sc_hd__a22oi_2 _14261_ (.A1(_03446_),
    .A2(_03715_),
    .B1(_03728_),
    .B2(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand3_4 _14262_ (.A(_03718_),
    .B(_03724_),
    .C(_03725_),
    .Y(_03732_));
 sky130_fd_sc_hd__o21ai_4 _14263_ (.A1(_03720_),
    .A2(_03729_),
    .B1(_03717_),
    .Y(_03733_));
 sky130_fd_sc_hd__o211ai_4 _14264_ (.A1(_03720_),
    .A2(_03729_),
    .B1(_03717_),
    .C1(_03728_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _14265_ (.A(net60),
    .B(net11),
    .Y(_03735_));
 sky130_fd_sc_hd__nand2_2 _14266_ (.A(net59),
    .B(net14),
    .Y(_03736_));
 sky130_fd_sc_hd__and4_1 _14267_ (.A(net58),
    .B(net59),
    .C(net13),
    .D(net14),
    .X(_03737_));
 sky130_fd_sc_hd__a22oi_4 _14268_ (.A1(net59),
    .A2(net13),
    .B1(net14),
    .B2(net58),
    .Y(_03739_));
 sky130_fd_sc_hd__a22o_1 _14269_ (.A1(net59),
    .A2(net13),
    .B1(net14),
    .B2(net58),
    .X(_03740_));
 sky130_fd_sc_hd__o221ai_1 _14270_ (.A1(_01835_),
    .A2(_02032_),
    .B1(_03459_),
    .B2(_03736_),
    .C1(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__o21bai_1 _14271_ (.A1(_03737_),
    .A2(_03739_),
    .B1_N(_03735_),
    .Y(_03742_));
 sky130_fd_sc_hd__o22a_1 _14272_ (.A1(_01835_),
    .A2(_02032_),
    .B1(_03737_),
    .B2(_03739_),
    .X(_03743_));
 sky130_fd_sc_hd__o22ai_2 _14273_ (.A1(_01835_),
    .A2(_02032_),
    .B1(_03737_),
    .B2(_03739_),
    .Y(_03744_));
 sky130_fd_sc_hd__o2111a_1 _14274_ (.A1(_03459_),
    .A2(_03736_),
    .B1(net60),
    .C1(net11),
    .D1(_03740_),
    .X(_03745_));
 sky130_fd_sc_hd__o2111ai_4 _14275_ (.A1(_03459_),
    .A2(_03736_),
    .B1(net60),
    .C1(net11),
    .D1(_03740_),
    .Y(_03746_));
 sky130_fd_sc_hd__nand2_1 _14276_ (.A(_03744_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand2_1 _14277_ (.A(_03741_),
    .B(_03742_),
    .Y(_03748_));
 sky130_fd_sc_hd__a21o_1 _14278_ (.A1(_03732_),
    .A2(_03734_),
    .B1(_03747_),
    .X(_03750_));
 sky130_fd_sc_hd__o221ai_2 _14279_ (.A1(_03726_),
    .A2(_03733_),
    .B1(_03743_),
    .B2(_03745_),
    .C1(_03732_),
    .Y(_03751_));
 sky130_fd_sc_hd__o2bb2ai_2 _14280_ (.A1_N(_03732_),
    .A2_N(_03734_),
    .B1(_03743_),
    .B2(_03745_),
    .Y(_03752_));
 sky130_fd_sc_hd__nand4_4 _14281_ (.A(_03732_),
    .B(_03734_),
    .C(_03744_),
    .D(_03746_),
    .Y(_03753_));
 sky130_fd_sc_hd__a32oi_2 _14282_ (.A1(_03441_),
    .A2(_03451_),
    .A3(_03452_),
    .B1(_03455_),
    .B2(_03474_),
    .Y(_03754_));
 sky130_fd_sc_hd__o2bb2ai_2 _14283_ (.A1_N(_03451_),
    .A2_N(_03456_),
    .B1(_03473_),
    .B2(_03453_),
    .Y(_03755_));
 sky130_fd_sc_hd__a21oi_4 _14284_ (.A1(_03752_),
    .A2(_03753_),
    .B1(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand3_2 _14285_ (.A(_03750_),
    .B(_03751_),
    .C(_03754_),
    .Y(_03757_));
 sky130_fd_sc_hd__nand3_4 _14286_ (.A(_03752_),
    .B(_03753_),
    .C(_03755_),
    .Y(_03758_));
 sky130_fd_sc_hd__a21o_2 _14287_ (.A1(_03757_),
    .A2(_03758_),
    .B1(_03714_),
    .X(_03759_));
 sky130_fd_sc_hd__o211ai_4 _14288_ (.A1(_03710_),
    .A2(_03712_),
    .B1(_03757_),
    .C1(_03758_),
    .Y(_03761_));
 sky130_fd_sc_hd__a22o_1 _14289_ (.A1(_03711_),
    .A2(_03713_),
    .B1(_03757_),
    .B2(_03758_),
    .X(_03762_));
 sky130_fd_sc_hd__nand3_1 _14290_ (.A(_03711_),
    .B(_03713_),
    .C(_03758_),
    .Y(_03763_));
 sky130_fd_sc_hd__a21oi_4 _14291_ (.A1(_03507_),
    .A2(_03482_),
    .B1(_03483_),
    .Y(_03764_));
 sky130_fd_sc_hd__a22oi_4 _14292_ (.A1(_03484_),
    .A2(_03513_),
    .B1(_03759_),
    .B2(_03761_),
    .Y(_03765_));
 sky130_fd_sc_hd__o221ai_4 _14293_ (.A1(_03756_),
    .A2(_03763_),
    .B1(_03483_),
    .B2(_03512_),
    .C1(_03762_),
    .Y(_03766_));
 sky130_fd_sc_hd__and3_1 _14294_ (.A(_03759_),
    .B(_03764_),
    .C(_03761_),
    .X(_03767_));
 sky130_fd_sc_hd__nand3_4 _14295_ (.A(_03759_),
    .B(_03761_),
    .C(_03764_),
    .Y(_03768_));
 sky130_fd_sc_hd__nor2_1 _14296_ (.A(_03501_),
    .B(_03504_),
    .Y(_03769_));
 sky130_fd_sc_hd__a31o_1 _14297_ (.A1(_03187_),
    .A2(_03486_),
    .A3(_03503_),
    .B1(_03501_),
    .X(_03770_));
 sky130_fd_sc_hd__nand2_1 _14298_ (.A(net2),
    .B(net38),
    .Y(_03772_));
 sky130_fd_sc_hd__a22oi_4 _14299_ (.A1(net4),
    .A2(net36),
    .B1(net37),
    .B2(net3),
    .Y(_03773_));
 sky130_fd_sc_hd__a22o_1 _14300_ (.A1(net4),
    .A2(net36),
    .B1(net37),
    .B2(net3),
    .X(_03774_));
 sky130_fd_sc_hd__nand4_4 _14301_ (.A(net3),
    .B(net4),
    .C(net36),
    .D(net37),
    .Y(_03775_));
 sky130_fd_sc_hd__a22oi_4 _14302_ (.A1(net2),
    .A2(net38),
    .B1(_03774_),
    .B2(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__and4_1 _14303_ (.A(_03774_),
    .B(_03775_),
    .C(net2),
    .D(net38),
    .X(_03777_));
 sky130_fd_sc_hd__nor2_1 _14304_ (.A(_03776_),
    .B(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__nor2_1 _14305_ (.A(_03407_),
    .B(_03411_),
    .Y(_03779_));
 sky130_fd_sc_hd__a31o_1 _14306_ (.A1(_03412_),
    .A2(net4),
    .A3(net35),
    .B1(_03408_),
    .X(_03780_));
 sky130_fd_sc_hd__o31a_1 _14307_ (.A1(_01934_),
    .A2(_01945_),
    .A3(_03411_),
    .B1(_03409_),
    .X(_03781_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(net35),
    .B(net5),
    .Y(_03783_));
 sky130_fd_sc_hd__nand4_4 _14309_ (.A(net64),
    .B(net34),
    .C(net6),
    .D(net7),
    .Y(_03784_));
 sky130_fd_sc_hd__a22oi_1 _14310_ (.A1(net34),
    .A2(net6),
    .B1(net7),
    .B2(net64),
    .Y(_03785_));
 sky130_fd_sc_hd__a22o_1 _14311_ (.A1(net34),
    .A2(net6),
    .B1(net7),
    .B2(net64),
    .X(_03786_));
 sky130_fd_sc_hd__o211ai_1 _14312_ (.A1(_01934_),
    .A2(_01956_),
    .B1(_03784_),
    .C1(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__a21o_1 _14313_ (.A1(_03784_),
    .A2(_03786_),
    .B1(_03783_),
    .X(_03788_));
 sky130_fd_sc_hd__nand4_2 _14314_ (.A(_03786_),
    .B(net5),
    .C(net35),
    .D(_03784_),
    .Y(_03789_));
 sky130_fd_sc_hd__o2bb2ai_2 _14315_ (.A1_N(_03784_),
    .A2_N(_03786_),
    .B1(_01934_),
    .B2(_01956_),
    .Y(_03790_));
 sky130_fd_sc_hd__o211a_2 _14316_ (.A1(_03408_),
    .A2(_03779_),
    .B1(_03789_),
    .C1(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__o211ai_1 _14317_ (.A1(_03408_),
    .A2(_03779_),
    .B1(_03789_),
    .C1(_03790_),
    .Y(_03792_));
 sky130_fd_sc_hd__a21oi_2 _14318_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03780_),
    .Y(_03794_));
 sky130_fd_sc_hd__nand3_1 _14319_ (.A(_03781_),
    .B(_03787_),
    .C(_03788_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _14320_ (.A(_03778_),
    .B(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__nand3_1 _14321_ (.A(_03778_),
    .B(_03792_),
    .C(_03795_),
    .Y(_03797_));
 sky130_fd_sc_hd__o22ai_4 _14322_ (.A1(_03776_),
    .A2(_03777_),
    .B1(_03791_),
    .B2(_03794_),
    .Y(_03798_));
 sky130_fd_sc_hd__o21a_1 _14323_ (.A1(_03791_),
    .A2(_03796_),
    .B1(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__o21ai_2 _14324_ (.A1(_03791_),
    .A2(_03796_),
    .B1(_03798_),
    .Y(_03800_));
 sky130_fd_sc_hd__a21oi_1 _14325_ (.A1(_03797_),
    .A2(_03798_),
    .B1(_03770_),
    .Y(_03801_));
 sky130_fd_sc_hd__a21o_1 _14326_ (.A1(_03797_),
    .A2(_03798_),
    .B1(_03770_),
    .X(_03802_));
 sky130_fd_sc_hd__o221a_2 _14327_ (.A1(_03501_),
    .A2(_03504_),
    .B1(_03791_),
    .B2(_03796_),
    .C1(_03798_),
    .X(_03803_));
 sky130_fd_sc_hd__o211ai_2 _14328_ (.A1(_03501_),
    .A2(_03504_),
    .B1(_03797_),
    .C1(_03798_),
    .Y(_03805_));
 sky130_fd_sc_hd__o31a_1 _14329_ (.A1(_03400_),
    .A2(_03401_),
    .A3(_03419_),
    .B1(_03418_),
    .X(_03806_));
 sky130_fd_sc_hd__nand2_1 _14330_ (.A(_03418_),
    .B(_03424_),
    .Y(_03807_));
 sky130_fd_sc_hd__a21oi_1 _14331_ (.A1(_03802_),
    .A2(_03805_),
    .B1(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__o21ai_2 _14332_ (.A1(_03801_),
    .A2(_03803_),
    .B1(_03806_),
    .Y(_03809_));
 sky130_fd_sc_hd__a22oi_4 _14333_ (.A1(_03418_),
    .A2(_03424_),
    .B1(_03800_),
    .B2(_03769_),
    .Y(_03810_));
 sky130_fd_sc_hd__and3_1 _14334_ (.A(_03802_),
    .B(_03805_),
    .C(_03807_),
    .X(_03811_));
 sky130_fd_sc_hd__o21ai_2 _14335_ (.A1(_03769_),
    .A2(_03800_),
    .B1(_03810_),
    .Y(_03812_));
 sky130_fd_sc_hd__nand3_1 _14336_ (.A(_03802_),
    .B(_03805_),
    .C(_03806_),
    .Y(_03813_));
 sky130_fd_sc_hd__o2bb2ai_1 _14337_ (.A1_N(_03418_),
    .A2_N(_03424_),
    .B1(_03801_),
    .B2(_03803_),
    .Y(_03814_));
 sky130_fd_sc_hd__o2bb2ai_4 _14338_ (.A1_N(_03766_),
    .A2_N(_03768_),
    .B1(_03808_),
    .B2(_03811_),
    .Y(_03816_));
 sky130_fd_sc_hd__a32oi_4 _14339_ (.A1(_03759_),
    .A2(_03764_),
    .A3(_03761_),
    .B1(_03814_),
    .B2(_03813_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand3_1 _14340_ (.A(_03768_),
    .B(_03809_),
    .C(_03812_),
    .Y(_03818_));
 sky130_fd_sc_hd__and4_2 _14341_ (.A(_03766_),
    .B(_03768_),
    .C(_03809_),
    .D(_03812_),
    .X(_03819_));
 sky130_fd_sc_hd__nand4_2 _14342_ (.A(_03766_),
    .B(_03768_),
    .C(_03809_),
    .D(_03812_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21oi_4 _14343_ (.A1(_03816_),
    .A2(_03820_),
    .B1(_03523_),
    .Y(_03821_));
 sky130_fd_sc_hd__a21o_2 _14344_ (.A1(_03816_),
    .A2(_03820_),
    .B1(_03523_),
    .X(_03822_));
 sky130_fd_sc_hd__nand2_2 _14345_ (.A(_03523_),
    .B(_03816_),
    .Y(_03823_));
 sky130_fd_sc_hd__o211a_1 _14346_ (.A1(_03765_),
    .A2(_03818_),
    .B1(_03816_),
    .C1(_03523_),
    .X(_03824_));
 sky130_fd_sc_hd__o211ai_2 _14347_ (.A1(_03765_),
    .A2(_03818_),
    .B1(_03816_),
    .C1(_03523_),
    .Y(_03825_));
 sky130_fd_sc_hd__o221ai_4 _14348_ (.A1(_03686_),
    .A2(_03690_),
    .B1(_03819_),
    .B2(_03823_),
    .C1(_03822_),
    .Y(_03827_));
 sky130_fd_sc_hd__o21ai_4 _14349_ (.A1(_03821_),
    .A2(_03824_),
    .B1(_03691_),
    .Y(_03828_));
 sky130_fd_sc_hd__o22ai_2 _14350_ (.A1(_03686_),
    .A2(_03690_),
    .B1(_03821_),
    .B2(_03824_),
    .Y(_03829_));
 sky130_fd_sc_hd__nand3_1 _14351_ (.A(_03691_),
    .B(_03822_),
    .C(_03825_),
    .Y(_03830_));
 sky130_fd_sc_hd__a22oi_1 _14352_ (.A1(_03534_),
    .A2(_03614_),
    .B1(_03829_),
    .B2(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__o211ai_4 _14353_ (.A1(_03533_),
    .A2(_03613_),
    .B1(_03827_),
    .C1(_03828_),
    .Y(_03832_));
 sky130_fd_sc_hd__a2bb2oi_4 _14354_ (.A1_N(_03535_),
    .A2_N(_03539_),
    .B1(_03827_),
    .B2(_03828_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand3_2 _14355_ (.A(_03615_),
    .B(_03829_),
    .C(_03830_),
    .Y(_03834_));
 sky130_fd_sc_hd__o22ai_1 _14356_ (.A1(_03608_),
    .A2(_03609_),
    .B1(_03831_),
    .B2(_03833_),
    .Y(_03835_));
 sky130_fd_sc_hd__a41oi_4 _14357_ (.A1(_03536_),
    .A2(_03540_),
    .A3(_03827_),
    .A4(_03828_),
    .B1(_03612_),
    .Y(_03836_));
 sky130_fd_sc_hd__nand4_1 _14358_ (.A(_03607_),
    .B(_03610_),
    .C(_03832_),
    .D(_03834_),
    .Y(_03838_));
 sky130_fd_sc_hd__a21o_1 _14359_ (.A1(_03832_),
    .A2(_03834_),
    .B1(_03612_),
    .X(_03839_));
 sky130_fd_sc_hd__o211ai_4 _14360_ (.A1(_03608_),
    .A2(_03609_),
    .B1(_03832_),
    .C1(_03834_),
    .Y(_03840_));
 sky130_fd_sc_hd__a32oi_4 _14361_ (.A1(_03538_),
    .A2(_03541_),
    .A3(_03545_),
    .B1(_03548_),
    .B2(_03559_),
    .Y(_03841_));
 sky130_fd_sc_hd__a21oi_1 _14362_ (.A1(_03546_),
    .A2(_03560_),
    .B1(_03547_),
    .Y(_03842_));
 sky130_fd_sc_hd__a21oi_2 _14363_ (.A1(_03839_),
    .A2(_03840_),
    .B1(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand3_1 _14364_ (.A(_03835_),
    .B(_03838_),
    .C(_03842_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand3_2 _14365_ (.A(_03839_),
    .B(_03840_),
    .C(_03841_),
    .Y(_03845_));
 sky130_fd_sc_hd__o2bb2ai_2 _14366_ (.A1_N(_03844_),
    .A2_N(_03845_),
    .B1(_03550_),
    .B2(_03552_),
    .Y(_03846_));
 sky130_fd_sc_hd__a31oi_2 _14367_ (.A1(_03839_),
    .A2(_03841_),
    .A3(_03840_),
    .B1(_03555_),
    .Y(_03847_));
 sky130_fd_sc_hd__a31o_1 _14368_ (.A1(_03839_),
    .A2(_03840_),
    .A3(_03841_),
    .B1(_03555_),
    .X(_03849_));
 sky130_fd_sc_hd__nand3_1 _14369_ (.A(_03845_),
    .B(_03554_),
    .C(_03844_),
    .Y(_03850_));
 sky130_fd_sc_hd__o21ai_1 _14370_ (.A1(_03843_),
    .A2(_03849_),
    .B1(_03846_),
    .Y(_03851_));
 sky130_fd_sc_hd__o32a_1 _14371_ (.A1(_03561_),
    .A2(_03563_),
    .A3(_03570_),
    .B1(_03285_),
    .B2(_03571_),
    .X(_03852_));
 sky130_fd_sc_hd__o32ai_4 _14372_ (.A1(_03561_),
    .A2(_03570_),
    .A3(_03563_),
    .B1(_03285_),
    .B2(_03571_),
    .Y(_03853_));
 sky130_fd_sc_hd__a21oi_1 _14373_ (.A1(_03846_),
    .A2(_03850_),
    .B1(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__a21o_1 _14374_ (.A1(_03846_),
    .A2(_03850_),
    .B1(_03853_),
    .X(_03855_));
 sky130_fd_sc_hd__o211a_1 _14375_ (.A1(_03843_),
    .A2(_03849_),
    .B1(_03853_),
    .C1(_03846_),
    .X(_03856_));
 sky130_fd_sc_hd__o211ai_1 _14376_ (.A1(_03843_),
    .A2(_03849_),
    .B1(_03853_),
    .C1(_03846_),
    .Y(_03857_));
 sky130_fd_sc_hd__o22ai_2 _14377_ (.A1(_03580_),
    .A2(_03581_),
    .B1(_03854_),
    .B2(_03856_),
    .Y(_03858_));
 sky130_fd_sc_hd__a21oi_1 _14378_ (.A1(_03851_),
    .A2(_03852_),
    .B1(_03584_),
    .Y(_03860_));
 sky130_fd_sc_hd__nand3_1 _14379_ (.A(_03855_),
    .B(_03857_),
    .C(_03583_),
    .Y(_03861_));
 sky130_fd_sc_hd__nand2_1 _14380_ (.A(_03858_),
    .B(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand4_2 _14381_ (.A(_03309_),
    .B(_03311_),
    .C(_03587_),
    .D(_03588_),
    .Y(_03863_));
 sky130_fd_sc_hd__nor3_4 _14382_ (.A(_02794_),
    .B(_03053_),
    .C(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__nand4_2 _14383_ (.A(_02793_),
    .B(_03052_),
    .C(_03313_),
    .D(_03589_),
    .Y(_03865_));
 sky130_fd_sc_hd__nand4_4 _14384_ (.A(_02792_),
    .B(_03052_),
    .C(_03313_),
    .D(_03589_),
    .Y(_03866_));
 sky130_fd_sc_hd__o2bb2a_2 _14385_ (.A1_N(_03306_),
    .A2_N(_03582_),
    .B1(_03585_),
    .B2(_03311_),
    .X(_03867_));
 sky130_fd_sc_hd__nand4_4 _14386_ (.A(_03054_),
    .B(_03589_),
    .C(_03311_),
    .D(_03309_),
    .Y(_03868_));
 sky130_fd_sc_hd__nand3_4 _14387_ (.A(_03866_),
    .B(_03867_),
    .C(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__o2111ai_4 _14388_ (.A1(_03865_),
    .A2(_01762_),
    .B1(_03867_),
    .C1(_03866_),
    .D1(_03868_),
    .Y(_03871_));
 sky130_fd_sc_hd__xnor2_1 _14389_ (.A(_03862_),
    .B(_03871_),
    .Y(net81));
 sky130_fd_sc_hd__a21oi_1 _14390_ (.A1(_03554_),
    .A2(_03845_),
    .B1(_03843_),
    .Y(_03872_));
 sky130_fd_sc_hd__a32o_1 _14391_ (.A1(_03835_),
    .A2(_03838_),
    .A3(_03842_),
    .B1(_03845_),
    .B2(_03554_),
    .X(_03873_));
 sky130_fd_sc_hd__o21ai_2 _14392_ (.A1(_03686_),
    .A2(_03690_),
    .B1(_03825_),
    .Y(_03874_));
 sky130_fd_sc_hd__o22ai_4 _14393_ (.A1(_03819_),
    .A2(_03823_),
    .B1(_03821_),
    .B2(_03692_),
    .Y(_03875_));
 sky130_fd_sc_hd__a21oi_1 _14394_ (.A1(_03809_),
    .A2(_03812_),
    .B1(_03765_),
    .Y(_03876_));
 sky130_fd_sc_hd__a31oi_2 _14395_ (.A1(_03768_),
    .A2(_03809_),
    .A3(_03812_),
    .B1(_03765_),
    .Y(_03877_));
 sky130_fd_sc_hd__o2bb2ai_2 _14396_ (.A1_N(_03709_),
    .A2_N(_03706_),
    .B1(_03703_),
    .B2(_03707_),
    .Y(_03878_));
 sky130_fd_sc_hd__o21ai_2 _14397_ (.A1(_03783_),
    .A2(_03785_),
    .B1(_03784_),
    .Y(_03879_));
 sky130_fd_sc_hd__nand2_1 _14398_ (.A(net35),
    .B(net6),
    .Y(_03881_));
 sky130_fd_sc_hd__a22oi_4 _14399_ (.A1(net34),
    .A2(net7),
    .B1(net8),
    .B2(net64),
    .Y(_03882_));
 sky130_fd_sc_hd__a22o_2 _14400_ (.A1(net34),
    .A2(net7),
    .B1(net8),
    .B2(net64),
    .X(_03883_));
 sky130_fd_sc_hd__and4_1 _14401_ (.A(net64),
    .B(net34),
    .C(net7),
    .D(net8),
    .X(_03884_));
 sky130_fd_sc_hd__nand4_2 _14402_ (.A(net64),
    .B(net34),
    .C(net7),
    .D(net8),
    .Y(_03885_));
 sky130_fd_sc_hd__o211ai_2 _14403_ (.A1(_01934_),
    .A2(_01966_),
    .B1(_03883_),
    .C1(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__o21bai_1 _14404_ (.A1(_03882_),
    .A2(_03884_),
    .B1_N(_03881_),
    .Y(_03887_));
 sky130_fd_sc_hd__o21ai_1 _14405_ (.A1(_03882_),
    .A2(_03884_),
    .B1(_03881_),
    .Y(_03888_));
 sky130_fd_sc_hd__a41o_1 _14406_ (.A1(net64),
    .A2(net34),
    .A3(net7),
    .A4(net8),
    .B1(_03881_),
    .X(_03889_));
 sky130_fd_sc_hd__nand3b_4 _14407_ (.A_N(_03879_),
    .B(_03886_),
    .C(_03887_),
    .Y(_03890_));
 sky130_fd_sc_hd__o211ai_4 _14408_ (.A1(_03882_),
    .A2(_03889_),
    .B1(_03879_),
    .C1(_03888_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _14409_ (.A(net3),
    .B(net38),
    .Y(_03893_));
 sky130_fd_sc_hd__a22oi_4 _14410_ (.A1(net36),
    .A2(net5),
    .B1(net37),
    .B2(net4),
    .Y(_03894_));
 sky130_fd_sc_hd__and4_1 _14411_ (.A(net4),
    .B(net36),
    .C(net5),
    .D(net37),
    .X(_03895_));
 sky130_fd_sc_hd__nand4_1 _14412_ (.A(net4),
    .B(net36),
    .C(net5),
    .D(net37),
    .Y(_03896_));
 sky130_fd_sc_hd__a211oi_2 _14413_ (.A1(net3),
    .A2(net38),
    .B1(_03894_),
    .C1(_03895_),
    .Y(_03897_));
 sky130_fd_sc_hd__a211o_1 _14414_ (.A1(net3),
    .A2(net38),
    .B1(_03894_),
    .C1(_03895_),
    .X(_03898_));
 sky130_fd_sc_hd__o211a_1 _14415_ (.A1(_03894_),
    .A2(_03895_),
    .B1(net3),
    .C1(net38),
    .X(_03899_));
 sky130_fd_sc_hd__o211ai_1 _14416_ (.A1(_03894_),
    .A2(_03895_),
    .B1(net3),
    .C1(net38),
    .Y(_03900_));
 sky130_fd_sc_hd__nand2_2 _14417_ (.A(_03898_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__a21oi_2 _14418_ (.A1(_03890_),
    .A2(_03892_),
    .B1(_03901_),
    .Y(_03903_));
 sky130_fd_sc_hd__a21o_1 _14419_ (.A1(_03890_),
    .A2(_03892_),
    .B1(_03901_),
    .X(_03904_));
 sky130_fd_sc_hd__o211a_2 _14420_ (.A1(_03897_),
    .A2(_03899_),
    .B1(_03890_),
    .C1(_03892_),
    .X(_03905_));
 sky130_fd_sc_hd__o211ai_4 _14421_ (.A1(_03897_),
    .A2(_03899_),
    .B1(_03890_),
    .C1(_03892_),
    .Y(_03906_));
 sky130_fd_sc_hd__a21oi_1 _14422_ (.A1(_03904_),
    .A2(_03906_),
    .B1(_03878_),
    .Y(_03907_));
 sky130_fd_sc_hd__o21bai_4 _14423_ (.A1(_03903_),
    .A2(_03905_),
    .B1_N(_03878_),
    .Y(_03908_));
 sky130_fd_sc_hd__a21o_1 _14424_ (.A1(_03708_),
    .A2(_03713_),
    .B1(_03903_),
    .X(_03909_));
 sky130_fd_sc_hd__nand3_2 _14425_ (.A(_03878_),
    .B(_03904_),
    .C(_03906_),
    .Y(_03910_));
 sky130_fd_sc_hd__o31a_1 _14426_ (.A1(_03776_),
    .A2(_03777_),
    .A3(_03794_),
    .B1(_03792_),
    .X(_03911_));
 sky130_fd_sc_hd__a32o_2 _14427_ (.A1(_03780_),
    .A2(_03789_),
    .A3(_03790_),
    .B1(_03795_),
    .B2(_03778_),
    .X(_03912_));
 sky130_fd_sc_hd__a21oi_4 _14428_ (.A1(_03908_),
    .A2(_03910_),
    .B1(_03912_),
    .Y(_03914_));
 sky130_fd_sc_hd__a21o_1 _14429_ (.A1(_03908_),
    .A2(_03910_),
    .B1(_03912_),
    .X(_03915_));
 sky130_fd_sc_hd__and3_2 _14430_ (.A(_03908_),
    .B(_03910_),
    .C(_03912_),
    .X(_03916_));
 sky130_fd_sc_hd__o211ai_2 _14431_ (.A1(_03905_),
    .A2(_03909_),
    .B1(_03912_),
    .C1(_03908_),
    .Y(_03917_));
 sky130_fd_sc_hd__nand2_1 _14432_ (.A(_03915_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__a31o_2 _14433_ (.A1(_03700_),
    .A2(net8),
    .A3(net63),
    .B1(_03698_),
    .X(_03919_));
 sky130_fd_sc_hd__o22ai_2 _14434_ (.A1(_03459_),
    .A2(_03736_),
    .B1(_03735_),
    .B2(_03739_),
    .Y(_03920_));
 sky130_fd_sc_hd__and2_1 _14435_ (.A(net63),
    .B(net9),
    .X(_03921_));
 sky130_fd_sc_hd__nand2_2 _14436_ (.A(net62),
    .B(net11),
    .Y(_03922_));
 sky130_fd_sc_hd__nand2_2 _14437_ (.A(net61),
    .B(net11),
    .Y(_03923_));
 sky130_fd_sc_hd__a22oi_2 _14438_ (.A1(net62),
    .A2(net10),
    .B1(net11),
    .B2(net61),
    .Y(_03925_));
 sky130_fd_sc_hd__a22o_1 _14439_ (.A1(net62),
    .A2(net10),
    .B1(net11),
    .B2(net61),
    .X(_03926_));
 sky130_fd_sc_hd__o2bb2ai_1 _14440_ (.A1_N(_03696_),
    .A2_N(_03923_),
    .B1(_03922_),
    .B2(_03697_),
    .Y(_03927_));
 sky130_fd_sc_hd__o221ai_4 _14441_ (.A1(_01890_),
    .A2(_01999_),
    .B1(_03697_),
    .B2(_03922_),
    .C1(_03926_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand2_1 _14442_ (.A(_03927_),
    .B(_03921_),
    .Y(_03929_));
 sky130_fd_sc_hd__o211a_1 _14443_ (.A1(_03697_),
    .A2(_03922_),
    .B1(_03921_),
    .C1(_03926_),
    .X(_03930_));
 sky130_fd_sc_hd__o2111ai_1 _14444_ (.A1(_03697_),
    .A2(_03922_),
    .B1(net63),
    .C1(net9),
    .D1(_03926_),
    .Y(_03931_));
 sky130_fd_sc_hd__o21ai_1 _14445_ (.A1(_01890_),
    .A2(_01999_),
    .B1(_03927_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _14446_ (.A(_03932_),
    .B(_03920_),
    .Y(_03933_));
 sky130_fd_sc_hd__and3_1 _14447_ (.A(_03932_),
    .B(_03920_),
    .C(_03931_),
    .X(_03934_));
 sky130_fd_sc_hd__nand3_1 _14448_ (.A(_03932_),
    .B(_03920_),
    .C(_03931_),
    .Y(_03936_));
 sky130_fd_sc_hd__nand3b_4 _14449_ (.A_N(_03920_),
    .B(_03928_),
    .C(_03929_),
    .Y(_03937_));
 sky130_fd_sc_hd__a21bo_1 _14450_ (.A1(_03936_),
    .A2(_03937_),
    .B1_N(_03919_),
    .X(_03938_));
 sky130_fd_sc_hd__nand3b_1 _14451_ (.A_N(_03919_),
    .B(_03936_),
    .C(_03937_),
    .Y(_03939_));
 sky130_fd_sc_hd__nand2_1 _14452_ (.A(_03937_),
    .B(_03919_),
    .Y(_03940_));
 sky130_fd_sc_hd__o211ai_1 _14453_ (.A1(_03930_),
    .A2(_03933_),
    .B1(_03937_),
    .C1(_03919_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21o_1 _14454_ (.A1(_03936_),
    .A2(_03937_),
    .B1(_03919_),
    .X(_03942_));
 sky130_fd_sc_hd__o21ai_2 _14455_ (.A1(_03934_),
    .A2(_03940_),
    .B1(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__o21ai_2 _14456_ (.A1(_01780_),
    .A2(_02076_),
    .B1(_03723_),
    .Y(_03944_));
 sky130_fd_sc_hd__o21a_1 _14457_ (.A1(_03719_),
    .A2(_03720_),
    .B1(_03723_),
    .X(_03945_));
 sky130_fd_sc_hd__nand2_1 _14458_ (.A(net55),
    .B(net16),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_2 _14459_ (.A(net33),
    .B(net18),
    .Y(_03948_));
 sky130_fd_sc_hd__a22oi_4 _14460_ (.A1(net44),
    .A2(net17),
    .B1(net18),
    .B2(net33),
    .Y(_03949_));
 sky130_fd_sc_hd__a22o_1 _14461_ (.A1(net44),
    .A2(net17),
    .B1(net18),
    .B2(net33),
    .X(_03950_));
 sky130_fd_sc_hd__and4_1 _14462_ (.A(net33),
    .B(net44),
    .C(net17),
    .D(net18),
    .X(_03951_));
 sky130_fd_sc_hd__nand4_4 _14463_ (.A(net33),
    .B(net44),
    .C(net17),
    .D(net18),
    .Y(_03952_));
 sky130_fd_sc_hd__o211ai_2 _14464_ (.A1(_01780_),
    .A2(_02098_),
    .B1(_03950_),
    .C1(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__o21bai_1 _14465_ (.A1(_03949_),
    .A2(_03951_),
    .B1_N(_03947_),
    .Y(_03954_));
 sky130_fd_sc_hd__o22a_2 _14466_ (.A1(_01780_),
    .A2(_02098_),
    .B1(_03949_),
    .B2(_03951_),
    .X(_03955_));
 sky130_fd_sc_hd__o22ai_2 _14467_ (.A1(_01780_),
    .A2(_02098_),
    .B1(_03949_),
    .B2(_03951_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand4_4 _14468_ (.A(_03950_),
    .B(_03952_),
    .C(net55),
    .D(net16),
    .Y(_03958_));
 sky130_fd_sc_hd__a22oi_1 _14469_ (.A1(_03721_),
    .A2(_03944_),
    .B1(_03956_),
    .B2(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__nand3_4 _14470_ (.A(_03945_),
    .B(_03953_),
    .C(_03954_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand3_2 _14471_ (.A(_03721_),
    .B(_03944_),
    .C(_03958_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand4_4 _14472_ (.A(_03721_),
    .B(_03944_),
    .C(_03956_),
    .D(_03958_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_2 _14473_ (.A(net60),
    .B(net13),
    .Y(_03963_));
 sky130_fd_sc_hd__a22oi_4 _14474_ (.A1(net59),
    .A2(net14),
    .B1(net15),
    .B2(net58),
    .Y(_03964_));
 sky130_fd_sc_hd__a22o_1 _14475_ (.A1(net59),
    .A2(net14),
    .B1(net15),
    .B2(net58),
    .X(_03965_));
 sky130_fd_sc_hd__and4_1 _14476_ (.A(net58),
    .B(net59),
    .C(net14),
    .D(net15),
    .X(_03966_));
 sky130_fd_sc_hd__nand4_2 _14477_ (.A(net58),
    .B(net59),
    .C(net14),
    .D(net15),
    .Y(_03967_));
 sky130_fd_sc_hd__and3_1 _14478_ (.A(_03963_),
    .B(_03965_),
    .C(_03967_),
    .X(_03969_));
 sky130_fd_sc_hd__o211ai_1 _14479_ (.A1(_01835_),
    .A2(_02043_),
    .B1(_03965_),
    .C1(_03967_),
    .Y(_03970_));
 sky130_fd_sc_hd__o211a_1 _14480_ (.A1(_03964_),
    .A2(_03966_),
    .B1(net60),
    .C1(net13),
    .X(_03971_));
 sky130_fd_sc_hd__o21bai_1 _14481_ (.A1(_03964_),
    .A2(_03966_),
    .B1_N(_03963_),
    .Y(_03972_));
 sky130_fd_sc_hd__o22a_2 _14482_ (.A1(_01835_),
    .A2(_02043_),
    .B1(_03964_),
    .B2(_03966_),
    .X(_03973_));
 sky130_fd_sc_hd__o21ai_2 _14483_ (.A1(_03964_),
    .A2(_03966_),
    .B1(_03963_),
    .Y(_03974_));
 sky130_fd_sc_hd__a41o_1 _14484_ (.A1(net58),
    .A2(net59),
    .A3(net14),
    .A4(net15),
    .B1(_03963_),
    .X(_03975_));
 sky130_fd_sc_hd__and4_2 _14485_ (.A(_03965_),
    .B(_03967_),
    .C(net60),
    .D(net13),
    .X(_03976_));
 sky130_fd_sc_hd__o21ai_1 _14486_ (.A1(_03964_),
    .A2(_03975_),
    .B1(_03974_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand2_1 _14487_ (.A(_03970_),
    .B(_03972_),
    .Y(_03978_));
 sky130_fd_sc_hd__o2bb2ai_2 _14488_ (.A1_N(_03960_),
    .A2_N(_03962_),
    .B1(_03969_),
    .B2(_03971_),
    .Y(_03980_));
 sky130_fd_sc_hd__o221ai_4 _14489_ (.A1(_03973_),
    .A2(_03976_),
    .B1(_03955_),
    .B2(_03961_),
    .C1(_03960_),
    .Y(_03981_));
 sky130_fd_sc_hd__o2bb2ai_4 _14490_ (.A1_N(_03960_),
    .A2_N(_03962_),
    .B1(_03973_),
    .B2(_03976_),
    .Y(_03982_));
 sky130_fd_sc_hd__o21ai_1 _14491_ (.A1(_03969_),
    .A2(_03971_),
    .B1(_03960_),
    .Y(_03983_));
 sky130_fd_sc_hd__o2111ai_4 _14492_ (.A1(_03964_),
    .A2(_03975_),
    .B1(_03974_),
    .C1(_03960_),
    .D1(_03962_),
    .Y(_03984_));
 sky130_fd_sc_hd__a2bb2oi_2 _14493_ (.A1_N(_03733_),
    .A2_N(_03726_),
    .B1(_03732_),
    .B2(_03748_),
    .Y(_03985_));
 sky130_fd_sc_hd__o22ai_4 _14494_ (.A1(_03726_),
    .A2(_03733_),
    .B1(_03747_),
    .B2(_03731_),
    .Y(_03986_));
 sky130_fd_sc_hd__a21oi_4 _14495_ (.A1(_03982_),
    .A2(_03984_),
    .B1(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand3_1 _14496_ (.A(_03980_),
    .B(_03985_),
    .C(_03981_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand3_4 _14497_ (.A(_03982_),
    .B(_03984_),
    .C(_03986_),
    .Y(_03989_));
 sky130_fd_sc_hd__a32o_1 _14498_ (.A1(_03982_),
    .A2(_03984_),
    .A3(_03986_),
    .B1(_03939_),
    .B2(_03938_),
    .X(_03991_));
 sky130_fd_sc_hd__o2111ai_4 _14499_ (.A1(_03934_),
    .A2(_03940_),
    .B1(_03942_),
    .C1(_03988_),
    .D1(_03989_),
    .Y(_03992_));
 sky130_fd_sc_hd__a22o_2 _14500_ (.A1(_03941_),
    .A2(_03942_),
    .B1(_03988_),
    .B2(_03989_),
    .X(_03993_));
 sky130_fd_sc_hd__o21a_1 _14501_ (.A1(_03987_),
    .A2(_03991_),
    .B1(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__o21a_1 _14502_ (.A1(_03710_),
    .A2(_03712_),
    .B1(_03758_),
    .X(_03995_));
 sky130_fd_sc_hd__o21ai_4 _14503_ (.A1(_03714_),
    .A2(_03756_),
    .B1(_03758_),
    .Y(_03996_));
 sky130_fd_sc_hd__a21oi_1 _14504_ (.A1(_03992_),
    .A2(_03993_),
    .B1(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__o2bb2ai_4 _14505_ (.A1_N(_03992_),
    .A2_N(_03993_),
    .B1(_03995_),
    .B2(_03756_),
    .Y(_03998_));
 sky130_fd_sc_hd__o211a_1 _14506_ (.A1(_03987_),
    .A2(_03991_),
    .B1(_03993_),
    .C1(_03996_),
    .X(_03999_));
 sky130_fd_sc_hd__o211ai_4 _14507_ (.A1(_03987_),
    .A2(_03991_),
    .B1(_03993_),
    .C1(_03996_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand2_1 _14508_ (.A(_03998_),
    .B(_04000_),
    .Y(_04002_));
 sky130_fd_sc_hd__nand4_4 _14509_ (.A(_03915_),
    .B(_03917_),
    .C(_03998_),
    .D(_04000_),
    .Y(_04003_));
 sky130_fd_sc_hd__o22ai_4 _14510_ (.A1(_03914_),
    .A2(_03916_),
    .B1(_03997_),
    .B2(_03999_),
    .Y(_04004_));
 sky130_fd_sc_hd__o211ai_2 _14511_ (.A1(_03914_),
    .A2(_03916_),
    .B1(_03998_),
    .C1(_04000_),
    .Y(_04005_));
 sky130_fd_sc_hd__a21o_1 _14512_ (.A1(_03998_),
    .A2(_04000_),
    .B1(_03918_),
    .X(_04006_));
 sky130_fd_sc_hd__a2bb2oi_4 _14513_ (.A1_N(_03765_),
    .A2_N(_03817_),
    .B1(_03918_),
    .B2(_04002_),
    .Y(_04007_));
 sky130_fd_sc_hd__o211a_1 _14514_ (.A1(_03765_),
    .A2(_03817_),
    .B1(_04003_),
    .C1(_04004_),
    .X(_04008_));
 sky130_fd_sc_hd__o211ai_4 _14515_ (.A1(_03765_),
    .A2(_03817_),
    .B1(_04003_),
    .C1(_04004_),
    .Y(_04009_));
 sky130_fd_sc_hd__a2bb2oi_1 _14516_ (.A1_N(_03767_),
    .A2_N(_03876_),
    .B1(_04003_),
    .B2(_04004_),
    .Y(_04010_));
 sky130_fd_sc_hd__nand3_4 _14517_ (.A(_04006_),
    .B(_03877_),
    .C(_04005_),
    .Y(_04011_));
 sky130_fd_sc_hd__a21oi_2 _14518_ (.A1(_03642_),
    .A2(_03673_),
    .B1(_03644_),
    .Y(_04013_));
 sky130_fd_sc_hd__a2bb2o_1 _14519_ (.A1_N(_03638_),
    .A2_N(_03643_),
    .B1(_03673_),
    .B2(_03642_),
    .X(_04014_));
 sky130_fd_sc_hd__nand2_1 _14520_ (.A(_03805_),
    .B(_03806_),
    .Y(_04015_));
 sky130_fd_sc_hd__o21ai_2 _14521_ (.A1(_03770_),
    .A2(_03799_),
    .B1(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__o2bb2ai_4 _14522_ (.A1_N(_03635_),
    .A2_N(_03631_),
    .B1(_03629_),
    .B2(_03632_),
    .Y(_04017_));
 sky130_fd_sc_hd__o22a_1 _14523_ (.A1(_01868_),
    .A2(_02010_),
    .B1(_03321_),
    .B2(_03621_),
    .X(_04018_));
 sky130_fd_sc_hd__and3_1 _14524_ (.A(_03625_),
    .B(net41),
    .C(net30),
    .X(_04019_));
 sky130_fd_sc_hd__and2_1 _14525_ (.A(_03772_),
    .B(_03775_),
    .X(_04020_));
 sky130_fd_sc_hd__o21ai_2 _14526_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03775_),
    .Y(_04021_));
 sky130_fd_sc_hd__o21a_1 _14527_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03775_),
    .X(_04022_));
 sky130_fd_sc_hd__and4_1 _14528_ (.A(net2),
    .B(net32),
    .C(net39),
    .D(net40),
    .X(_04024_));
 sky130_fd_sc_hd__nand4_2 _14529_ (.A(net2),
    .B(net32),
    .C(net39),
    .D(net40),
    .Y(_04025_));
 sky130_fd_sc_hd__a22oi_4 _14530_ (.A1(net2),
    .A2(net39),
    .B1(net40),
    .B2(net32),
    .Y(_04026_));
 sky130_fd_sc_hd__a22o_1 _14531_ (.A1(net2),
    .A2(net39),
    .B1(net40),
    .B2(net32),
    .X(_04027_));
 sky130_fd_sc_hd__a2bb2oi_1 _14532_ (.A1_N(_01879_),
    .A2_N(_02010_),
    .B1(_04025_),
    .B2(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__o22ai_4 _14533_ (.A1(_01879_),
    .A2(_02010_),
    .B1(_04024_),
    .B2(_04026_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand3_2 _14534_ (.A(_04025_),
    .B(net41),
    .C(net31),
    .Y(_04030_));
 sky130_fd_sc_hd__nor2_1 _14535_ (.A(_04026_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__o21ai_1 _14536_ (.A1(_04026_),
    .A2(_04030_),
    .B1(_04029_),
    .Y(_04032_));
 sky130_fd_sc_hd__o211a_1 _14537_ (.A1(_04026_),
    .A2(_04030_),
    .B1(_04021_),
    .C1(_04029_),
    .X(_04033_));
 sky130_fd_sc_hd__o211ai_4 _14538_ (.A1(_04026_),
    .A2(_04030_),
    .B1(_04021_),
    .C1(_04029_),
    .Y(_04035_));
 sky130_fd_sc_hd__o22ai_4 _14539_ (.A1(_03773_),
    .A2(_04020_),
    .B1(_04028_),
    .B2(_04031_),
    .Y(_04036_));
 sky130_fd_sc_hd__a2bb2oi_1 _14540_ (.A1_N(_03622_),
    .A2_N(_04019_),
    .B1(_04022_),
    .B2(_04032_),
    .Y(_04037_));
 sky130_fd_sc_hd__o21ai_4 _14541_ (.A1(_03622_),
    .A2(_04019_),
    .B1(_04036_),
    .Y(_04038_));
 sky130_fd_sc_hd__o211a_1 _14542_ (.A1(_03622_),
    .A2(_04019_),
    .B1(_04035_),
    .C1(_04036_),
    .X(_04039_));
 sky130_fd_sc_hd__a2bb2oi_2 _14543_ (.A1_N(_03624_),
    .A2_N(_04018_),
    .B1(_04035_),
    .B2(_04036_),
    .Y(_04040_));
 sky130_fd_sc_hd__a2bb2o_1 _14544_ (.A1_N(_03624_),
    .A2_N(_04018_),
    .B1(_04035_),
    .B2(_04036_),
    .X(_04041_));
 sky130_fd_sc_hd__a21oi_2 _14545_ (.A1(_04037_),
    .A2(_04035_),
    .B1(_04040_),
    .Y(_04042_));
 sky130_fd_sc_hd__o211a_2 _14546_ (.A1(_04038_),
    .A2(_04033_),
    .B1(_04017_),
    .C1(_04041_),
    .X(_04043_));
 sky130_fd_sc_hd__o211ai_4 _14547_ (.A1(_04038_),
    .A2(_04033_),
    .B1(_04017_),
    .C1(_04041_),
    .Y(_04044_));
 sky130_fd_sc_hd__o21bai_4 _14548_ (.A1(_04039_),
    .A2(_04040_),
    .B1_N(_04017_),
    .Y(_04046_));
 sky130_fd_sc_hd__o21ai_4 _14549_ (.A1(_03648_),
    .A2(_03649_),
    .B1(_03653_),
    .Y(_04047_));
 sky130_fd_sc_hd__o31a_1 _14550_ (.A1(_01769_),
    .A2(_02054_),
    .A3(_03649_),
    .B1(_03653_),
    .X(_04048_));
 sky130_fd_sc_hd__nand2_1 _14551_ (.A(net28),
    .B(net45),
    .Y(_04049_));
 sky130_fd_sc_hd__and4_1 _14552_ (.A(net29),
    .B(net30),
    .C(net42),
    .D(net43),
    .X(_04050_));
 sky130_fd_sc_hd__nand4_4 _14553_ (.A(net29),
    .B(net30),
    .C(net42),
    .D(net43),
    .Y(_04051_));
 sky130_fd_sc_hd__a22oi_4 _14554_ (.A1(net30),
    .A2(net42),
    .B1(net43),
    .B2(net29),
    .Y(_04052_));
 sky130_fd_sc_hd__a22o_1 _14555_ (.A1(net30),
    .A2(net42),
    .B1(net43),
    .B2(net29),
    .X(_04053_));
 sky130_fd_sc_hd__o211ai_2 _14556_ (.A1(_01748_),
    .A2(_02054_),
    .B1(_04051_),
    .C1(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__o21bai_1 _14557_ (.A1(_04050_),
    .A2(_04052_),
    .B1_N(_04049_),
    .Y(_04055_));
 sky130_fd_sc_hd__o22ai_4 _14558_ (.A1(_01748_),
    .A2(_02054_),
    .B1(_04050_),
    .B2(_04052_),
    .Y(_04057_));
 sky130_fd_sc_hd__nand4_4 _14559_ (.A(_04053_),
    .B(net45),
    .C(net28),
    .D(_04051_),
    .Y(_04058_));
 sky130_fd_sc_hd__a21oi_1 _14560_ (.A1(_04057_),
    .A2(_04058_),
    .B1(_04047_),
    .Y(_04059_));
 sky130_fd_sc_hd__a21o_1 _14561_ (.A1(_04057_),
    .A2(_04058_),
    .B1(_04047_),
    .X(_04060_));
 sky130_fd_sc_hd__nand3_4 _14562_ (.A(_04057_),
    .B(_04058_),
    .C(_04047_),
    .Y(_04061_));
 sky130_fd_sc_hd__nand2_1 _14563_ (.A(net23),
    .B(net48),
    .Y(_04062_));
 sky130_fd_sc_hd__nand2_1 _14564_ (.A(net27),
    .B(net47),
    .Y(_04063_));
 sky130_fd_sc_hd__and4_1 _14565_ (.A(net27),
    .B(net26),
    .C(net46),
    .D(net47),
    .X(_04064_));
 sky130_fd_sc_hd__nand4_4 _14566_ (.A(net27),
    .B(net26),
    .C(net46),
    .D(net47),
    .Y(_04065_));
 sky130_fd_sc_hd__a22oi_2 _14567_ (.A1(net27),
    .A2(net46),
    .B1(net47),
    .B2(net26),
    .Y(_04066_));
 sky130_fd_sc_hd__a22o_1 _14568_ (.A1(net27),
    .A2(net46),
    .B1(net47),
    .B2(net26),
    .X(_04068_));
 sky130_fd_sc_hd__o2bb2ai_4 _14569_ (.A1_N(_04065_),
    .A2_N(_04068_),
    .B1(_01802_),
    .B2(_02109_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand4_4 _14570_ (.A(_04068_),
    .B(net48),
    .C(net23),
    .D(_04065_),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_2 _14571_ (.A(_04069_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__and4_2 _14572_ (.A(_04060_),
    .B(_04061_),
    .C(_04069_),
    .D(_04070_),
    .X(_04072_));
 sky130_fd_sc_hd__a22oi_4 _14573_ (.A1(_04060_),
    .A2(_04061_),
    .B1(_04069_),
    .B2(_04070_),
    .Y(_04073_));
 sky130_fd_sc_hd__a21oi_4 _14574_ (.A1(_04060_),
    .A2(_04061_),
    .B1(_04071_),
    .Y(_04074_));
 sky130_fd_sc_hd__and3_2 _14575_ (.A(_04060_),
    .B(_04061_),
    .C(_04071_),
    .X(_04075_));
 sky130_fd_sc_hd__o211ai_4 _14576_ (.A1(_04072_),
    .A2(_04073_),
    .B1(_04044_),
    .C1(_04046_),
    .Y(_04076_));
 sky130_fd_sc_hd__o2bb2ai_2 _14577_ (.A1_N(_04044_),
    .A2_N(_04046_),
    .B1(_04074_),
    .B2(_04075_),
    .Y(_04077_));
 sky130_fd_sc_hd__o2bb2ai_2 _14578_ (.A1_N(_04044_),
    .A2_N(_04046_),
    .B1(_04072_),
    .B2(_04073_),
    .Y(_04079_));
 sky130_fd_sc_hd__o22a_2 _14579_ (.A1(_04074_),
    .A2(_04075_),
    .B1(_04017_),
    .B2(_04042_),
    .X(_04080_));
 sky130_fd_sc_hd__o22ai_4 _14580_ (.A1(_04074_),
    .A2(_04075_),
    .B1(_04017_),
    .B2(_04042_),
    .Y(_04081_));
 sky130_fd_sc_hd__o221a_1 _14581_ (.A1(_04074_),
    .A2(_04075_),
    .B1(_04017_),
    .B2(_04042_),
    .C1(_04044_),
    .X(_04082_));
 sky130_fd_sc_hd__nand3_1 _14582_ (.A(_04077_),
    .B(_04016_),
    .C(_04076_),
    .Y(_04083_));
 sky130_fd_sc_hd__o21ai_1 _14583_ (.A1(_03803_),
    .A2(_03810_),
    .B1(_04079_),
    .Y(_04084_));
 sky130_fd_sc_hd__o221a_2 _14584_ (.A1(_04043_),
    .A2(_04081_),
    .B1(_03803_),
    .B2(_03810_),
    .C1(_04079_),
    .X(_04085_));
 sky130_fd_sc_hd__o221ai_4 _14585_ (.A1(_04043_),
    .A2(_04081_),
    .B1(_03803_),
    .B2(_03810_),
    .C1(_04079_),
    .Y(_04086_));
 sky130_fd_sc_hd__a21oi_2 _14586_ (.A1(_04083_),
    .A2(_04086_),
    .B1(_04014_),
    .Y(_04087_));
 sky130_fd_sc_hd__a21o_1 _14587_ (.A1(_04083_),
    .A2(_04086_),
    .B1(_04014_),
    .X(_04088_));
 sky130_fd_sc_hd__a31oi_4 _14588_ (.A1(_04077_),
    .A2(_04016_),
    .A3(_04076_),
    .B1(_04013_),
    .Y(_04090_));
 sky130_fd_sc_hd__a31o_2 _14589_ (.A1(_04077_),
    .A2(_04016_),
    .A3(_04076_),
    .B1(_04013_),
    .X(_04091_));
 sky130_fd_sc_hd__o21ai_2 _14590_ (.A1(_04082_),
    .A2(_04084_),
    .B1(_04090_),
    .Y(_04092_));
 sky130_fd_sc_hd__inv_2 _14591_ (.A(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__a21oi_1 _14592_ (.A1(_04086_),
    .A2(_04090_),
    .B1(_04087_),
    .Y(_04094_));
 sky130_fd_sc_hd__o21ai_1 _14593_ (.A1(_04085_),
    .A2(_04091_),
    .B1(_04088_),
    .Y(_04095_));
 sky130_fd_sc_hd__o2bb2ai_4 _14594_ (.A1_N(_04009_),
    .A2_N(_04011_),
    .B1(_04087_),
    .B2(_04093_),
    .Y(_04096_));
 sky130_fd_sc_hd__nand3_4 _14595_ (.A(_04011_),
    .B(_04088_),
    .C(_04092_),
    .Y(_04097_));
 sky130_fd_sc_hd__o2111ai_4 _14596_ (.A1(_04085_),
    .A2(_04091_),
    .B1(_04088_),
    .C1(_04009_),
    .D1(_04011_),
    .Y(_04098_));
 sky130_fd_sc_hd__a22oi_4 _14597_ (.A1(_03822_),
    .A2(_03874_),
    .B1(_04096_),
    .B2(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__a22o_1 _14598_ (.A1(_03822_),
    .A2(_03874_),
    .B1(_04096_),
    .B2(_04098_),
    .X(_04101_));
 sky130_fd_sc_hd__o211a_1 _14599_ (.A1(_04008_),
    .A2(_04097_),
    .B1(_03875_),
    .C1(_04096_),
    .X(_04102_));
 sky130_fd_sc_hd__o211ai_4 _14600_ (.A1(_04008_),
    .A2(_04097_),
    .B1(_03875_),
    .C1(_04096_),
    .Y(_04103_));
 sky130_fd_sc_hd__o21ai_2 _14601_ (.A1(_03663_),
    .A2(_03664_),
    .B1(_03666_),
    .Y(_04104_));
 sky130_fd_sc_hd__inv_2 _14602_ (.A(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__nand2_1 _14603_ (.A(net12),
    .B(net50),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_4 _14604_ (.A(net12),
    .B(net49),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _14605_ (.A(net1),
    .B(net50),
    .Y(_04108_));
 sky130_fd_sc_hd__and4_1 _14606_ (.A(net12),
    .B(net1),
    .C(net49),
    .D(net50),
    .X(_04109_));
 sky130_fd_sc_hd__nand4_1 _14607_ (.A(net12),
    .B(net1),
    .C(net49),
    .D(net50),
    .Y(_04110_));
 sky130_fd_sc_hd__o21a_1 _14608_ (.A1(_01824_),
    .A2(_02120_),
    .B1(_04108_),
    .X(_04112_));
 sky130_fd_sc_hd__a22o_1 _14609_ (.A1(net12),
    .A2(net49),
    .B1(net50),
    .B2(net1),
    .X(_04113_));
 sky130_fd_sc_hd__a31o_1 _14610_ (.A1(net12),
    .A2(net50),
    .A3(_03594_),
    .B1(_04112_),
    .X(_04114_));
 sky130_fd_sc_hd__o311a_1 _14611_ (.A1(_01846_),
    .A2(_02120_),
    .A3(_04106_),
    .B1(_04113_),
    .C1(_04104_),
    .X(_04115_));
 sky130_fd_sc_hd__nand3_1 _14612_ (.A(_04104_),
    .B(_04110_),
    .C(_04113_),
    .Y(_04116_));
 sky130_fd_sc_hd__a21o_1 _14613_ (.A1(_04110_),
    .A2(_04113_),
    .B1(_04104_),
    .X(_04117_));
 sky130_fd_sc_hd__o21a_1 _14614_ (.A1(_04109_),
    .A2(_04112_),
    .B1(_04104_),
    .X(_04118_));
 sky130_fd_sc_hd__and4_1 _14615_ (.A(_03666_),
    .B(_03668_),
    .C(_04110_),
    .D(_04113_),
    .X(_04119_));
 sky130_fd_sc_hd__nand2_1 _14616_ (.A(_04116_),
    .B(_04117_),
    .Y(_04120_));
 sky130_fd_sc_hd__o22ai_2 _14617_ (.A1(_03656_),
    .A2(_03660_),
    .B1(_03669_),
    .B2(_03658_),
    .Y(_04121_));
 sky130_fd_sc_hd__o211a_1 _14618_ (.A1(_03669_),
    .A2(_03658_),
    .B1(_03662_),
    .C1(_04120_),
    .X(_04123_));
 sky130_fd_sc_hd__o211ai_2 _14619_ (.A1(_03669_),
    .A2(_03658_),
    .B1(_03662_),
    .C1(_04120_),
    .Y(_04124_));
 sky130_fd_sc_hd__o21ai_4 _14620_ (.A1(_04118_),
    .A2(_04119_),
    .B1(_04121_),
    .Y(_04125_));
 sky130_fd_sc_hd__a32o_2 _14621_ (.A1(net1),
    .A2(_03595_),
    .A3(net49),
    .B1(_04125_),
    .B2(_04124_),
    .X(_04126_));
 sky130_fd_sc_hd__o211a_1 _14622_ (.A1(_03362_),
    .A2(_03364_),
    .B1(_04124_),
    .C1(_04125_),
    .X(_04127_));
 sky130_fd_sc_hd__o2111ai_2 _14623_ (.A1(_03362_),
    .A2(_03364_),
    .B1(_03594_),
    .C1(_04124_),
    .D1(_04125_),
    .Y(_04128_));
 sky130_fd_sc_hd__a21oi_1 _14624_ (.A1(_04126_),
    .A2(_04128_),
    .B1(_03599_),
    .Y(_04129_));
 sky130_fd_sc_hd__a32o_1 _14625_ (.A1(_03593_),
    .A2(_03596_),
    .A3(_03597_),
    .B1(_04126_),
    .B2(_04128_),
    .X(_04130_));
 sky130_fd_sc_hd__and4_1 _14626_ (.A(_03593_),
    .B(_03596_),
    .C(_03597_),
    .D(_04126_),
    .X(_04131_));
 sky130_fd_sc_hd__nand2_1 _14627_ (.A(_04126_),
    .B(_03599_),
    .Y(_04132_));
 sky130_fd_sc_hd__a21oi_1 _14628_ (.A1(_03599_),
    .A2(_04126_),
    .B1(_04129_),
    .Y(_04134_));
 sky130_fd_sc_hd__a21o_1 _14629_ (.A1(_03599_),
    .A2(_04126_),
    .B1(_04129_),
    .X(_04135_));
 sky130_fd_sc_hd__o22ai_2 _14630_ (.A1(_03676_),
    .A2(_03680_),
    .B1(_03684_),
    .B2(_03678_),
    .Y(_04136_));
 sky130_fd_sc_hd__and3_1 _14631_ (.A(_04130_),
    .B(_04132_),
    .C(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__nand2_1 _14632_ (.A(_04136_),
    .B(_04134_),
    .Y(_04138_));
 sky130_fd_sc_hd__o211ai_4 _14633_ (.A1(_03678_),
    .A2(_03684_),
    .B1(_04135_),
    .C1(_03682_),
    .Y(_04139_));
 sky130_fd_sc_hd__inv_2 _14634_ (.A(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__a22oi_1 _14635_ (.A1(_03549_),
    .A2(_03601_),
    .B1(_04138_),
    .B2(_04139_),
    .Y(_04141_));
 sky130_fd_sc_hd__a22o_1 _14636_ (.A1(_03549_),
    .A2(_03601_),
    .B1(_04138_),
    .B2(_04139_),
    .X(_04142_));
 sky130_fd_sc_hd__nand4_2 _14637_ (.A(_04138_),
    .B(_04139_),
    .C(_03549_),
    .D(_03601_),
    .Y(_04143_));
 sky130_fd_sc_hd__a21boi_1 _14638_ (.A1(_04136_),
    .A2(_04134_),
    .B1_N(_03602_),
    .Y(_04145_));
 sky130_fd_sc_hd__a21oi_1 _14639_ (.A1(_04139_),
    .A2(_04145_),
    .B1(_04141_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_2 _14640_ (.A(_04142_),
    .B(_04143_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand4_2 _14641_ (.A(_04101_),
    .B(_04103_),
    .C(_04142_),
    .D(_04143_),
    .Y(_04148_));
 sky130_fd_sc_hd__o21bai_2 _14642_ (.A1(_04099_),
    .A2(_04102_),
    .B1_N(_04146_),
    .Y(_04149_));
 sky130_fd_sc_hd__o21bai_4 _14643_ (.A1(_04099_),
    .A2(_04102_),
    .B1_N(_04147_),
    .Y(_04150_));
 sky130_fd_sc_hd__nand3_4 _14644_ (.A(_04101_),
    .B(_04103_),
    .C(_04147_),
    .Y(_04151_));
 sky130_fd_sc_hd__a21oi_4 _14645_ (.A1(_03832_),
    .A2(_03611_),
    .B1(_03833_),
    .Y(_04152_));
 sky130_fd_sc_hd__nand3_2 _14646_ (.A(_04150_),
    .B(_04151_),
    .C(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__a21oi_4 _14647_ (.A1(_04150_),
    .A2(_04151_),
    .B1(_04152_),
    .Y(_04154_));
 sky130_fd_sc_hd__o211ai_4 _14648_ (.A1(_03833_),
    .A2(_03836_),
    .B1(_04148_),
    .C1(_04149_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _14649_ (.A(_04153_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__o2bb2ai_1 _14650_ (.A1_N(_04153_),
    .A2_N(_04156_),
    .B1(_03592_),
    .B2(_03605_),
    .Y(_04158_));
 sky130_fd_sc_hd__a31oi_2 _14651_ (.A1(_04150_),
    .A2(_04151_),
    .A3(_04152_),
    .B1(_03610_),
    .Y(_04159_));
 sky130_fd_sc_hd__a31o_1 _14652_ (.A1(_04150_),
    .A2(_04151_),
    .A3(_04152_),
    .B1(_03610_),
    .X(_04160_));
 sky130_fd_sc_hd__nand3_1 _14653_ (.A(_04156_),
    .B(_03609_),
    .C(_04153_),
    .Y(_04161_));
 sky130_fd_sc_hd__a21o_1 _14654_ (.A1(_04153_),
    .A2(_04156_),
    .B1(_03610_),
    .X(_04162_));
 sky130_fd_sc_hd__o211ai_1 _14655_ (.A1(_03592_),
    .A2(_03605_),
    .B1(_04153_),
    .C1(_04156_),
    .Y(_04163_));
 sky130_fd_sc_hd__o21ai_1 _14656_ (.A1(_04154_),
    .A2(_04160_),
    .B1(_04158_),
    .Y(_04164_));
 sky130_fd_sc_hd__a21oi_1 _14657_ (.A1(_04158_),
    .A2(_04161_),
    .B1(_03873_),
    .Y(_04165_));
 sky130_fd_sc_hd__nand3_1 _14658_ (.A(_04162_),
    .B(_04163_),
    .C(_03872_),
    .Y(_04167_));
 sky130_fd_sc_hd__a2bb2oi_2 _14659_ (.A1_N(_03843_),
    .A2_N(_03847_),
    .B1(_04157_),
    .B2(_03610_),
    .Y(_04168_));
 sky130_fd_sc_hd__o221a_1 _14660_ (.A1(_03843_),
    .A2(_03847_),
    .B1(_04154_),
    .B2(_04160_),
    .C1(_04158_),
    .X(_04169_));
 sky130_fd_sc_hd__a21oi_1 _14661_ (.A1(_04161_),
    .A2(_04168_),
    .B1(_04165_),
    .Y(_04170_));
 sky130_fd_sc_hd__o22ai_1 _14662_ (.A1(_03852_),
    .A2(_03851_),
    .B1(_04169_),
    .B2(_04165_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand2_1 _14663_ (.A(_03856_),
    .B(_04167_),
    .Y(_04172_));
 sky130_fd_sc_hd__o21a_1 _14664_ (.A1(_04169_),
    .A2(_04172_),
    .B1(_04171_),
    .X(_04173_));
 sky130_fd_sc_hd__o21ai_1 _14665_ (.A1(_04169_),
    .A2(_04172_),
    .B1(_04171_),
    .Y(_04174_));
 sky130_fd_sc_hd__a22o_1 _14666_ (.A1(_03857_),
    .A2(_03860_),
    .B1(_03871_),
    .B2(_03858_),
    .X(_04175_));
 sky130_fd_sc_hd__xor2_1 _14667_ (.A(_04173_),
    .B(_04175_),
    .X(net82));
 sky130_fd_sc_hd__a31oi_2 _14668_ (.A1(_03875_),
    .A2(_04096_),
    .A3(_04098_),
    .B1(_04146_),
    .Y(_04177_));
 sky130_fd_sc_hd__a21oi_2 _14669_ (.A1(_04103_),
    .A2(_04147_),
    .B1(_04099_),
    .Y(_04178_));
 sky130_fd_sc_hd__a32oi_4 _14670_ (.A1(_04057_),
    .A2(_04058_),
    .A3(_04047_),
    .B1(_04069_),
    .B2(_04070_),
    .Y(_04179_));
 sky130_fd_sc_hd__a32oi_4 _14671_ (.A1(_04048_),
    .A2(_04054_),
    .A3(_04055_),
    .B1(_04061_),
    .B2(_04071_),
    .Y(_04180_));
 sky130_fd_sc_hd__nor2_1 _14672_ (.A(_04062_),
    .B(_04066_),
    .Y(_04181_));
 sky130_fd_sc_hd__o21ai_1 _14673_ (.A1(_04062_),
    .A2(_04066_),
    .B1(_04065_),
    .Y(_04182_));
 sky130_fd_sc_hd__o21a_1 _14674_ (.A1(_04062_),
    .A2(_04066_),
    .B1(_04065_),
    .X(_04183_));
 sky130_fd_sc_hd__and2_1 _14675_ (.A(net1),
    .B(net51),
    .X(_04184_));
 sky130_fd_sc_hd__nand2_4 _14676_ (.A(net23),
    .B(net50),
    .Y(_04185_));
 sky130_fd_sc_hd__nand2_1 _14677_ (.A(net23),
    .B(net49),
    .Y(_04186_));
 sky130_fd_sc_hd__a22oi_4 _14678_ (.A1(net23),
    .A2(net49),
    .B1(net50),
    .B2(net12),
    .Y(_04188_));
 sky130_fd_sc_hd__a22o_1 _14679_ (.A1(net23),
    .A2(net49),
    .B1(net50),
    .B2(net12),
    .X(_04189_));
 sky130_fd_sc_hd__o2bb2ai_1 _14680_ (.A1_N(_04106_),
    .A2_N(_04186_),
    .B1(_04185_),
    .B2(_04107_),
    .Y(_04190_));
 sky130_fd_sc_hd__o221ai_4 _14681_ (.A1(_01846_),
    .A2(_02152_),
    .B1(_04107_),
    .B2(_04185_),
    .C1(_04189_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_1 _14682_ (.A(_04190_),
    .B(_04184_),
    .Y(_04192_));
 sky130_fd_sc_hd__o2111ai_2 _14683_ (.A1(_04107_),
    .A2(_04185_),
    .B1(net1),
    .C1(net51),
    .D1(_04189_),
    .Y(_04193_));
 sky130_fd_sc_hd__o21ai_1 _14684_ (.A1(_01846_),
    .A2(_02152_),
    .B1(_04190_),
    .Y(_04194_));
 sky130_fd_sc_hd__a2bb2oi_2 _14685_ (.A1_N(_04064_),
    .A2_N(_04181_),
    .B1(_04191_),
    .B2(_04192_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand3_2 _14686_ (.A(_04194_),
    .B(_04182_),
    .C(_04193_),
    .Y(_04196_));
 sky130_fd_sc_hd__a21oi_1 _14687_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04182_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand3_2 _14688_ (.A(_04183_),
    .B(_04191_),
    .C(_04192_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _14689_ (.A(_04199_),
    .B(_04109_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand3_1 _14690_ (.A(_04199_),
    .B(_04109_),
    .C(_04196_),
    .Y(_04201_));
 sky130_fd_sc_hd__o2bb2ai_2 _14691_ (.A1_N(_04196_),
    .A2_N(_04199_),
    .B1(_04107_),
    .B2(_04108_),
    .Y(_04202_));
 sky130_fd_sc_hd__o21ai_1 _14692_ (.A1(_04195_),
    .A2(_04197_),
    .B1(_04109_),
    .Y(_04203_));
 sky130_fd_sc_hd__o211ai_1 _14693_ (.A1(_04107_),
    .A2(_04108_),
    .B1(_04196_),
    .C1(_04199_),
    .Y(_04204_));
 sky130_fd_sc_hd__o211a_1 _14694_ (.A1(_04195_),
    .A2(_04200_),
    .B1(_04180_),
    .C1(_04202_),
    .X(_04205_));
 sky130_fd_sc_hd__o211ai_2 _14695_ (.A1(_04195_),
    .A2(_04200_),
    .B1(_04180_),
    .C1(_04202_),
    .Y(_04206_));
 sky130_fd_sc_hd__a2bb2oi_2 _14696_ (.A1_N(_04059_),
    .A2_N(_04179_),
    .B1(_04201_),
    .B2(_04202_),
    .Y(_04207_));
 sky130_fd_sc_hd__o211ai_1 _14697_ (.A1(_04059_),
    .A2(_04179_),
    .B1(_04203_),
    .C1(_04204_),
    .Y(_04208_));
 sky130_fd_sc_hd__o22ai_4 _14698_ (.A1(_04114_),
    .A2(_04105_),
    .B1(_04207_),
    .B2(_04205_),
    .Y(_04210_));
 sky130_fd_sc_hd__nor2_1 _14699_ (.A(_04116_),
    .B(_04207_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand3_2 _14700_ (.A(_04208_),
    .B(_04115_),
    .C(_04206_),
    .Y(_04212_));
 sky130_fd_sc_hd__o21ai_2 _14701_ (.A1(_03596_),
    .A2(_04123_),
    .B1(_04125_),
    .Y(_04213_));
 sky130_fd_sc_hd__a22oi_1 _14702_ (.A1(_03594_),
    .A2(_04127_),
    .B1(_04210_),
    .B2(_04212_),
    .Y(_04214_));
 sky130_fd_sc_hd__a21oi_2 _14703_ (.A1(_04210_),
    .A2(_04212_),
    .B1(_04213_),
    .Y(_04215_));
 sky130_fd_sc_hd__and3_4 _14704_ (.A(_04210_),
    .B(_04212_),
    .C(_04213_),
    .X(_04216_));
 sky130_fd_sc_hd__nand3_2 _14705_ (.A(_04210_),
    .B(_04212_),
    .C(_04213_),
    .Y(_04217_));
 sky130_fd_sc_hd__a21boi_2 _14706_ (.A1(_04214_),
    .A2(_04125_),
    .B1_N(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__o2bb2ai_1 _14707_ (.A1_N(_04014_),
    .A2_N(_04083_),
    .B1(_04084_),
    .B2(_04082_),
    .Y(_04219_));
 sky130_fd_sc_hd__o21a_1 _14708_ (.A1(_04085_),
    .A2(_04090_),
    .B1(_04218_),
    .X(_04221_));
 sky130_fd_sc_hd__o21ai_2 _14709_ (.A1(_04085_),
    .A2(_04090_),
    .B1(_04218_),
    .Y(_04222_));
 sky130_fd_sc_hd__o211a_1 _14710_ (.A1(_04215_),
    .A2(_04216_),
    .B1(_04086_),
    .C1(_04091_),
    .X(_04223_));
 sky130_fd_sc_hd__o211ai_4 _14711_ (.A1(_04215_),
    .A2(_04216_),
    .B1(_04086_),
    .C1(_04091_),
    .Y(_04224_));
 sky130_fd_sc_hd__a22oi_4 _14712_ (.A1(_03599_),
    .A2(_04126_),
    .B1(_04222_),
    .B2(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__a22o_1 _14713_ (.A1(_03599_),
    .A2(_04126_),
    .B1(_04222_),
    .B2(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__a21oi_1 _14714_ (.A1(_04219_),
    .A2(_04218_),
    .B1(_04132_),
    .Y(_04227_));
 sky130_fd_sc_hd__a21o_1 _14715_ (.A1(_04219_),
    .A2(_04218_),
    .B1(_04132_),
    .X(_04228_));
 sky130_fd_sc_hd__and3_2 _14716_ (.A(_04222_),
    .B(_04224_),
    .C(_04131_),
    .X(_04229_));
 sky130_fd_sc_hd__a21oi_1 _14717_ (.A1(_04224_),
    .A2(_04227_),
    .B1(_04225_),
    .Y(_04230_));
 sky130_fd_sc_hd__o21ai_2 _14718_ (.A1(_04223_),
    .A2(_04228_),
    .B1(_04226_),
    .Y(_04232_));
 sky130_fd_sc_hd__o2bb2ai_4 _14719_ (.A1_N(_04003_),
    .A2_N(_04007_),
    .B1(_04095_),
    .B2(_04010_),
    .Y(_04233_));
 sky130_fd_sc_hd__a22oi_4 _14720_ (.A1(_04003_),
    .A2(_04007_),
    .B1(_04094_),
    .B2(_04011_),
    .Y(_04234_));
 sky130_fd_sc_hd__o22ai_4 _14721_ (.A1(_03905_),
    .A2(_03909_),
    .B1(_03911_),
    .B2(_03907_),
    .Y(_04235_));
 sky130_fd_sc_hd__o21ai_2 _14722_ (.A1(_04049_),
    .A2(_04052_),
    .B1(_04051_),
    .Y(_04236_));
 sky130_fd_sc_hd__nand2_1 _14723_ (.A(net29),
    .B(net45),
    .Y(_04237_));
 sky130_fd_sc_hd__and4_1 _14724_ (.A(net30),
    .B(net31),
    .C(net42),
    .D(net43),
    .X(_04238_));
 sky130_fd_sc_hd__nand4_2 _14725_ (.A(net30),
    .B(net31),
    .C(net42),
    .D(net43),
    .Y(_04239_));
 sky130_fd_sc_hd__a22oi_4 _14726_ (.A1(net31),
    .A2(net42),
    .B1(net43),
    .B2(net30),
    .Y(_04240_));
 sky130_fd_sc_hd__a22o_1 _14727_ (.A1(net31),
    .A2(net42),
    .B1(net43),
    .B2(net30),
    .X(_04241_));
 sky130_fd_sc_hd__o211ai_1 _14728_ (.A1(_01857_),
    .A2(_02054_),
    .B1(_04239_),
    .C1(_04241_),
    .Y(_04243_));
 sky130_fd_sc_hd__o21bai_1 _14729_ (.A1(_04238_),
    .A2(_04240_),
    .B1_N(_04237_),
    .Y(_04244_));
 sky130_fd_sc_hd__a22o_1 _14730_ (.A1(net29),
    .A2(net45),
    .B1(_04239_),
    .B2(_04241_),
    .X(_04245_));
 sky130_fd_sc_hd__a41o_1 _14731_ (.A1(net30),
    .A2(net31),
    .A3(net42),
    .A4(net43),
    .B1(_04237_),
    .X(_04246_));
 sky130_fd_sc_hd__nand3b_2 _14732_ (.A_N(_04236_),
    .B(_04243_),
    .C(_04244_),
    .Y(_04247_));
 sky130_fd_sc_hd__o211a_1 _14733_ (.A1(_04240_),
    .A2(_04246_),
    .B1(_04236_),
    .C1(_04245_),
    .X(_04248_));
 sky130_fd_sc_hd__o211ai_2 _14734_ (.A1(_04240_),
    .A2(_04246_),
    .B1(_04236_),
    .C1(_04245_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_1 _14735_ (.A(net26),
    .B(net48),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2_2 _14736_ (.A(net28),
    .B(net46),
    .Y(_04251_));
 sky130_fd_sc_hd__a22oi_4 _14737_ (.A1(net28),
    .A2(net46),
    .B1(net47),
    .B2(net27),
    .Y(_04252_));
 sky130_fd_sc_hd__and4_2 _14738_ (.A(net28),
    .B(net27),
    .C(net46),
    .D(net47),
    .X(_04253_));
 sky130_fd_sc_hd__a211oi_1 _14739_ (.A1(net26),
    .A2(net48),
    .B1(_04252_),
    .C1(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__a211o_1 _14740_ (.A1(net26),
    .A2(net48),
    .B1(_04252_),
    .C1(_04253_),
    .X(_04255_));
 sky130_fd_sc_hd__o211a_1 _14741_ (.A1(_04252_),
    .A2(_04253_),
    .B1(net26),
    .C1(net48),
    .X(_04256_));
 sky130_fd_sc_hd__o211ai_1 _14742_ (.A1(_04252_),
    .A2(_04253_),
    .B1(net26),
    .C1(net48),
    .Y(_04257_));
 sky130_fd_sc_hd__nand2_1 _14743_ (.A(_04255_),
    .B(_04257_),
    .Y(_04258_));
 sky130_fd_sc_hd__o21a_1 _14744_ (.A1(_04254_),
    .A2(_04256_),
    .B1(_04247_),
    .X(_04259_));
 sky130_fd_sc_hd__and3_1 _14745_ (.A(_04247_),
    .B(_04249_),
    .C(_04258_),
    .X(_04260_));
 sky130_fd_sc_hd__a21oi_2 _14746_ (.A1(_04247_),
    .A2(_04249_),
    .B1(_04258_),
    .Y(_04261_));
 sky130_fd_sc_hd__and4_1 _14747_ (.A(_04247_),
    .B(_04249_),
    .C(_04255_),
    .D(_04257_),
    .X(_04262_));
 sky130_fd_sc_hd__o2bb2a_1 _14748_ (.A1_N(_04247_),
    .A2_N(_04249_),
    .B1(_04254_),
    .B2(_04256_),
    .X(_04264_));
 sky130_fd_sc_hd__a21oi_1 _14749_ (.A1(_04259_),
    .A2(_04249_),
    .B1(_04261_),
    .Y(_04265_));
 sky130_fd_sc_hd__o21ai_2 _14750_ (.A1(_04022_),
    .A2(_04032_),
    .B1(_04038_),
    .Y(_04266_));
 sky130_fd_sc_hd__o21a_1 _14751_ (.A1(_01879_),
    .A2(_02010_),
    .B1(_04025_),
    .X(_04267_));
 sky130_fd_sc_hd__a31o_1 _14752_ (.A1(_04027_),
    .A2(net41),
    .A3(net31),
    .B1(_04024_),
    .X(_04268_));
 sky130_fd_sc_hd__o31a_1 _14753_ (.A1(_01879_),
    .A2(_02010_),
    .A3(_04026_),
    .B1(_04025_),
    .X(_04269_));
 sky130_fd_sc_hd__o21ai_2 _14754_ (.A1(_03893_),
    .A2(_03894_),
    .B1(_03896_),
    .Y(_04270_));
 sky130_fd_sc_hd__o21a_1 _14755_ (.A1(_03893_),
    .A2(_03894_),
    .B1(_03896_),
    .X(_04271_));
 sky130_fd_sc_hd__nand2_1 _14756_ (.A(net32),
    .B(net41),
    .Y(_04272_));
 sky130_fd_sc_hd__nand2_2 _14757_ (.A(net3),
    .B(net39),
    .Y(_04273_));
 sky130_fd_sc_hd__a22oi_4 _14758_ (.A1(net3),
    .A2(net39),
    .B1(net40),
    .B2(net2),
    .Y(_04275_));
 sky130_fd_sc_hd__a22o_1 _14759_ (.A1(net3),
    .A2(net39),
    .B1(net40),
    .B2(net2),
    .X(_04276_));
 sky130_fd_sc_hd__nand2_1 _14760_ (.A(net3),
    .B(net40),
    .Y(_04277_));
 sky130_fd_sc_hd__and4_2 _14761_ (.A(net2),
    .B(net3),
    .C(net39),
    .D(net40),
    .X(_04278_));
 sky130_fd_sc_hd__nand4_4 _14762_ (.A(net2),
    .B(net3),
    .C(net39),
    .D(net40),
    .Y(_04279_));
 sky130_fd_sc_hd__o211ai_2 _14763_ (.A1(_01912_),
    .A2(_02010_),
    .B1(_04276_),
    .C1(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__o21bai_2 _14764_ (.A1(_04275_),
    .A2(_04278_),
    .B1_N(_04272_),
    .Y(_04281_));
 sky130_fd_sc_hd__o22ai_4 _14765_ (.A1(_01912_),
    .A2(_02010_),
    .B1(_04275_),
    .B2(_04278_),
    .Y(_04282_));
 sky130_fd_sc_hd__a41o_1 _14766_ (.A1(net2),
    .A2(net3),
    .A3(net39),
    .A4(net40),
    .B1(_04272_),
    .X(_04283_));
 sky130_fd_sc_hd__nand4_1 _14767_ (.A(_04276_),
    .B(_04279_),
    .C(net32),
    .D(net41),
    .Y(_04284_));
 sky130_fd_sc_hd__o211a_1 _14768_ (.A1(_04275_),
    .A2(_04283_),
    .B1(_04270_),
    .C1(_04282_),
    .X(_04286_));
 sky130_fd_sc_hd__o211ai_4 _14769_ (.A1(_04275_),
    .A2(_04283_),
    .B1(_04270_),
    .C1(_04282_),
    .Y(_04287_));
 sky130_fd_sc_hd__a21oi_1 _14770_ (.A1(_04282_),
    .A2(_04284_),
    .B1(_04270_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand3_1 _14771_ (.A(_04271_),
    .B(_04280_),
    .C(_04281_),
    .Y(_04289_));
 sky130_fd_sc_hd__a31oi_4 _14772_ (.A1(_04271_),
    .A2(_04280_),
    .A3(_04281_),
    .B1(_04269_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _14773_ (.A(_04290_),
    .B(_04287_),
    .Y(_04291_));
 sky130_fd_sc_hd__a2bb2oi_2 _14774_ (.A1_N(_04026_),
    .A2_N(_04267_),
    .B1(_04287_),
    .B2(_04289_),
    .Y(_04292_));
 sky130_fd_sc_hd__o22ai_2 _14775_ (.A1(_04026_),
    .A2(_04267_),
    .B1(_04286_),
    .B2(_04288_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21oi_1 _14776_ (.A1(_04287_),
    .A2(_04290_),
    .B1(_04292_),
    .Y(_04294_));
 sky130_fd_sc_hd__a221oi_4 _14777_ (.A1(_04290_),
    .A2(_04287_),
    .B1(_04038_),
    .B2(_04035_),
    .C1(_04292_),
    .Y(_04295_));
 sky130_fd_sc_hd__a221o_1 _14778_ (.A1(_04290_),
    .A2(_04287_),
    .B1(_04038_),
    .B2(_04035_),
    .C1(_04292_),
    .X(_04297_));
 sky130_fd_sc_hd__a21oi_2 _14779_ (.A1(_04291_),
    .A2(_04293_),
    .B1(_04266_),
    .Y(_04298_));
 sky130_fd_sc_hd__a21o_1 _14780_ (.A1(_04291_),
    .A2(_04293_),
    .B1(_04266_),
    .X(_04299_));
 sky130_fd_sc_hd__o21ai_1 _14781_ (.A1(_04266_),
    .A2(_04294_),
    .B1(_04265_),
    .Y(_04300_));
 sky130_fd_sc_hd__and3_2 _14782_ (.A(_04299_),
    .B(_04265_),
    .C(_04297_),
    .X(_04301_));
 sky130_fd_sc_hd__o211ai_2 _14783_ (.A1(_04262_),
    .A2(_04264_),
    .B1(_04297_),
    .C1(_04299_),
    .Y(_04302_));
 sky130_fd_sc_hd__o22ai_4 _14784_ (.A1(_04260_),
    .A2(_04261_),
    .B1(_04295_),
    .B2(_04298_),
    .Y(_04303_));
 sky130_fd_sc_hd__nand2_2 _14785_ (.A(_04235_),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__o211a_2 _14786_ (.A1(_04295_),
    .A2(_04300_),
    .B1(_04303_),
    .C1(_04235_),
    .X(_04305_));
 sky130_fd_sc_hd__a21oi_4 _14787_ (.A1(_04302_),
    .A2(_04303_),
    .B1(_04235_),
    .Y(_04306_));
 sky130_fd_sc_hd__a21o_1 _14788_ (.A1(_04302_),
    .A2(_04303_),
    .B1(_04235_),
    .X(_04308_));
 sky130_fd_sc_hd__a21oi_2 _14789_ (.A1(_04017_),
    .A2(_04042_),
    .B1(_04080_),
    .Y(_04309_));
 sky130_fd_sc_hd__o22a_2 _14790_ (.A1(_04043_),
    .A2(_04080_),
    .B1(_04305_),
    .B2(_04306_),
    .X(_04310_));
 sky130_fd_sc_hd__o22ai_4 _14791_ (.A1(_04043_),
    .A2(_04080_),
    .B1(_04305_),
    .B2(_04306_),
    .Y(_04311_));
 sky130_fd_sc_hd__o211a_2 _14792_ (.A1(_04304_),
    .A2(_04301_),
    .B1(_04309_),
    .C1(_04308_),
    .X(_04312_));
 sky130_fd_sc_hd__o211ai_4 _14793_ (.A1(_04304_),
    .A2(_04301_),
    .B1(_04309_),
    .C1(_04308_),
    .Y(_04313_));
 sky130_fd_sc_hd__o21a_1 _14794_ (.A1(_04305_),
    .A2(_04306_),
    .B1(_04309_),
    .X(_04314_));
 sky130_fd_sc_hd__a21oi_2 _14795_ (.A1(_04044_),
    .A2(_04081_),
    .B1(_04306_),
    .Y(_04315_));
 sky130_fd_sc_hd__o221a_1 _14796_ (.A1(_04043_),
    .A2(_04080_),
    .B1(_04301_),
    .B2(_04304_),
    .C1(_04308_),
    .X(_04316_));
 sky130_fd_sc_hd__o21ai_4 _14797_ (.A1(_03914_),
    .A2(_03916_),
    .B1(_04000_),
    .Y(_04317_));
 sky130_fd_sc_hd__o21ai_4 _14798_ (.A1(_03994_),
    .A2(_03996_),
    .B1(_04317_),
    .Y(_04319_));
 sky130_fd_sc_hd__o21ai_4 _14799_ (.A1(_01934_),
    .A2(_01966_),
    .B1(_03885_),
    .Y(_04320_));
 sky130_fd_sc_hd__a22oi_4 _14800_ (.A1(net34),
    .A2(net8),
    .B1(net9),
    .B2(net64),
    .Y(_04321_));
 sky130_fd_sc_hd__a22o_1 _14801_ (.A1(net34),
    .A2(net8),
    .B1(net9),
    .B2(net64),
    .X(_04322_));
 sky130_fd_sc_hd__and4_2 _14802_ (.A(net64),
    .B(net34),
    .C(net8),
    .D(net9),
    .X(_04323_));
 sky130_fd_sc_hd__nand4_2 _14803_ (.A(net64),
    .B(net34),
    .C(net8),
    .D(net9),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _14804_ (.A(net35),
    .B(net7),
    .Y(_04325_));
 sky130_fd_sc_hd__o22ai_4 _14805_ (.A1(_01934_),
    .A2(_01977_),
    .B1(_04321_),
    .B2(_04323_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand3_2 _14806_ (.A(_04324_),
    .B(net7),
    .C(net35),
    .Y(_04327_));
 sky130_fd_sc_hd__nand4_2 _14807_ (.A(_04322_),
    .B(_04324_),
    .C(net35),
    .D(net7),
    .Y(_04328_));
 sky130_fd_sc_hd__a22oi_4 _14808_ (.A1(_03883_),
    .A2(_04320_),
    .B1(_04326_),
    .B2(_04328_),
    .Y(_04330_));
 sky130_fd_sc_hd__a22o_1 _14809_ (.A1(_03883_),
    .A2(_04320_),
    .B1(_04326_),
    .B2(_04328_),
    .X(_04331_));
 sky130_fd_sc_hd__o2111a_2 _14810_ (.A1(_04327_),
    .A2(_04321_),
    .B1(_04320_),
    .C1(_03883_),
    .D1(_04326_),
    .X(_04332_));
 sky130_fd_sc_hd__o2111ai_4 _14811_ (.A1(_04327_),
    .A2(_04321_),
    .B1(_04320_),
    .C1(_03883_),
    .D1(_04326_),
    .Y(_04333_));
 sky130_fd_sc_hd__a22oi_1 _14812_ (.A1(net5),
    .A2(net37),
    .B1(net6),
    .B2(net36),
    .Y(_04334_));
 sky130_fd_sc_hd__a22o_2 _14813_ (.A1(net5),
    .A2(net37),
    .B1(net6),
    .B2(net36),
    .X(_04335_));
 sky130_fd_sc_hd__and4_1 _14814_ (.A(net36),
    .B(net5),
    .C(net37),
    .D(net6),
    .X(_04336_));
 sky130_fd_sc_hd__nand4_2 _14815_ (.A(net36),
    .B(net5),
    .C(net37),
    .D(net6),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_1 _14816_ (.A(net4),
    .B(net38),
    .Y(_04338_));
 sky130_fd_sc_hd__a22oi_2 _14817_ (.A1(net4),
    .A2(net38),
    .B1(_04335_),
    .B2(_04337_),
    .Y(_04339_));
 sky130_fd_sc_hd__and3_1 _14818_ (.A(_04337_),
    .B(net38),
    .C(net4),
    .X(_04341_));
 sky130_fd_sc_hd__a21oi_2 _14819_ (.A1(_04341_),
    .A2(_04335_),
    .B1(_04339_),
    .Y(_04342_));
 sky130_fd_sc_hd__a21o_2 _14820_ (.A1(_04341_),
    .A2(_04335_),
    .B1(_04339_),
    .X(_04343_));
 sky130_fd_sc_hd__o21ai_4 _14821_ (.A1(_04330_),
    .A2(_04332_),
    .B1(_04342_),
    .Y(_04344_));
 sky130_fd_sc_hd__nand3_4 _14822_ (.A(_04331_),
    .B(_04333_),
    .C(_04343_),
    .Y(_04345_));
 sky130_fd_sc_hd__o21ai_2 _14823_ (.A1(_04330_),
    .A2(_04332_),
    .B1(_04343_),
    .Y(_04346_));
 sky130_fd_sc_hd__nand3_1 _14824_ (.A(_04331_),
    .B(_04333_),
    .C(_04342_),
    .Y(_04347_));
 sky130_fd_sc_hd__o2bb2ai_2 _14825_ (.A1_N(_03919_),
    .A2_N(_03937_),
    .B1(_03933_),
    .B2(_03930_),
    .Y(_04348_));
 sky130_fd_sc_hd__a21boi_4 _14826_ (.A1(_03937_),
    .A2(_03919_),
    .B1_N(_03936_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand3_4 _14827_ (.A(_04344_),
    .B(_04345_),
    .C(_04349_),
    .Y(_04350_));
 sky130_fd_sc_hd__and3_1 _14828_ (.A(_04346_),
    .B(_04347_),
    .C(_04348_),
    .X(_04352_));
 sky130_fd_sc_hd__nand3_4 _14829_ (.A(_04346_),
    .B(_04347_),
    .C(_04348_),
    .Y(_04353_));
 sky130_fd_sc_hd__a21boi_4 _14830_ (.A1(_03890_),
    .A2(_03901_),
    .B1_N(_03892_),
    .Y(_04354_));
 sky130_fd_sc_hd__nand2_1 _14831_ (.A(_03892_),
    .B(_03906_),
    .Y(_04355_));
 sky130_fd_sc_hd__a21oi_4 _14832_ (.A1(_04350_),
    .A2(_04353_),
    .B1(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__a21o_1 _14833_ (.A1(_04350_),
    .A2(_04353_),
    .B1(_04355_),
    .X(_04357_));
 sky130_fd_sc_hd__a31o_1 _14834_ (.A1(_04344_),
    .A2(_04345_),
    .A3(_04349_),
    .B1(_04354_),
    .X(_04358_));
 sky130_fd_sc_hd__and3_2 _14835_ (.A(_04350_),
    .B(_04353_),
    .C(_04355_),
    .X(_04359_));
 sky130_fd_sc_hd__and3_1 _14836_ (.A(_04350_),
    .B(_04353_),
    .C(_04354_),
    .X(_04360_));
 sky130_fd_sc_hd__nand4_1 _14837_ (.A(_03892_),
    .B(_03906_),
    .C(_04350_),
    .D(_04353_),
    .Y(_04361_));
 sky130_fd_sc_hd__a21oi_1 _14838_ (.A1(_04350_),
    .A2(_04353_),
    .B1(_04354_),
    .Y(_04363_));
 sky130_fd_sc_hd__a22o_1 _14839_ (.A1(_03892_),
    .A2(_03906_),
    .B1(_04350_),
    .B2(_04353_),
    .X(_04364_));
 sky130_fd_sc_hd__o21ai_2 _14840_ (.A1(_04352_),
    .A2(_04358_),
    .B1(_04357_),
    .Y(_04365_));
 sky130_fd_sc_hd__a32oi_4 _14841_ (.A1(_03980_),
    .A2(_03981_),
    .A3(_03985_),
    .B1(_03943_),
    .B2(_03989_),
    .Y(_04366_));
 sky130_fd_sc_hd__a31o_1 _14842_ (.A1(_03938_),
    .A2(_03939_),
    .A3(_03989_),
    .B1(_03987_),
    .X(_04367_));
 sky130_fd_sc_hd__o21ai_1 _14843_ (.A1(_01780_),
    .A2(_02098_),
    .B1(_03952_),
    .Y(_04368_));
 sky130_fd_sc_hd__o21ai_4 _14844_ (.A1(_03947_),
    .A2(_03949_),
    .B1(_03952_),
    .Y(_04369_));
 sky130_fd_sc_hd__o21a_1 _14845_ (.A1(_03947_),
    .A2(_03949_),
    .B1(_03952_),
    .X(_04370_));
 sky130_fd_sc_hd__nand2_2 _14846_ (.A(net55),
    .B(net17),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_2 _14847_ (.A(net33),
    .B(net19),
    .Y(_04372_));
 sky130_fd_sc_hd__a22oi_4 _14848_ (.A1(net44),
    .A2(net18),
    .B1(net19),
    .B2(net33),
    .Y(_04374_));
 sky130_fd_sc_hd__a22o_2 _14849_ (.A1(net44),
    .A2(net18),
    .B1(net19),
    .B2(net33),
    .X(_04375_));
 sky130_fd_sc_hd__nand2_2 _14850_ (.A(net44),
    .B(net19),
    .Y(_04376_));
 sky130_fd_sc_hd__and4_1 _14851_ (.A(net33),
    .B(net44),
    .C(net18),
    .D(net19),
    .X(_04377_));
 sky130_fd_sc_hd__o211ai_2 _14852_ (.A1(_03948_),
    .A2(_04376_),
    .B1(_04375_),
    .C1(_04371_),
    .Y(_04378_));
 sky130_fd_sc_hd__o21bai_1 _14853_ (.A1(_04374_),
    .A2(_04377_),
    .B1_N(_04371_),
    .Y(_04379_));
 sky130_fd_sc_hd__o2bb2ai_4 _14854_ (.A1_N(net55),
    .A2_N(net17),
    .B1(_04374_),
    .B2(_04377_),
    .Y(_04380_));
 sky130_fd_sc_hd__o2111ai_4 _14855_ (.A1(_03948_),
    .A2(_04376_),
    .B1(net55),
    .C1(net17),
    .D1(_04375_),
    .Y(_04381_));
 sky130_fd_sc_hd__a22oi_1 _14856_ (.A1(_03950_),
    .A2(_04368_),
    .B1(_04380_),
    .B2(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand3_4 _14857_ (.A(_04370_),
    .B(_04378_),
    .C(_04379_),
    .Y(_04383_));
 sky130_fd_sc_hd__o31a_1 _14858_ (.A1(_04371_),
    .A2(_04374_),
    .A3(_04377_),
    .B1(_04369_),
    .X(_04385_));
 sky130_fd_sc_hd__nand3_4 _14859_ (.A(_04380_),
    .B(_04381_),
    .C(_04369_),
    .Y(_04386_));
 sky130_fd_sc_hd__nand2_1 _14860_ (.A(net60),
    .B(net14),
    .Y(_04387_));
 sky130_fd_sc_hd__a22oi_4 _14861_ (.A1(net59),
    .A2(net15),
    .B1(net16),
    .B2(net58),
    .Y(_04388_));
 sky130_fd_sc_hd__a22o_1 _14862_ (.A1(net59),
    .A2(net15),
    .B1(net16),
    .B2(net58),
    .X(_04389_));
 sky130_fd_sc_hd__and4_1 _14863_ (.A(net58),
    .B(net59),
    .C(net15),
    .D(net16),
    .X(_04390_));
 sky130_fd_sc_hd__nand4_2 _14864_ (.A(net58),
    .B(net59),
    .C(net15),
    .D(net16),
    .Y(_04391_));
 sky130_fd_sc_hd__and3_1 _14865_ (.A(_04387_),
    .B(_04389_),
    .C(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__o211ai_2 _14866_ (.A1(_01835_),
    .A2(_02065_),
    .B1(_04389_),
    .C1(_04391_),
    .Y(_04393_));
 sky130_fd_sc_hd__o211a_1 _14867_ (.A1(_04388_),
    .A2(_04390_),
    .B1(net60),
    .C1(net14),
    .X(_04394_));
 sky130_fd_sc_hd__o21bai_2 _14868_ (.A1(_04388_),
    .A2(_04390_),
    .B1_N(_04387_),
    .Y(_04396_));
 sky130_fd_sc_hd__o22a_1 _14869_ (.A1(_01835_),
    .A2(_02065_),
    .B1(_04388_),
    .B2(_04390_),
    .X(_04397_));
 sky130_fd_sc_hd__o21ai_2 _14870_ (.A1(_04388_),
    .A2(_04390_),
    .B1(_04387_),
    .Y(_04398_));
 sky130_fd_sc_hd__a41o_1 _14871_ (.A1(net58),
    .A2(net59),
    .A3(net15),
    .A4(net16),
    .B1(_04387_),
    .X(_04399_));
 sky130_fd_sc_hd__and4_1 _14872_ (.A(_04389_),
    .B(_04391_),
    .C(net60),
    .D(net14),
    .X(_04400_));
 sky130_fd_sc_hd__o21ai_1 _14873_ (.A1(_04388_),
    .A2(_04399_),
    .B1(_04398_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _14874_ (.A(_04393_),
    .B(_04396_),
    .Y(_04402_));
 sky130_fd_sc_hd__o2bb2ai_4 _14875_ (.A1_N(_04383_),
    .A2_N(_04386_),
    .B1(_04392_),
    .B2(_04394_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand4_4 _14876_ (.A(_04383_),
    .B(_04386_),
    .C(_04393_),
    .D(_04396_),
    .Y(_04404_));
 sky130_fd_sc_hd__o2bb2ai_1 _14877_ (.A1_N(_04383_),
    .A2_N(_04386_),
    .B1(_04397_),
    .B2(_04400_),
    .Y(_04405_));
 sky130_fd_sc_hd__o2111ai_4 _14878_ (.A1(_04388_),
    .A2(_04399_),
    .B1(_04398_),
    .C1(_04383_),
    .D1(_04386_),
    .Y(_04407_));
 sky130_fd_sc_hd__a2bb2oi_2 _14879_ (.A1_N(_03955_),
    .A2_N(_03961_),
    .B1(_03978_),
    .B2(_03960_),
    .Y(_04408_));
 sky130_fd_sc_hd__o22ai_2 _14880_ (.A1(_03955_),
    .A2(_03961_),
    .B1(_03977_),
    .B2(_03959_),
    .Y(_04409_));
 sky130_fd_sc_hd__a22oi_4 _14881_ (.A1(_03962_),
    .A2(_03983_),
    .B1(_04403_),
    .B2(_04404_),
    .Y(_04410_));
 sky130_fd_sc_hd__nand3_4 _14882_ (.A(_04405_),
    .B(_04407_),
    .C(_04409_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand3_4 _14883_ (.A(_04403_),
    .B(_04408_),
    .C(_04404_),
    .Y(_04412_));
 sky130_fd_sc_hd__o21ai_1 _14884_ (.A1(_03963_),
    .A2(_03964_),
    .B1(_03967_),
    .Y(_04413_));
 sky130_fd_sc_hd__o21a_1 _14885_ (.A1(_03963_),
    .A2(_03964_),
    .B1(_03967_),
    .X(_04414_));
 sky130_fd_sc_hd__nand2_1 _14886_ (.A(net62),
    .B(net13),
    .Y(_04415_));
 sky130_fd_sc_hd__nand4_4 _14887_ (.A(net61),
    .B(net62),
    .C(net11),
    .D(net13),
    .Y(_04416_));
 sky130_fd_sc_hd__nand2_1 _14888_ (.A(net61),
    .B(net13),
    .Y(_04418_));
 sky130_fd_sc_hd__a22oi_2 _14889_ (.A1(net62),
    .A2(net11),
    .B1(net13),
    .B2(net61),
    .Y(_04419_));
 sky130_fd_sc_hd__a22o_1 _14890_ (.A1(net62),
    .A2(net11),
    .B1(net13),
    .B2(net61),
    .X(_04420_));
 sky130_fd_sc_hd__o2bb2ai_1 _14891_ (.A1_N(_03922_),
    .A2_N(_04418_),
    .B1(_04415_),
    .B2(_03923_),
    .Y(_04421_));
 sky130_fd_sc_hd__o221ai_4 _14892_ (.A1(_01890_),
    .A2(_02021_),
    .B1(_03923_),
    .B2(_04415_),
    .C1(_04420_),
    .Y(_04422_));
 sky130_fd_sc_hd__nand3_2 _14893_ (.A(_04421_),
    .B(net10),
    .C(net63),
    .Y(_04423_));
 sky130_fd_sc_hd__a22o_1 _14894_ (.A1(net63),
    .A2(net10),
    .B1(_04416_),
    .B2(_04420_),
    .X(_04424_));
 sky130_fd_sc_hd__and4_1 _14895_ (.A(_04420_),
    .B(net10),
    .C(net63),
    .D(_04416_),
    .X(_04425_));
 sky130_fd_sc_hd__o2111ai_1 _14896_ (.A1(_03923_),
    .A2(_04415_),
    .B1(net63),
    .C1(net10),
    .D1(_04420_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand3_4 _14897_ (.A(_04414_),
    .B(_04422_),
    .C(_04423_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_1 _14898_ (.A(_04424_),
    .B(_04413_),
    .Y(_04429_));
 sky130_fd_sc_hd__a21oi_4 _14899_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04414_),
    .Y(_04430_));
 sky130_fd_sc_hd__nand3_2 _14900_ (.A(_04424_),
    .B(_04426_),
    .C(_04413_),
    .Y(_04431_));
 sky130_fd_sc_hd__o22a_1 _14901_ (.A1(_01890_),
    .A2(_01999_),
    .B1(_03697_),
    .B2(_03922_),
    .X(_04432_));
 sky130_fd_sc_hd__a2bb2o_2 _14902_ (.A1_N(_03697_),
    .A2_N(_03922_),
    .B1(_03921_),
    .B2(_03926_),
    .X(_04433_));
 sky130_fd_sc_hd__o2bb2a_1 _14903_ (.A1_N(_04427_),
    .A2_N(_04431_),
    .B1(_04432_),
    .B2(_03925_),
    .X(_04434_));
 sky130_fd_sc_hd__o2bb2ai_4 _14904_ (.A1_N(_04427_),
    .A2_N(_04431_),
    .B1(_04432_),
    .B2(_03925_),
    .Y(_04435_));
 sky130_fd_sc_hd__nand2_2 _14905_ (.A(_04427_),
    .B(_04433_),
    .Y(_04436_));
 sky130_fd_sc_hd__and3_1 _14906_ (.A(_04427_),
    .B(_04431_),
    .C(_04433_),
    .X(_04437_));
 sky130_fd_sc_hd__o211ai_2 _14907_ (.A1(_04425_),
    .A2(_04429_),
    .B1(_04433_),
    .C1(_04427_),
    .Y(_04438_));
 sky130_fd_sc_hd__o21ai_1 _14908_ (.A1(_04430_),
    .A2(_04436_),
    .B1(_04435_),
    .Y(_04440_));
 sky130_fd_sc_hd__o211ai_2 _14909_ (.A1(_04434_),
    .A2(_04437_),
    .B1(_04411_),
    .C1(_04412_),
    .Y(_04441_));
 sky130_fd_sc_hd__a21o_1 _14910_ (.A1(_04411_),
    .A2(_04412_),
    .B1(_04440_),
    .X(_04442_));
 sky130_fd_sc_hd__o2bb2ai_4 _14911_ (.A1_N(_04411_),
    .A2_N(_04412_),
    .B1(_04434_),
    .B2(_04437_),
    .Y(_04443_));
 sky130_fd_sc_hd__a31oi_2 _14912_ (.A1(_04403_),
    .A2(_04404_),
    .A3(_04408_),
    .B1(_04440_),
    .Y(_04444_));
 sky130_fd_sc_hd__o211ai_4 _14913_ (.A1(_04430_),
    .A2(_04436_),
    .B1(_04435_),
    .C1(_04412_),
    .Y(_04445_));
 sky130_fd_sc_hd__o2111ai_4 _14914_ (.A1(_04430_),
    .A2(_04436_),
    .B1(_04435_),
    .C1(_04411_),
    .D1(_04412_),
    .Y(_04446_));
 sky130_fd_sc_hd__o21ai_1 _14915_ (.A1(_04410_),
    .A2(_04445_),
    .B1(_04443_),
    .Y(_04447_));
 sky130_fd_sc_hd__a21oi_4 _14916_ (.A1(_04443_),
    .A2(_04446_),
    .B1(_04366_),
    .Y(_04448_));
 sky130_fd_sc_hd__o2111ai_4 _14917_ (.A1(_03943_),
    .A2(_03987_),
    .B1(_03989_),
    .C1(_04441_),
    .D1(_04442_),
    .Y(_04449_));
 sky130_fd_sc_hd__o211a_2 _14918_ (.A1(_04410_),
    .A2(_04445_),
    .B1(_04443_),
    .C1(_04366_),
    .X(_04451_));
 sky130_fd_sc_hd__o211ai_4 _14919_ (.A1(_04410_),
    .A2(_04445_),
    .B1(_04443_),
    .C1(_04366_),
    .Y(_04452_));
 sky130_fd_sc_hd__o211ai_4 _14920_ (.A1(_04356_),
    .A2(_04359_),
    .B1(_04449_),
    .C1(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__o22ai_4 _14921_ (.A1(_04360_),
    .A2(_04363_),
    .B1(_04448_),
    .B2(_04451_),
    .Y(_04454_));
 sky130_fd_sc_hd__o22ai_4 _14922_ (.A1(_04356_),
    .A2(_04359_),
    .B1(_04448_),
    .B2(_04451_),
    .Y(_04455_));
 sky130_fd_sc_hd__a22oi_2 _14923_ (.A1(_04361_),
    .A2(_04364_),
    .B1(_04447_),
    .B2(_04367_),
    .Y(_04456_));
 sky130_fd_sc_hd__o2111ai_4 _14924_ (.A1(_04358_),
    .A2(_04352_),
    .B1(_04357_),
    .C1(_04449_),
    .D1(_04452_),
    .Y(_04457_));
 sky130_fd_sc_hd__nand2_2 _14925_ (.A(_04455_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__a22oi_4 _14926_ (.A1(_03998_),
    .A2(_04317_),
    .B1(_04455_),
    .B2(_04457_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand3_2 _14927_ (.A(_04319_),
    .B(_04453_),
    .C(_04454_),
    .Y(_04460_));
 sky130_fd_sc_hd__a21oi_4 _14928_ (.A1(_04453_),
    .A2(_04454_),
    .B1(_04319_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand4_4 _14929_ (.A(_03998_),
    .B(_04317_),
    .C(_04455_),
    .D(_04457_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand4_4 _14930_ (.A(_04311_),
    .B(_04313_),
    .C(_04460_),
    .D(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__o22ai_4 _14931_ (.A1(_04310_),
    .A2(_04312_),
    .B1(_04459_),
    .B2(_04462_),
    .Y(_04465_));
 sky130_fd_sc_hd__a32oi_4 _14932_ (.A1(_04319_),
    .A2(_04453_),
    .A3(_04454_),
    .B1(_04313_),
    .B2(_04311_),
    .Y(_04466_));
 sky130_fd_sc_hd__o2bb2ai_4 _14933_ (.A1_N(_04319_),
    .A2_N(_04458_),
    .B1(_04310_),
    .B2(_04312_),
    .Y(_04467_));
 sky130_fd_sc_hd__o211ai_4 _14934_ (.A1(_04310_),
    .A2(_04312_),
    .B1(_04460_),
    .C1(_04463_),
    .Y(_04468_));
 sky130_fd_sc_hd__o22ai_4 _14935_ (.A1(_04314_),
    .A2(_04316_),
    .B1(_04459_),
    .B2(_04462_),
    .Y(_04469_));
 sky130_fd_sc_hd__a22oi_4 _14936_ (.A1(_04009_),
    .A2(_04097_),
    .B1(_04464_),
    .B2(_04465_),
    .Y(_04470_));
 sky130_fd_sc_hd__o211ai_4 _14937_ (.A1(_04462_),
    .A2(_04467_),
    .B1(_04469_),
    .C1(_04233_),
    .Y(_04471_));
 sky130_fd_sc_hd__a21oi_4 _14938_ (.A1(_04468_),
    .A2(_04469_),
    .B1(_04233_),
    .Y(_04473_));
 sky130_fd_sc_hd__nand3_2 _14939_ (.A(_04234_),
    .B(_04464_),
    .C(_04465_),
    .Y(_04474_));
 sky130_fd_sc_hd__o211ai_4 _14940_ (.A1(_04225_),
    .A2(_04229_),
    .B1(_04471_),
    .C1(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__a21o_1 _14941_ (.A1(_04471_),
    .A2(_04474_),
    .B1(_04232_),
    .X(_04476_));
 sky130_fd_sc_hd__o22ai_4 _14942_ (.A1(_04225_),
    .A2(_04229_),
    .B1(_04470_),
    .B2(_04473_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_2 _14943_ (.A(_04474_),
    .B(_04230_),
    .Y(_04478_));
 sky130_fd_sc_hd__o2111ai_1 _14944_ (.A1(_04228_),
    .A2(_04223_),
    .B1(_04226_),
    .C1(_04471_),
    .D1(_04474_),
    .Y(_04479_));
 sky130_fd_sc_hd__o211a_1 _14945_ (.A1(_04099_),
    .A2(_04177_),
    .B1(_04475_),
    .C1(_04476_),
    .X(_04480_));
 sky130_fd_sc_hd__o211ai_4 _14946_ (.A1(_04099_),
    .A2(_04177_),
    .B1(_04475_),
    .C1(_04476_),
    .Y(_04481_));
 sky130_fd_sc_hd__and3_1 _14947_ (.A(_04178_),
    .B(_04477_),
    .C(_04479_),
    .X(_04482_));
 sky130_fd_sc_hd__o211ai_4 _14948_ (.A1(_04478_),
    .A2(_04470_),
    .B1(_04178_),
    .C1(_04477_),
    .Y(_04484_));
 sky130_fd_sc_hd__o31a_1 _14949_ (.A1(_03063_),
    .A2(_03076_),
    .A3(_03600_),
    .B1(_04138_),
    .X(_04485_));
 sky130_fd_sc_hd__o311a_1 _14950_ (.A1(_03681_),
    .A2(_03688_),
    .A3(_04134_),
    .B1(_03601_),
    .C1(_03549_),
    .X(_04486_));
 sky130_fd_sc_hd__a31o_1 _14951_ (.A1(_03549_),
    .A2(_03601_),
    .A3(_04139_),
    .B1(_04137_),
    .X(_04487_));
 sky130_fd_sc_hd__o2bb2ai_1 _14952_ (.A1_N(_04481_),
    .A2_N(_04484_),
    .B1(_04486_),
    .B2(_04137_),
    .Y(_04488_));
 sky130_fd_sc_hd__a31oi_1 _14953_ (.A1(_04178_),
    .A2(_04477_),
    .A3(_04479_),
    .B1(_04487_),
    .Y(_04489_));
 sky130_fd_sc_hd__o21ai_4 _14954_ (.A1(_04140_),
    .A2(_04485_),
    .B1(_04484_),
    .Y(_04490_));
 sky130_fd_sc_hd__o2bb2ai_2 _14955_ (.A1_N(_04481_),
    .A2_N(_04484_),
    .B1(_04485_),
    .B2(_04140_),
    .Y(_04491_));
 sky130_fd_sc_hd__o21ai_1 _14956_ (.A1(_04137_),
    .A2(_04486_),
    .B1(_04481_),
    .Y(_04492_));
 sky130_fd_sc_hd__o211ai_2 _14957_ (.A1(_04137_),
    .A2(_04486_),
    .B1(_04484_),
    .C1(_04481_),
    .Y(_04493_));
 sky130_fd_sc_hd__o21ai_1 _14958_ (.A1(_04482_),
    .A2(_04492_),
    .B1(_04491_),
    .Y(_04495_));
 sky130_fd_sc_hd__a21oi_2 _14959_ (.A1(_03609_),
    .A2(_04153_),
    .B1(_04154_),
    .Y(_04496_));
 sky130_fd_sc_hd__o211ai_4 _14960_ (.A1(_04490_),
    .A2(_04480_),
    .B1(_04488_),
    .C1(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__o211a_1 _14961_ (.A1(_04154_),
    .A2(_04159_),
    .B1(_04491_),
    .C1(_04493_),
    .X(_04498_));
 sky130_fd_sc_hd__o211ai_4 _14962_ (.A1(_04154_),
    .A2(_04159_),
    .B1(_04491_),
    .C1(_04493_),
    .Y(_04499_));
 sky130_fd_sc_hd__o2bb2ai_2 _14963_ (.A1_N(_04497_),
    .A2_N(_04499_),
    .B1(_03872_),
    .B2(_04164_),
    .Y(_04500_));
 sky130_fd_sc_hd__o211ai_2 _14964_ (.A1(_04154_),
    .A2(_04160_),
    .B1(_04168_),
    .C1(_04497_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand4_2 _14965_ (.A(_04161_),
    .B(_04497_),
    .C(_04499_),
    .D(_04168_),
    .Y(_04502_));
 sky130_fd_sc_hd__o21ai_2 _14966_ (.A1(_04498_),
    .A2(_04501_),
    .B1(_04500_),
    .Y(_04503_));
 sky130_fd_sc_hd__and3_1 _14967_ (.A(_04173_),
    .B(_03861_),
    .C(_03858_),
    .X(_04504_));
 sky130_fd_sc_hd__o21ai_2 _14968_ (.A1(_03856_),
    .A2(_03860_),
    .B1(_04170_),
    .Y(_04506_));
 sky130_fd_sc_hd__a21boi_4 _14969_ (.A1(_03871_),
    .A2(_04504_),
    .B1_N(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__xor2_1 _14970_ (.A(_04503_),
    .B(_04507_),
    .X(net83));
 sky130_fd_sc_hd__a21o_1 _14971_ (.A1(_04481_),
    .A2(_04487_),
    .B1(_04482_),
    .X(_04508_));
 sky130_fd_sc_hd__a21oi_1 _14972_ (.A1(_04481_),
    .A2(_04487_),
    .B1(_04482_),
    .Y(_04509_));
 sky130_fd_sc_hd__a21oi_1 _14973_ (.A1(_04131_),
    .A2(_04224_),
    .B1(_04221_),
    .Y(_04510_));
 sky130_fd_sc_hd__a31o_1 _14974_ (.A1(_03599_),
    .A2(_04126_),
    .A3(_04224_),
    .B1(_04221_),
    .X(_04511_));
 sky130_fd_sc_hd__a31oi_2 _14975_ (.A1(_04233_),
    .A2(_04468_),
    .A3(_04469_),
    .B1(_04230_),
    .Y(_04512_));
 sky130_fd_sc_hd__a32oi_4 _14976_ (.A1(_04234_),
    .A2(_04464_),
    .A3(_04465_),
    .B1(_04471_),
    .B2(_04232_),
    .Y(_04513_));
 sky130_fd_sc_hd__a21oi_1 _14977_ (.A1(_04289_),
    .A2(_04268_),
    .B1(_04286_),
    .Y(_04514_));
 sky130_fd_sc_hd__o21a_1 _14978_ (.A1(_01912_),
    .A2(_02010_),
    .B1(_04279_),
    .X(_04516_));
 sky130_fd_sc_hd__and3_1 _14979_ (.A(_04276_),
    .B(net41),
    .C(net32),
    .X(_04517_));
 sky130_fd_sc_hd__o31a_1 _14980_ (.A1(_01912_),
    .A2(_02010_),
    .A3(_04275_),
    .B1(_04279_),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _14981_ (.A(_04337_),
    .B(_04338_),
    .Y(_04519_));
 sky130_fd_sc_hd__nor2_1 _14982_ (.A(_04338_),
    .B(_04334_),
    .Y(_04520_));
 sky130_fd_sc_hd__o21ai_1 _14983_ (.A1(_04338_),
    .A2(_04334_),
    .B1(_04337_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand2_2 _14984_ (.A(net4),
    .B(net40),
    .Y(_04522_));
 sky130_fd_sc_hd__and4_1 _14985_ (.A(net3),
    .B(net4),
    .C(net39),
    .D(net40),
    .X(_04523_));
 sky130_fd_sc_hd__nand2_1 _14986_ (.A(net4),
    .B(net39),
    .Y(_04524_));
 sky130_fd_sc_hd__a22o_1 _14987_ (.A1(net4),
    .A2(net39),
    .B1(net40),
    .B2(net3),
    .X(_04525_));
 sky130_fd_sc_hd__o2bb2ai_1 _14988_ (.A1_N(_04277_),
    .A2_N(_04524_),
    .B1(_04522_),
    .B2(_04273_),
    .Y(_04527_));
 sky130_fd_sc_hd__o221ai_2 _14989_ (.A1(_01901_),
    .A2(_02010_),
    .B1(_04273_),
    .B2(_04522_),
    .C1(_04525_),
    .Y(_04528_));
 sky130_fd_sc_hd__nand3_1 _14990_ (.A(_04527_),
    .B(net41),
    .C(net2),
    .Y(_04529_));
 sky130_fd_sc_hd__o2111ai_4 _14991_ (.A1(_04273_),
    .A2(_04522_),
    .B1(net2),
    .C1(net41),
    .D1(_04525_),
    .Y(_04530_));
 sky130_fd_sc_hd__o21ai_2 _14992_ (.A1(_01901_),
    .A2(_02010_),
    .B1(_04527_),
    .Y(_04531_));
 sky130_fd_sc_hd__a2bb2oi_1 _14993_ (.A1_N(_04336_),
    .A2_N(_04520_),
    .B1(_04528_),
    .B2(_04529_),
    .Y(_04532_));
 sky130_fd_sc_hd__o211ai_4 _14994_ (.A1(_04336_),
    .A2(_04520_),
    .B1(_04530_),
    .C1(_04531_),
    .Y(_04533_));
 sky130_fd_sc_hd__a22oi_4 _14995_ (.A1(_04335_),
    .A2(_04519_),
    .B1(_04530_),
    .B2(_04531_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand3b_1 _14996_ (.A_N(_04521_),
    .B(_04528_),
    .C(_04529_),
    .Y(_04535_));
 sky130_fd_sc_hd__o211ai_2 _14997_ (.A1(_04278_),
    .A2(_04517_),
    .B1(_04533_),
    .C1(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__o22ai_2 _14998_ (.A1(_04275_),
    .A2(_04516_),
    .B1(_04532_),
    .B2(_04534_),
    .Y(_04538_));
 sky130_fd_sc_hd__o22ai_1 _14999_ (.A1(_04278_),
    .A2(_04517_),
    .B1(_04532_),
    .B2(_04534_),
    .Y(_04539_));
 sky130_fd_sc_hd__o2111ai_2 _15000_ (.A1(_04272_),
    .A2(_04275_),
    .B1(_04279_),
    .C1(_04533_),
    .D1(_04535_),
    .Y(_04540_));
 sky130_fd_sc_hd__and3_2 _15001_ (.A(_04539_),
    .B(_04540_),
    .C(_04514_),
    .X(_04541_));
 sky130_fd_sc_hd__nand3_2 _15002_ (.A(_04539_),
    .B(_04540_),
    .C(_04514_),
    .Y(_04542_));
 sky130_fd_sc_hd__o211ai_4 _15003_ (.A1(_04286_),
    .A2(_04290_),
    .B1(_04536_),
    .C1(_04538_),
    .Y(_04543_));
 sky130_fd_sc_hd__o21ai_2 _15004_ (.A1(_04237_),
    .A2(_04240_),
    .B1(_04239_),
    .Y(_04544_));
 sky130_fd_sc_hd__a22oi_4 _15005_ (.A1(net32),
    .A2(net42),
    .B1(net43),
    .B2(net31),
    .Y(_04545_));
 sky130_fd_sc_hd__a22o_1 _15006_ (.A1(net32),
    .A2(net42),
    .B1(net43),
    .B2(net31),
    .X(_04546_));
 sky130_fd_sc_hd__and4_1 _15007_ (.A(net31),
    .B(net32),
    .C(net42),
    .D(net43),
    .X(_04547_));
 sky130_fd_sc_hd__nand4_2 _15008_ (.A(net31),
    .B(net32),
    .C(net42),
    .D(net43),
    .Y(_04549_));
 sky130_fd_sc_hd__o22ai_4 _15009_ (.A1(_01868_),
    .A2(_02054_),
    .B1(_04545_),
    .B2(_04547_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand4_4 _15010_ (.A(_04546_),
    .B(_04549_),
    .C(net30),
    .D(net45),
    .Y(_04551_));
 sky130_fd_sc_hd__a21oi_2 _15011_ (.A1(_04550_),
    .A2(_04551_),
    .B1(_04544_),
    .Y(_04552_));
 sky130_fd_sc_hd__a21o_2 _15012_ (.A1(_04550_),
    .A2(_04551_),
    .B1(_04544_),
    .X(_04553_));
 sky130_fd_sc_hd__nand3_4 _15013_ (.A(_04550_),
    .B(_04551_),
    .C(_04544_),
    .Y(_04554_));
 sky130_fd_sc_hd__nand2_1 _15014_ (.A(net27),
    .B(net48),
    .Y(_04555_));
 sky130_fd_sc_hd__a22oi_4 _15015_ (.A1(net29),
    .A2(net46),
    .B1(net47),
    .B2(net28),
    .Y(_04556_));
 sky130_fd_sc_hd__nand2_1 _15016_ (.A(net29),
    .B(net47),
    .Y(_04557_));
 sky130_fd_sc_hd__and4_1 _15017_ (.A(net28),
    .B(net29),
    .C(net46),
    .D(net47),
    .X(_04558_));
 sky130_fd_sc_hd__a211o_2 _15018_ (.A1(net27),
    .A2(net48),
    .B1(_04556_),
    .C1(_04558_),
    .X(_04560_));
 sky130_fd_sc_hd__o211ai_4 _15019_ (.A1(_04556_),
    .A2(_04558_),
    .B1(net27),
    .C1(net48),
    .Y(_04561_));
 sky130_fd_sc_hd__nand2_1 _15020_ (.A(_04560_),
    .B(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__and3_1 _15021_ (.A(_04553_),
    .B(_04554_),
    .C(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__a21oi_1 _15022_ (.A1(_04553_),
    .A2(_04554_),
    .B1(_04562_),
    .Y(_04564_));
 sky130_fd_sc_hd__and4_1 _15023_ (.A(_04553_),
    .B(_04554_),
    .C(_04560_),
    .D(_04561_),
    .X(_04565_));
 sky130_fd_sc_hd__nand4_4 _15024_ (.A(_04553_),
    .B(_04554_),
    .C(_04560_),
    .D(_04561_),
    .Y(_04566_));
 sky130_fd_sc_hd__a22oi_2 _15025_ (.A1(_04553_),
    .A2(_04554_),
    .B1(_04560_),
    .B2(_04561_),
    .Y(_04567_));
 sky130_fd_sc_hd__a22o_1 _15026_ (.A1(_04553_),
    .A2(_04554_),
    .B1(_04560_),
    .B2(_04561_),
    .X(_04568_));
 sky130_fd_sc_hd__o2bb2ai_1 _15027_ (.A1_N(_04542_),
    .A2_N(_04543_),
    .B1(_04565_),
    .B2(_04567_),
    .Y(_04569_));
 sky130_fd_sc_hd__nand3_2 _15028_ (.A(_04543_),
    .B(_04566_),
    .C(_04568_),
    .Y(_04571_));
 sky130_fd_sc_hd__o2bb2ai_1 _15029_ (.A1_N(_04542_),
    .A2_N(_04543_),
    .B1(_04563_),
    .B2(_04564_),
    .Y(_04572_));
 sky130_fd_sc_hd__o211ai_2 _15030_ (.A1(_04565_),
    .A2(_04567_),
    .B1(_04542_),
    .C1(_04543_),
    .Y(_04573_));
 sky130_fd_sc_hd__a32oi_4 _15031_ (.A1(_04344_),
    .A2(_04345_),
    .A3(_04349_),
    .B1(_04353_),
    .B2(_04354_),
    .Y(_04574_));
 sky130_fd_sc_hd__a32o_1 _15032_ (.A1(_04344_),
    .A2(_04345_),
    .A3(_04349_),
    .B1(_04353_),
    .B2(_04354_),
    .X(_04575_));
 sky130_fd_sc_hd__a21oi_1 _15033_ (.A1(_04572_),
    .A2(_04573_),
    .B1(_04574_),
    .Y(_04576_));
 sky130_fd_sc_hd__o211ai_4 _15034_ (.A1(_04571_),
    .A2(_04541_),
    .B1(_04569_),
    .C1(_04575_),
    .Y(_04577_));
 sky130_fd_sc_hd__and3_2 _15035_ (.A(_04572_),
    .B(_04574_),
    .C(_04573_),
    .X(_04578_));
 sky130_fd_sc_hd__nand3_1 _15036_ (.A(_04572_),
    .B(_04574_),
    .C(_04573_),
    .Y(_04579_));
 sky130_fd_sc_hd__o31a_1 _15037_ (.A1(_04260_),
    .A2(_04261_),
    .A3(_04298_),
    .B1(_04297_),
    .X(_04580_));
 sky130_fd_sc_hd__a21o_1 _15038_ (.A1(_04299_),
    .A2(_04265_),
    .B1(_04295_),
    .X(_04582_));
 sky130_fd_sc_hd__a21o_2 _15039_ (.A1(_04577_),
    .A2(_04579_),
    .B1(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__nand2_2 _15040_ (.A(_04577_),
    .B(_04582_),
    .Y(_04584_));
 sky130_fd_sc_hd__o211ai_1 _15041_ (.A1(_04295_),
    .A2(_04301_),
    .B1(_04577_),
    .C1(_04579_),
    .Y(_04585_));
 sky130_fd_sc_hd__o21ai_4 _15042_ (.A1(_04578_),
    .A2(_04584_),
    .B1(_04583_),
    .Y(_04586_));
 sky130_fd_sc_hd__o31a_1 _15043_ (.A1(_04356_),
    .A2(_04359_),
    .A3(_04448_),
    .B1(_04452_),
    .X(_04587_));
 sky130_fd_sc_hd__a31oi_2 _15044_ (.A1(_04412_),
    .A2(_04435_),
    .A3(_04438_),
    .B1(_04410_),
    .Y(_04588_));
 sky130_fd_sc_hd__a31o_1 _15045_ (.A1(_04412_),
    .A2(_04435_),
    .A3(_04438_),
    .B1(_04410_),
    .X(_04589_));
 sky130_fd_sc_hd__o21ai_1 _15046_ (.A1(_04387_),
    .A2(_04388_),
    .B1(_04391_),
    .Y(_04590_));
 sky130_fd_sc_hd__o31a_1 _15047_ (.A1(_01835_),
    .A2(_02065_),
    .A3(_04388_),
    .B1(_04391_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_1 _15048_ (.A(net63),
    .B(net11),
    .Y(_04593_));
 sky130_fd_sc_hd__a22oi_4 _15049_ (.A1(net62),
    .A2(net13),
    .B1(net14),
    .B2(net61),
    .Y(_04594_));
 sky130_fd_sc_hd__a22o_1 _15050_ (.A1(net62),
    .A2(net13),
    .B1(net14),
    .B2(net61),
    .X(_04595_));
 sky130_fd_sc_hd__and4_1 _15051_ (.A(net61),
    .B(net62),
    .C(net13),
    .D(net14),
    .X(_04596_));
 sky130_fd_sc_hd__nand4_2 _15052_ (.A(net61),
    .B(net62),
    .C(net13),
    .D(net14),
    .Y(_04597_));
 sky130_fd_sc_hd__o211ai_4 _15053_ (.A1(_01890_),
    .A2(_02032_),
    .B1(_04595_),
    .C1(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__o21bai_2 _15054_ (.A1(_04594_),
    .A2(_04596_),
    .B1_N(_04593_),
    .Y(_04599_));
 sky130_fd_sc_hd__o21ai_1 _15055_ (.A1(_04594_),
    .A2(_04596_),
    .B1(_04593_),
    .Y(_04600_));
 sky130_fd_sc_hd__nand4_1 _15056_ (.A(_04595_),
    .B(_04597_),
    .C(net63),
    .D(net11),
    .Y(_04601_));
 sky130_fd_sc_hd__nand3_1 _15057_ (.A(_04591_),
    .B(_04598_),
    .C(_04599_),
    .Y(_04602_));
 sky130_fd_sc_hd__and3_4 _15058_ (.A(_04600_),
    .B(_04601_),
    .C(_04590_),
    .X(_04604_));
 sky130_fd_sc_hd__nand3_1 _15059_ (.A(_04600_),
    .B(_04601_),
    .C(_04590_),
    .Y(_04605_));
 sky130_fd_sc_hd__or3_1 _15060_ (.A(_01890_),
    .B(_02021_),
    .C(_04419_),
    .X(_04606_));
 sky130_fd_sc_hd__o31ai_2 _15061_ (.A1(_01890_),
    .A2(_02021_),
    .A3(_04419_),
    .B1(_04416_),
    .Y(_04607_));
 sky130_fd_sc_hd__a21o_2 _15062_ (.A1(_04602_),
    .A2(_04605_),
    .B1(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__a32oi_4 _15063_ (.A1(_04591_),
    .A2(_04598_),
    .A3(_04599_),
    .B1(_04606_),
    .B2(_04416_),
    .Y(_04609_));
 sky130_fd_sc_hd__a32o_2 _15064_ (.A1(_04591_),
    .A2(_04598_),
    .A3(_04599_),
    .B1(_04606_),
    .B2(_04416_),
    .X(_04610_));
 sky130_fd_sc_hd__nand2_1 _15065_ (.A(_04609_),
    .B(_04605_),
    .Y(_04611_));
 sky130_fd_sc_hd__o21ai_4 _15066_ (.A1(_04604_),
    .A2(_04610_),
    .B1(_04608_),
    .Y(_04612_));
 sky130_fd_sc_hd__o21ai_1 _15067_ (.A1(_03948_),
    .A2(_04376_),
    .B1(_04371_),
    .Y(_04613_));
 sky130_fd_sc_hd__o22ai_4 _15068_ (.A1(_03948_),
    .A2(_04376_),
    .B1(_04371_),
    .B2(_04374_),
    .Y(_04615_));
 sky130_fd_sc_hd__o22a_1 _15069_ (.A1(_03948_),
    .A2(_04376_),
    .B1(_04371_),
    .B2(_04374_),
    .X(_04616_));
 sky130_fd_sc_hd__and2_1 _15070_ (.A(net55),
    .B(net18),
    .X(_04617_));
 sky130_fd_sc_hd__nand2_2 _15071_ (.A(net55),
    .B(net18),
    .Y(_04618_));
 sky130_fd_sc_hd__a22oi_4 _15072_ (.A1(net44),
    .A2(net19),
    .B1(net20),
    .B2(net33),
    .Y(_04619_));
 sky130_fd_sc_hd__a22o_2 _15073_ (.A1(net44),
    .A2(net19),
    .B1(net20),
    .B2(net33),
    .X(_04620_));
 sky130_fd_sc_hd__nand2_2 _15074_ (.A(net44),
    .B(net20),
    .Y(_04621_));
 sky130_fd_sc_hd__and4_1 _15075_ (.A(net33),
    .B(net44),
    .C(net19),
    .D(net20),
    .X(_04622_));
 sky130_fd_sc_hd__nand4_2 _15076_ (.A(net33),
    .B(net44),
    .C(net19),
    .D(net20),
    .Y(_04623_));
 sky130_fd_sc_hd__o221ai_4 _15077_ (.A1(_01780_),
    .A2(_02131_),
    .B1(_04372_),
    .B2(_04621_),
    .C1(_04620_),
    .Y(_04624_));
 sky130_fd_sc_hd__o21bai_1 _15078_ (.A1(_04619_),
    .A2(_04622_),
    .B1_N(_04618_),
    .Y(_04626_));
 sky130_fd_sc_hd__o22a_2 _15079_ (.A1(_01780_),
    .A2(_02131_),
    .B1(_04619_),
    .B2(_04622_),
    .X(_04627_));
 sky130_fd_sc_hd__o21ai_4 _15080_ (.A1(_04619_),
    .A2(_04622_),
    .B1(_04618_),
    .Y(_04628_));
 sky130_fd_sc_hd__nand3_4 _15081_ (.A(_04620_),
    .B(_04623_),
    .C(_04617_),
    .Y(_04629_));
 sky130_fd_sc_hd__a22oi_4 _15082_ (.A1(_04375_),
    .A2(_04613_),
    .B1(_04628_),
    .B2(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__nand3_4 _15083_ (.A(_04616_),
    .B(_04624_),
    .C(_04626_),
    .Y(_04631_));
 sky130_fd_sc_hd__nand2_2 _15084_ (.A(_04615_),
    .B(_04629_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand3_2 _15085_ (.A(_04628_),
    .B(_04629_),
    .C(_04615_),
    .Y(_04633_));
 sky130_fd_sc_hd__nand2_1 _15086_ (.A(net60),
    .B(net15),
    .Y(_04634_));
 sky130_fd_sc_hd__a22oi_4 _15087_ (.A1(net59),
    .A2(net16),
    .B1(net17),
    .B2(net58),
    .Y(_04635_));
 sky130_fd_sc_hd__a22o_1 _15088_ (.A1(net59),
    .A2(net16),
    .B1(net17),
    .B2(net58),
    .X(_04637_));
 sky130_fd_sc_hd__and4_1 _15089_ (.A(net58),
    .B(net59),
    .C(net16),
    .D(net17),
    .X(_04638_));
 sky130_fd_sc_hd__nand4_4 _15090_ (.A(net58),
    .B(net59),
    .C(net16),
    .D(net17),
    .Y(_04639_));
 sky130_fd_sc_hd__and3_1 _15091_ (.A(_04634_),
    .B(_04637_),
    .C(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__o211ai_2 _15092_ (.A1(_01835_),
    .A2(_02076_),
    .B1(_04637_),
    .C1(_04639_),
    .Y(_04641_));
 sky130_fd_sc_hd__o211a_1 _15093_ (.A1(_04635_),
    .A2(_04638_),
    .B1(net60),
    .C1(net15),
    .X(_04642_));
 sky130_fd_sc_hd__a21o_1 _15094_ (.A1(_04637_),
    .A2(_04639_),
    .B1(_04634_),
    .X(_04643_));
 sky130_fd_sc_hd__o22a_1 _15095_ (.A1(_01835_),
    .A2(_02076_),
    .B1(_04635_),
    .B2(_04638_),
    .X(_04644_));
 sky130_fd_sc_hd__o21ai_1 _15096_ (.A1(_04635_),
    .A2(_04638_),
    .B1(_04634_),
    .Y(_04645_));
 sky130_fd_sc_hd__a41o_1 _15097_ (.A1(net58),
    .A2(net59),
    .A3(net16),
    .A4(net17),
    .B1(_04634_),
    .X(_04646_));
 sky130_fd_sc_hd__and4_1 _15098_ (.A(_04637_),
    .B(_04639_),
    .C(net60),
    .D(net15),
    .X(_04648_));
 sky130_fd_sc_hd__o21ai_1 _15099_ (.A1(_04635_),
    .A2(_04646_),
    .B1(_04645_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_1 _15100_ (.A(_04641_),
    .B(_04643_),
    .Y(_04650_));
 sky130_fd_sc_hd__o2bb2ai_2 _15101_ (.A1_N(_04641_),
    .A2_N(_04643_),
    .B1(_04627_),
    .B2(_04632_),
    .Y(_04651_));
 sky130_fd_sc_hd__o2bb2ai_2 _15102_ (.A1_N(_04631_),
    .A2_N(_04633_),
    .B1(_04644_),
    .B2(_04648_),
    .Y(_04652_));
 sky130_fd_sc_hd__o221ai_4 _15103_ (.A1(_04644_),
    .A2(_04648_),
    .B1(_04627_),
    .B2(_04632_),
    .C1(_04631_),
    .Y(_04653_));
 sky130_fd_sc_hd__o2bb2ai_4 _15104_ (.A1_N(_04631_),
    .A2_N(_04633_),
    .B1(_04640_),
    .B2(_04642_),
    .Y(_04654_));
 sky130_fd_sc_hd__a32oi_4 _15105_ (.A1(_04369_),
    .A2(_04380_),
    .A3(_04381_),
    .B1(_04383_),
    .B2(_04402_),
    .Y(_04655_));
 sky130_fd_sc_hd__o2bb2ai_2 _15106_ (.A1_N(_04380_),
    .A2_N(_04385_),
    .B1(_04401_),
    .B2(_04382_),
    .Y(_04656_));
 sky130_fd_sc_hd__and3_1 _15107_ (.A(_04655_),
    .B(_04654_),
    .C(_04653_),
    .X(_04657_));
 sky130_fd_sc_hd__nand3_2 _15108_ (.A(_04653_),
    .B(_04654_),
    .C(_04655_),
    .Y(_04659_));
 sky130_fd_sc_hd__o211a_1 _15109_ (.A1(_04651_),
    .A2(_04630_),
    .B1(_04656_),
    .C1(_04652_),
    .X(_04660_));
 sky130_fd_sc_hd__o211ai_4 _15110_ (.A1(_04651_),
    .A2(_04630_),
    .B1(_04656_),
    .C1(_04652_),
    .Y(_04661_));
 sky130_fd_sc_hd__nand3_1 _15111_ (.A(_04612_),
    .B(_04659_),
    .C(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__a21o_1 _15112_ (.A1(_04659_),
    .A2(_04661_),
    .B1(_04612_),
    .X(_04663_));
 sky130_fd_sc_hd__a22o_2 _15113_ (.A1(_04608_),
    .A2(_04611_),
    .B1(_04659_),
    .B2(_04661_),
    .X(_04664_));
 sky130_fd_sc_hd__o211ai_2 _15114_ (.A1(_04610_),
    .A2(_04604_),
    .B1(_04608_),
    .C1(_04659_),
    .Y(_04665_));
 sky130_fd_sc_hd__o2111ai_4 _15115_ (.A1(_04610_),
    .A2(_04604_),
    .B1(_04608_),
    .C1(_04659_),
    .D1(_04661_),
    .Y(_04666_));
 sky130_fd_sc_hd__and3_1 _15116_ (.A(_04663_),
    .B(_04588_),
    .C(_04662_),
    .X(_04667_));
 sky130_fd_sc_hd__nand3_4 _15117_ (.A(_04663_),
    .B(_04588_),
    .C(_04662_),
    .Y(_04668_));
 sky130_fd_sc_hd__o221ai_4 _15118_ (.A1(_04660_),
    .A2(_04665_),
    .B1(_04410_),
    .B2(_04444_),
    .C1(_04664_),
    .Y(_04670_));
 sky130_fd_sc_hd__o21ai_2 _15119_ (.A1(_01934_),
    .A2(_01977_),
    .B1(_04324_),
    .Y(_04671_));
 sky130_fd_sc_hd__nor2_1 _15120_ (.A(_04325_),
    .B(_04321_),
    .Y(_04672_));
 sky130_fd_sc_hd__nand2_1 _15121_ (.A(net64),
    .B(net10),
    .Y(_04673_));
 sky130_fd_sc_hd__a22oi_4 _15122_ (.A1(net34),
    .A2(net9),
    .B1(net10),
    .B2(net64),
    .Y(_04674_));
 sky130_fd_sc_hd__a22o_1 _15123_ (.A1(net34),
    .A2(net9),
    .B1(net10),
    .B2(net64),
    .X(_04675_));
 sky130_fd_sc_hd__and4_1 _15124_ (.A(net64),
    .B(net34),
    .C(net9),
    .D(net10),
    .X(_04676_));
 sky130_fd_sc_hd__nand4_2 _15125_ (.A(net64),
    .B(net34),
    .C(net9),
    .D(net10),
    .Y(_04677_));
 sky130_fd_sc_hd__o22ai_4 _15126_ (.A1(_01934_),
    .A2(_01988_),
    .B1(_04674_),
    .B2(_04676_),
    .Y(_04678_));
 sky130_fd_sc_hd__nand4_4 _15127_ (.A(_04675_),
    .B(_04677_),
    .C(net35),
    .D(net8),
    .Y(_04679_));
 sky130_fd_sc_hd__a22oi_4 _15128_ (.A1(_04322_),
    .A2(_04671_),
    .B1(_04678_),
    .B2(_04679_),
    .Y(_04681_));
 sky130_fd_sc_hd__a22o_1 _15129_ (.A1(_04322_),
    .A2(_04671_),
    .B1(_04678_),
    .B2(_04679_),
    .X(_04682_));
 sky130_fd_sc_hd__o211a_1 _15130_ (.A1(_04323_),
    .A2(_04672_),
    .B1(_04678_),
    .C1(_04679_),
    .X(_04683_));
 sky130_fd_sc_hd__o211ai_4 _15131_ (.A1(_04323_),
    .A2(_04672_),
    .B1(_04678_),
    .C1(_04679_),
    .Y(_04684_));
 sky130_fd_sc_hd__a22oi_4 _15132_ (.A1(net37),
    .A2(net6),
    .B1(net7),
    .B2(net36),
    .Y(_04685_));
 sky130_fd_sc_hd__a22o_1 _15133_ (.A1(net37),
    .A2(net6),
    .B1(net7),
    .B2(net36),
    .X(_04686_));
 sky130_fd_sc_hd__nand4_1 _15134_ (.A(net36),
    .B(net37),
    .C(net6),
    .D(net7),
    .Y(_04687_));
 sky130_fd_sc_hd__nand2_1 _15135_ (.A(net5),
    .B(net38),
    .Y(_04688_));
 sky130_fd_sc_hd__a22o_1 _15136_ (.A1(net5),
    .A2(net38),
    .B1(_04686_),
    .B2(_04687_),
    .X(_04689_));
 sky130_fd_sc_hd__a41o_1 _15137_ (.A1(net36),
    .A2(net37),
    .A3(net6),
    .A4(net7),
    .B1(_04688_),
    .X(_04690_));
 sky130_fd_sc_hd__o21a_1 _15138_ (.A1(_04685_),
    .A2(_04690_),
    .B1(_04689_),
    .X(_04692_));
 sky130_fd_sc_hd__o21ai_4 _15139_ (.A1(_04685_),
    .A2(_04690_),
    .B1(_04689_),
    .Y(_04693_));
 sky130_fd_sc_hd__o21ai_4 _15140_ (.A1(_04681_),
    .A2(_04683_),
    .B1(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__nand3_2 _15141_ (.A(_04682_),
    .B(_04684_),
    .C(_04693_),
    .Y(_04695_));
 sky130_fd_sc_hd__o21ai_1 _15142_ (.A1(_04681_),
    .A2(_04683_),
    .B1(_04693_),
    .Y(_04696_));
 sky130_fd_sc_hd__nand2_1 _15143_ (.A(_04692_),
    .B(_04682_),
    .Y(_04697_));
 sky130_fd_sc_hd__nand3_1 _15144_ (.A(_04682_),
    .B(_04692_),
    .C(_04684_),
    .Y(_04698_));
 sky130_fd_sc_hd__a21oi_4 _15145_ (.A1(_04427_),
    .A2(_04433_),
    .B1(_04430_),
    .Y(_04699_));
 sky130_fd_sc_hd__o2bb2ai_2 _15146_ (.A1_N(_04433_),
    .A2_N(_04427_),
    .B1(_04425_),
    .B2(_04429_),
    .Y(_04700_));
 sky130_fd_sc_hd__nand3_4 _15147_ (.A(_04694_),
    .B(_04699_),
    .C(_04695_),
    .Y(_04701_));
 sky130_fd_sc_hd__a21oi_1 _15148_ (.A1(_04694_),
    .A2(_04695_),
    .B1(_04699_),
    .Y(_04703_));
 sky130_fd_sc_hd__nand3_4 _15149_ (.A(_04696_),
    .B(_04698_),
    .C(_04700_),
    .Y(_04704_));
 sky130_fd_sc_hd__a21oi_2 _15150_ (.A1(_04331_),
    .A2(_04342_),
    .B1(_04332_),
    .Y(_04705_));
 sky130_fd_sc_hd__o21ai_2 _15151_ (.A1(_04330_),
    .A2(_04343_),
    .B1(_04333_),
    .Y(_04706_));
 sky130_fd_sc_hd__a21oi_2 _15152_ (.A1(_04701_),
    .A2(_04704_),
    .B1(_04705_),
    .Y(_04707_));
 sky130_fd_sc_hd__a21o_1 _15153_ (.A1(_04701_),
    .A2(_04704_),
    .B1(_04705_),
    .X(_04708_));
 sky130_fd_sc_hd__and3_1 _15154_ (.A(_04701_),
    .B(_04704_),
    .C(_04705_),
    .X(_04709_));
 sky130_fd_sc_hd__o2111ai_4 _15155_ (.A1(_04343_),
    .A2(_04330_),
    .B1(_04333_),
    .C1(_04701_),
    .D1(_04704_),
    .Y(_04710_));
 sky130_fd_sc_hd__a21oi_1 _15156_ (.A1(_04701_),
    .A2(_04704_),
    .B1(_04706_),
    .Y(_04711_));
 sky130_fd_sc_hd__a21o_1 _15157_ (.A1(_04701_),
    .A2(_04704_),
    .B1(_04706_),
    .X(_04712_));
 sky130_fd_sc_hd__and3_1 _15158_ (.A(_04701_),
    .B(_04704_),
    .C(_04706_),
    .X(_04714_));
 sky130_fd_sc_hd__nand3_1 _15159_ (.A(_04701_),
    .B(_04704_),
    .C(_04706_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand2_1 _15160_ (.A(_04708_),
    .B(_04710_),
    .Y(_04716_));
 sky130_fd_sc_hd__o211ai_2 _15161_ (.A1(_04707_),
    .A2(_04709_),
    .B1(_04668_),
    .C1(_04670_),
    .Y(_04717_));
 sky130_fd_sc_hd__o2bb2ai_1 _15162_ (.A1_N(_04668_),
    .A2_N(_04670_),
    .B1(_04711_),
    .B2(_04714_),
    .Y(_04718_));
 sky130_fd_sc_hd__nand4_4 _15163_ (.A(_04668_),
    .B(_04670_),
    .C(_04708_),
    .D(_04710_),
    .Y(_04719_));
 sky130_fd_sc_hd__o2bb2ai_4 _15164_ (.A1_N(_04668_),
    .A2_N(_04670_),
    .B1(_04707_),
    .B2(_04709_),
    .Y(_04720_));
 sky130_fd_sc_hd__o2111a_2 _15165_ (.A1(_04365_),
    .A2(_04448_),
    .B1(_04452_),
    .C1(_04719_),
    .D1(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__o2111ai_4 _15166_ (.A1(_04365_),
    .A2(_04448_),
    .B1(_04452_),
    .C1(_04719_),
    .D1(_04720_),
    .Y(_04722_));
 sky130_fd_sc_hd__o211ai_4 _15167_ (.A1(_04451_),
    .A2(_04456_),
    .B1(_04717_),
    .C1(_04718_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand3_1 _15168_ (.A(_04586_),
    .B(_04722_),
    .C(_04723_),
    .Y(_04725_));
 sky130_fd_sc_hd__a21o_1 _15169_ (.A1(_04722_),
    .A2(_04723_),
    .B1(_04586_),
    .X(_04726_));
 sky130_fd_sc_hd__o211ai_4 _15170_ (.A1(_04584_),
    .A2(_04578_),
    .B1(_04583_),
    .C1(_04723_),
    .Y(_04727_));
 sky130_fd_sc_hd__a22o_1 _15171_ (.A1(_04583_),
    .A2(_04585_),
    .B1(_04722_),
    .B2(_04723_),
    .X(_04728_));
 sky130_fd_sc_hd__o221a_1 _15172_ (.A1(_04721_),
    .A2(_04727_),
    .B1(_04462_),
    .B2(_04466_),
    .C1(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__o221ai_4 _15173_ (.A1(_04721_),
    .A2(_04727_),
    .B1(_04462_),
    .B2(_04466_),
    .C1(_04728_),
    .Y(_04730_));
 sky130_fd_sc_hd__o2111ai_4 _15174_ (.A1(_04319_),
    .A2(_04458_),
    .B1(_04467_),
    .C1(_04725_),
    .D1(_04726_),
    .Y(_04731_));
 sky130_fd_sc_hd__o32a_2 _15175_ (.A1(_01802_),
    .A2(_02120_),
    .A3(_04106_),
    .B1(_02152_),
    .B2(_01846_),
    .X(_04732_));
 sky130_fd_sc_hd__o32a_2 _15176_ (.A1(_01846_),
    .A2(_02152_),
    .A3(_04188_),
    .B1(_04185_),
    .B2(_04107_),
    .X(_04733_));
 sky130_fd_sc_hd__o21a_1 _15177_ (.A1(_04063_),
    .A2(_04251_),
    .B1(_04250_),
    .X(_04734_));
 sky130_fd_sc_hd__a21oi_2 _15178_ (.A1(_04063_),
    .A2(_04251_),
    .B1(_04250_),
    .Y(_04736_));
 sky130_fd_sc_hd__nor2_1 _15179_ (.A(_04253_),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_1 _15180_ (.A(net12),
    .B(net51),
    .Y(_04738_));
 sky130_fd_sc_hd__nand2_2 _15181_ (.A(net26),
    .B(net49),
    .Y(_04739_));
 sky130_fd_sc_hd__and4_2 _15182_ (.A(net26),
    .B(net23),
    .C(net49),
    .D(net50),
    .X(_04740_));
 sky130_fd_sc_hd__nand4_4 _15183_ (.A(net26),
    .B(net23),
    .C(net49),
    .D(net50),
    .Y(_04741_));
 sky130_fd_sc_hd__o21a_1 _15184_ (.A1(_01791_),
    .A2(_02120_),
    .B1(_04185_),
    .X(_04742_));
 sky130_fd_sc_hd__nand2_2 _15185_ (.A(_04185_),
    .B(_04739_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _15186_ (.A(_04741_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__o211ai_1 _15187_ (.A1(_01824_),
    .A2(_02152_),
    .B1(_04741_),
    .C1(_04743_),
    .Y(_04745_));
 sky130_fd_sc_hd__a21o_1 _15188_ (.A1(_04741_),
    .A2(_04743_),
    .B1(_04738_),
    .X(_04747_));
 sky130_fd_sc_hd__nand4_4 _15189_ (.A(_04743_),
    .B(net51),
    .C(net12),
    .D(_04741_),
    .Y(_04748_));
 sky130_fd_sc_hd__o2bb2ai_2 _15190_ (.A1_N(_04741_),
    .A2_N(_04743_),
    .B1(_01824_),
    .B2(_02152_),
    .Y(_04749_));
 sky130_fd_sc_hd__a2bb2oi_1 _15191_ (.A1_N(_04253_),
    .A2_N(_04736_),
    .B1(_04738_),
    .B2(_04744_),
    .Y(_04750_));
 sky130_fd_sc_hd__o211a_1 _15192_ (.A1(_04253_),
    .A2(_04736_),
    .B1(_04748_),
    .C1(_04749_),
    .X(_04751_));
 sky130_fd_sc_hd__o211ai_4 _15193_ (.A1(_04253_),
    .A2(_04736_),
    .B1(_04748_),
    .C1(_04749_),
    .Y(_04752_));
 sky130_fd_sc_hd__a2bb2oi_2 _15194_ (.A1_N(_04252_),
    .A2_N(_04734_),
    .B1(_04748_),
    .B2(_04749_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand3_1 _15195_ (.A(_04737_),
    .B(_04745_),
    .C(_04747_),
    .Y(_04754_));
 sky130_fd_sc_hd__a31o_1 _15196_ (.A1(_04737_),
    .A2(_04745_),
    .A3(_04747_),
    .B1(_04733_),
    .X(_04755_));
 sky130_fd_sc_hd__a211oi_2 _15197_ (.A1(_04750_),
    .A2(_04748_),
    .B1(_04733_),
    .C1(_04753_),
    .Y(_04756_));
 sky130_fd_sc_hd__a2bb2oi_4 _15198_ (.A1_N(_04188_),
    .A2_N(_04732_),
    .B1(_04752_),
    .B2(_04754_),
    .Y(_04758_));
 sky130_fd_sc_hd__a2bb2o_1 _15199_ (.A1_N(_04188_),
    .A2_N(_04732_),
    .B1(_04752_),
    .B2(_04754_),
    .X(_04759_));
 sky130_fd_sc_hd__a21oi_1 _15200_ (.A1(_04247_),
    .A2(_04258_),
    .B1(_04248_),
    .Y(_04760_));
 sky130_fd_sc_hd__o21ai_4 _15201_ (.A1(_04756_),
    .A2(_04758_),
    .B1(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__o22ai_4 _15202_ (.A1(_04751_),
    .A2(_04755_),
    .B1(_04248_),
    .B2(_04259_),
    .Y(_04762_));
 sky130_fd_sc_hd__o221ai_2 _15203_ (.A1(_04751_),
    .A2(_04755_),
    .B1(_04248_),
    .B2(_04259_),
    .C1(_04759_),
    .Y(_04763_));
 sky130_fd_sc_hd__o31a_1 _15204_ (.A1(_01824_),
    .A2(_02120_),
    .A3(_04108_),
    .B1(_04196_),
    .X(_04764_));
 sky130_fd_sc_hd__a41o_2 _15205_ (.A1(_04199_),
    .A2(_03594_),
    .A3(net50),
    .A4(net12),
    .B1(_04195_),
    .X(_04765_));
 sky130_fd_sc_hd__o2bb2ai_2 _15206_ (.A1_N(_04761_),
    .A2_N(_04763_),
    .B1(_04764_),
    .B2(_04197_),
    .Y(_04766_));
 sky130_fd_sc_hd__o211ai_4 _15207_ (.A1(_04758_),
    .A2(_04762_),
    .B1(_04765_),
    .C1(_04761_),
    .Y(_04767_));
 sky130_fd_sc_hd__o31a_1 _15208_ (.A1(_04105_),
    .A2(_04109_),
    .A3(_04112_),
    .B1(_04206_),
    .X(_04769_));
 sky130_fd_sc_hd__o21ai_1 _15209_ (.A1(_04116_),
    .A2(_04207_),
    .B1(_04206_),
    .Y(_04770_));
 sky130_fd_sc_hd__a21oi_1 _15210_ (.A1(_04766_),
    .A2(_04767_),
    .B1(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__o2bb2ai_2 _15211_ (.A1_N(_04766_),
    .A2_N(_04767_),
    .B1(_04769_),
    .B2(_04207_),
    .Y(_04772_));
 sky130_fd_sc_hd__o211a_1 _15212_ (.A1(_04205_),
    .A2(_04211_),
    .B1(_04766_),
    .C1(_04767_),
    .X(_04773_));
 sky130_fd_sc_hd__o211ai_2 _15213_ (.A1(_04205_),
    .A2(_04211_),
    .B1(_04766_),
    .C1(_04767_),
    .Y(_04774_));
 sky130_fd_sc_hd__o22ai_4 _15214_ (.A1(_01846_),
    .A2(_02174_),
    .B1(_04771_),
    .B2(_04773_),
    .Y(_04775_));
 sky130_fd_sc_hd__nand4_4 _15215_ (.A(_04772_),
    .B(_04774_),
    .C(net1),
    .D(net52),
    .Y(_04776_));
 sky130_fd_sc_hd__o211a_1 _15216_ (.A1(_04301_),
    .A2(_04304_),
    .B1(_04044_),
    .C1(_04081_),
    .X(_04777_));
 sky130_fd_sc_hd__o22ai_1 _15217_ (.A1(_04301_),
    .A2(_04304_),
    .B1(_04309_),
    .B2(_04306_),
    .Y(_04778_));
 sky130_fd_sc_hd__a21oi_2 _15218_ (.A1(_04775_),
    .A2(_04776_),
    .B1(_04778_),
    .Y(_04780_));
 sky130_fd_sc_hd__o2bb2ai_4 _15219_ (.A1_N(_04775_),
    .A2_N(_04776_),
    .B1(_04777_),
    .B2(_04306_),
    .Y(_04781_));
 sky130_fd_sc_hd__o211a_4 _15220_ (.A1(_04305_),
    .A2(_04315_),
    .B1(_04775_),
    .C1(_04776_),
    .X(_04782_));
 sky130_fd_sc_hd__o211ai_4 _15221_ (.A1(_04305_),
    .A2(_04315_),
    .B1(_04775_),
    .C1(_04776_),
    .Y(_04783_));
 sky130_fd_sc_hd__a21oi_1 _15222_ (.A1(_04781_),
    .A2(_04783_),
    .B1(_04216_),
    .Y(_04784_));
 sky130_fd_sc_hd__o21ai_2 _15223_ (.A1(_04780_),
    .A2(_04782_),
    .B1(_04217_),
    .Y(_04785_));
 sky130_fd_sc_hd__nand2_2 _15224_ (.A(_04781_),
    .B(_04216_),
    .Y(_04786_));
 sky130_fd_sc_hd__inv_2 _15225_ (.A(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__and3_1 _15226_ (.A(_04781_),
    .B(_04783_),
    .C(_04216_),
    .X(_04788_));
 sky130_fd_sc_hd__nand3_1 _15227_ (.A(_04781_),
    .B(_04783_),
    .C(_04216_),
    .Y(_04789_));
 sky130_fd_sc_hd__a21oi_1 _15228_ (.A1(_04781_),
    .A2(_04783_),
    .B1(_04217_),
    .Y(_04791_));
 sky130_fd_sc_hd__o21ai_2 _15229_ (.A1(_04780_),
    .A2(_04782_),
    .B1(_04216_),
    .Y(_04792_));
 sky130_fd_sc_hd__nor3_1 _15230_ (.A(_04216_),
    .B(_04780_),
    .C(_04782_),
    .Y(_04793_));
 sky130_fd_sc_hd__nand3_2 _15231_ (.A(_04217_),
    .B(_04781_),
    .C(_04783_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand4_4 _15232_ (.A(_04730_),
    .B(_04731_),
    .C(_04792_),
    .D(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__o2bb2ai_2 _15233_ (.A1_N(_04730_),
    .A2_N(_04731_),
    .B1(_04791_),
    .B2(_04793_),
    .Y(_04796_));
 sky130_fd_sc_hd__o2bb2ai_2 _15234_ (.A1_N(_04730_),
    .A2_N(_04731_),
    .B1(_04784_),
    .B2(_04788_),
    .Y(_04797_));
 sky130_fd_sc_hd__o211ai_1 _15235_ (.A1(_04782_),
    .A2(_04786_),
    .B1(_04785_),
    .C1(_04731_),
    .Y(_04798_));
 sky130_fd_sc_hd__o2111ai_4 _15236_ (.A1(_04782_),
    .A2(_04786_),
    .B1(_04785_),
    .C1(_04730_),
    .D1(_04731_),
    .Y(_04799_));
 sky130_fd_sc_hd__o211a_2 _15237_ (.A1(_04729_),
    .A2(_04798_),
    .B1(_04797_),
    .C1(_04513_),
    .X(_04800_));
 sky130_fd_sc_hd__nand3_4 _15238_ (.A(_04513_),
    .B(_04797_),
    .C(_04799_),
    .Y(_04802_));
 sky130_fd_sc_hd__o211ai_4 _15239_ (.A1(_04473_),
    .A2(_04512_),
    .B1(_04795_),
    .C1(_04796_),
    .Y(_04803_));
 sky130_fd_sc_hd__a41oi_4 _15240_ (.A1(_04471_),
    .A2(_04478_),
    .A3(_04795_),
    .A4(_04796_),
    .B1(_04510_),
    .Y(_04804_));
 sky130_fd_sc_hd__o21ai_2 _15241_ (.A1(_04221_),
    .A2(_04229_),
    .B1(_04803_),
    .Y(_04805_));
 sky130_fd_sc_hd__o211a_1 _15242_ (.A1(_04221_),
    .A2(_04229_),
    .B1(_04802_),
    .C1(_04803_),
    .X(_04806_));
 sky130_fd_sc_hd__o211ai_1 _15243_ (.A1(_04221_),
    .A2(_04229_),
    .B1(_04802_),
    .C1(_04803_),
    .Y(_04807_));
 sky130_fd_sc_hd__a21oi_2 _15244_ (.A1(_04802_),
    .A2(_04803_),
    .B1(_04511_),
    .Y(_04808_));
 sky130_fd_sc_hd__a21o_1 _15245_ (.A1(_04802_),
    .A2(_04803_),
    .B1(_04511_),
    .X(_04809_));
 sky130_fd_sc_hd__a21oi_1 _15246_ (.A1(_04802_),
    .A2(_04804_),
    .B1(_04808_),
    .Y(_04810_));
 sky130_fd_sc_hd__o21ai_1 _15247_ (.A1(_04800_),
    .A2(_04805_),
    .B1(_04809_),
    .Y(_04811_));
 sky130_fd_sc_hd__a2bb2oi_1 _15248_ (.A1_N(_04480_),
    .A2_N(_04489_),
    .B1(_04807_),
    .B2(_04809_),
    .Y(_04813_));
 sky130_fd_sc_hd__o21ai_1 _15249_ (.A1(_04806_),
    .A2(_04808_),
    .B1(_04509_),
    .Y(_04814_));
 sky130_fd_sc_hd__a221oi_2 _15250_ (.A1(_04804_),
    .A2(_04802_),
    .B1(_04492_),
    .B2(_04484_),
    .C1(_04808_),
    .Y(_04815_));
 sky130_fd_sc_hd__o2111ai_4 _15251_ (.A1(_04805_),
    .A2(_04800_),
    .B1(_04490_),
    .C1(_04481_),
    .D1(_04809_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _15252_ (.A(_04814_),
    .B(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__o22ai_2 _15253_ (.A1(_04495_),
    .A2(_04496_),
    .B1(_04813_),
    .B2(_04815_),
    .Y(_04818_));
 sky130_fd_sc_hd__nand3_2 _15254_ (.A(_04498_),
    .B(_04814_),
    .C(_04816_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _15255_ (.A(_04818_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__o21ai_1 _15256_ (.A1(_04503_),
    .A2(_04507_),
    .B1(_04502_),
    .Y(_04821_));
 sky130_fd_sc_hd__xnor2_1 _15257_ (.A(_04820_),
    .B(_04821_),
    .Y(net84));
 sky130_fd_sc_hd__nand3_2 _15258_ (.A(_04730_),
    .B(_04792_),
    .C(_04794_),
    .Y(_04823_));
 sky130_fd_sc_hd__a31oi_1 _15259_ (.A1(_04731_),
    .A2(_04785_),
    .A3(_04789_),
    .B1(_04729_),
    .Y(_04824_));
 sky130_fd_sc_hd__a32oi_1 _15260_ (.A1(_04589_),
    .A2(_04664_),
    .A3(_04666_),
    .B1(_04712_),
    .B2(_04715_),
    .Y(_04825_));
 sky130_fd_sc_hd__a32oi_4 _15261_ (.A1(_04589_),
    .A2(_04664_),
    .A3(_04666_),
    .B1(_04668_),
    .B2(_04716_),
    .Y(_04826_));
 sky130_fd_sc_hd__a32o_1 _15262_ (.A1(_04589_),
    .A2(_04664_),
    .A3(_04666_),
    .B1(_04668_),
    .B2(_04716_),
    .X(_04827_));
 sky130_fd_sc_hd__o21a_1 _15263_ (.A1(_01835_),
    .A2(_02076_),
    .B1(_04639_),
    .X(_04828_));
 sky130_fd_sc_hd__o21ai_2 _15264_ (.A1(_04634_),
    .A2(_04635_),
    .B1(_04639_),
    .Y(_04829_));
 sky130_fd_sc_hd__nand2_1 _15265_ (.A(net63),
    .B(net13),
    .Y(_04830_));
 sky130_fd_sc_hd__nand2_1 _15266_ (.A(net62),
    .B(net15),
    .Y(_04831_));
 sky130_fd_sc_hd__and4_1 _15267_ (.A(net61),
    .B(net62),
    .C(net14),
    .D(net15),
    .X(_04832_));
 sky130_fd_sc_hd__nand4_4 _15268_ (.A(net61),
    .B(net62),
    .C(net14),
    .D(net15),
    .Y(_04834_));
 sky130_fd_sc_hd__a22oi_4 _15269_ (.A1(net62),
    .A2(net14),
    .B1(net15),
    .B2(net61),
    .Y(_04835_));
 sky130_fd_sc_hd__a22o_1 _15270_ (.A1(net62),
    .A2(net14),
    .B1(net15),
    .B2(net61),
    .X(_04836_));
 sky130_fd_sc_hd__a2bb2oi_1 _15271_ (.A1_N(_01890_),
    .A2_N(_02043_),
    .B1(_04834_),
    .B2(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__a22o_1 _15272_ (.A1(net63),
    .A2(net13),
    .B1(_04834_),
    .B2(_04836_),
    .X(_04838_));
 sky130_fd_sc_hd__nor3_4 _15273_ (.A(_04835_),
    .B(_04830_),
    .C(_04832_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand4_2 _15274_ (.A(_04836_),
    .B(net13),
    .C(net63),
    .D(_04834_),
    .Y(_04840_));
 sky130_fd_sc_hd__o22ai_4 _15275_ (.A1(_04635_),
    .A2(_04828_),
    .B1(_04837_),
    .B2(_04839_),
    .Y(_04841_));
 sky130_fd_sc_hd__nand2_2 _15276_ (.A(_04838_),
    .B(_04829_),
    .Y(_04842_));
 sky130_fd_sc_hd__and3_1 _15277_ (.A(_04838_),
    .B(_04840_),
    .C(_04829_),
    .X(_04843_));
 sky130_fd_sc_hd__nand3_4 _15278_ (.A(_04838_),
    .B(_04840_),
    .C(_04829_),
    .Y(_04845_));
 sky130_fd_sc_hd__o21a_1 _15279_ (.A1(_01890_),
    .A2(_02032_),
    .B1(_04597_),
    .X(_04846_));
 sky130_fd_sc_hd__a31o_2 _15280_ (.A1(_04595_),
    .A2(net11),
    .A3(net63),
    .B1(_04596_),
    .X(_04847_));
 sky130_fd_sc_hd__a21oi_2 _15281_ (.A1(_04841_),
    .A2(_04845_),
    .B1(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__o2bb2ai_2 _15282_ (.A1_N(_04841_),
    .A2_N(_04845_),
    .B1(_04846_),
    .B2(_04594_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_2 _15283_ (.A(_04841_),
    .B(_04847_),
    .Y(_04850_));
 sky130_fd_sc_hd__and3_1 _15284_ (.A(_04841_),
    .B(_04845_),
    .C(_04847_),
    .X(_04851_));
 sky130_fd_sc_hd__o211ai_4 _15285_ (.A1(_04839_),
    .A2(_04842_),
    .B1(_04847_),
    .C1(_04841_),
    .Y(_04852_));
 sky130_fd_sc_hd__o21ai_1 _15286_ (.A1(_04843_),
    .A2(_04850_),
    .B1(_04849_),
    .Y(_04853_));
 sky130_fd_sc_hd__o21ai_1 _15287_ (.A1(_04372_),
    .A2(_04621_),
    .B1(_04618_),
    .Y(_04854_));
 sky130_fd_sc_hd__o22ai_2 _15288_ (.A1(_04372_),
    .A2(_04621_),
    .B1(_04618_),
    .B2(_04619_),
    .Y(_04856_));
 sky130_fd_sc_hd__o22a_1 _15289_ (.A1(_04372_),
    .A2(_04621_),
    .B1(_04618_),
    .B2(_04619_),
    .X(_04857_));
 sky130_fd_sc_hd__nand2_1 _15290_ (.A(net55),
    .B(net19),
    .Y(_04858_));
 sky130_fd_sc_hd__a22oi_4 _15291_ (.A1(net44),
    .A2(net20),
    .B1(net21),
    .B2(net33),
    .Y(_04859_));
 sky130_fd_sc_hd__a22o_2 _15292_ (.A1(net44),
    .A2(net20),
    .B1(net21),
    .B2(net33),
    .X(_04860_));
 sky130_fd_sc_hd__and4_1 _15293_ (.A(net33),
    .B(net44),
    .C(net20),
    .D(net21),
    .X(_04861_));
 sky130_fd_sc_hd__nand4_4 _15294_ (.A(net33),
    .B(net44),
    .C(net20),
    .D(net21),
    .Y(_04862_));
 sky130_fd_sc_hd__o211ai_4 _15295_ (.A1(_01780_),
    .A2(_02142_),
    .B1(_04860_),
    .C1(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__o21bai_2 _15296_ (.A1(_04859_),
    .A2(_04861_),
    .B1_N(_04858_),
    .Y(_04864_));
 sky130_fd_sc_hd__o22a_2 _15297_ (.A1(_01780_),
    .A2(_02142_),
    .B1(_04859_),
    .B2(_04861_),
    .X(_04865_));
 sky130_fd_sc_hd__o21ai_2 _15298_ (.A1(_04859_),
    .A2(_04861_),
    .B1(_04858_),
    .Y(_04867_));
 sky130_fd_sc_hd__nand4_4 _15299_ (.A(_04860_),
    .B(_04862_),
    .C(net55),
    .D(net19),
    .Y(_04868_));
 sky130_fd_sc_hd__a22oi_4 _15300_ (.A1(_04620_),
    .A2(_04854_),
    .B1(_04867_),
    .B2(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand3_4 _15301_ (.A(_04857_),
    .B(_04863_),
    .C(_04864_),
    .Y(_04870_));
 sky130_fd_sc_hd__nand2_2 _15302_ (.A(_04868_),
    .B(_04856_),
    .Y(_04871_));
 sky130_fd_sc_hd__a21oi_1 _15303_ (.A1(_04863_),
    .A2(_04864_),
    .B1(_04857_),
    .Y(_04872_));
 sky130_fd_sc_hd__nand3_1 _15304_ (.A(_04867_),
    .B(_04868_),
    .C(_04856_),
    .Y(_04873_));
 sky130_fd_sc_hd__nand2_1 _15305_ (.A(net60),
    .B(net16),
    .Y(_04874_));
 sky130_fd_sc_hd__a22oi_4 _15306_ (.A1(net59),
    .A2(net17),
    .B1(net18),
    .B2(net58),
    .Y(_04875_));
 sky130_fd_sc_hd__a22o_1 _15307_ (.A1(net59),
    .A2(net17),
    .B1(net18),
    .B2(net58),
    .X(_04876_));
 sky130_fd_sc_hd__and4_1 _15308_ (.A(net58),
    .B(net59),
    .C(net17),
    .D(net18),
    .X(_04878_));
 sky130_fd_sc_hd__nand4_4 _15309_ (.A(net58),
    .B(net59),
    .C(net17),
    .D(net18),
    .Y(_04879_));
 sky130_fd_sc_hd__and3_1 _15310_ (.A(_04874_),
    .B(_04876_),
    .C(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__o211ai_2 _15311_ (.A1(_01835_),
    .A2(_02098_),
    .B1(_04876_),
    .C1(_04879_),
    .Y(_04881_));
 sky130_fd_sc_hd__o211a_1 _15312_ (.A1(_04875_),
    .A2(_04878_),
    .B1(net60),
    .C1(net16),
    .X(_04882_));
 sky130_fd_sc_hd__a21o_1 _15313_ (.A1(_04876_),
    .A2(_04879_),
    .B1(_04874_),
    .X(_04883_));
 sky130_fd_sc_hd__o22a_1 _15314_ (.A1(_01835_),
    .A2(_02098_),
    .B1(_04875_),
    .B2(_04878_),
    .X(_04884_));
 sky130_fd_sc_hd__a22o_1 _15315_ (.A1(net60),
    .A2(net16),
    .B1(_04876_),
    .B2(_04879_),
    .X(_04885_));
 sky130_fd_sc_hd__a41o_1 _15316_ (.A1(net58),
    .A2(net59),
    .A3(net17),
    .A4(net18),
    .B1(_04874_),
    .X(_04886_));
 sky130_fd_sc_hd__and4_1 _15317_ (.A(_04876_),
    .B(_04879_),
    .C(net60),
    .D(net16),
    .X(_04887_));
 sky130_fd_sc_hd__o21ai_1 _15318_ (.A1(_04875_),
    .A2(_04886_),
    .B1(_04885_),
    .Y(_04889_));
 sky130_fd_sc_hd__nand2_1 _15319_ (.A(_04881_),
    .B(_04883_),
    .Y(_04890_));
 sky130_fd_sc_hd__o2bb2ai_2 _15320_ (.A1_N(_04881_),
    .A2_N(_04883_),
    .B1(_04865_),
    .B2(_04871_),
    .Y(_04891_));
 sky130_fd_sc_hd__o2bb2ai_2 _15321_ (.A1_N(_04870_),
    .A2_N(_04873_),
    .B1(_04884_),
    .B2(_04887_),
    .Y(_04892_));
 sky130_fd_sc_hd__o221ai_4 _15322_ (.A1(_04884_),
    .A2(_04887_),
    .B1(_04865_),
    .B2(_04871_),
    .C1(_04870_),
    .Y(_04893_));
 sky130_fd_sc_hd__o2bb2ai_2 _15323_ (.A1_N(_04870_),
    .A2_N(_04873_),
    .B1(_04880_),
    .B2(_04882_),
    .Y(_04894_));
 sky130_fd_sc_hd__nand2_1 _15324_ (.A(_04893_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__o21ai_1 _15325_ (.A1(_04869_),
    .A2(_04891_),
    .B1(_04892_),
    .Y(_04896_));
 sky130_fd_sc_hd__a32oi_4 _15326_ (.A1(_04615_),
    .A2(_04628_),
    .A3(_04629_),
    .B1(_04631_),
    .B2(_04650_),
    .Y(_04897_));
 sky130_fd_sc_hd__o22ai_4 _15327_ (.A1(_04627_),
    .A2(_04632_),
    .B1(_04649_),
    .B2(_04630_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand3_4 _15328_ (.A(_04897_),
    .B(_04894_),
    .C(_04893_),
    .Y(_04900_));
 sky130_fd_sc_hd__o211a_2 _15329_ (.A1(_04891_),
    .A2(_04869_),
    .B1(_04898_),
    .C1(_04892_),
    .X(_04901_));
 sky130_fd_sc_hd__o211ai_4 _15330_ (.A1(_04891_),
    .A2(_04869_),
    .B1(_04898_),
    .C1(_04892_),
    .Y(_04902_));
 sky130_fd_sc_hd__a22o_1 _15331_ (.A1(_04849_),
    .A2(_04852_),
    .B1(_04900_),
    .B2(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__a21oi_2 _15332_ (.A1(_04896_),
    .A2(_04897_),
    .B1(_04853_),
    .Y(_04904_));
 sky130_fd_sc_hd__o211ai_2 _15333_ (.A1(_04850_),
    .A2(_04843_),
    .B1(_04849_),
    .C1(_04900_),
    .Y(_04905_));
 sky130_fd_sc_hd__o211ai_4 _15334_ (.A1(_04848_),
    .A2(_04851_),
    .B1(_04900_),
    .C1(_04902_),
    .Y(_04906_));
 sky130_fd_sc_hd__a21o_1 _15335_ (.A1(_04900_),
    .A2(_04902_),
    .B1(_04853_),
    .X(_04907_));
 sky130_fd_sc_hd__a32oi_4 _15336_ (.A1(_04653_),
    .A2(_04655_),
    .A3(_04654_),
    .B1(_04612_),
    .B2(_04661_),
    .Y(_04908_));
 sky130_fd_sc_hd__a32o_1 _15337_ (.A1(_04653_),
    .A2(_04655_),
    .A3(_04654_),
    .B1(_04612_),
    .B2(_04661_),
    .X(_04909_));
 sky130_fd_sc_hd__o2111ai_4 _15338_ (.A1(_04612_),
    .A2(_04657_),
    .B1(_04661_),
    .C1(_04906_),
    .D1(_04907_),
    .Y(_04911_));
 sky130_fd_sc_hd__o211ai_4 _15339_ (.A1(_04901_),
    .A2(_04905_),
    .B1(_04908_),
    .C1(_04903_),
    .Y(_04912_));
 sky130_fd_sc_hd__a21oi_2 _15340_ (.A1(_04602_),
    .A2(_04607_),
    .B1(_04604_),
    .Y(_04913_));
 sky130_fd_sc_hd__o21a_1 _15341_ (.A1(_01934_),
    .A2(_01988_),
    .B1(_04677_),
    .X(_04914_));
 sky130_fd_sc_hd__a31o_2 _15342_ (.A1(_04675_),
    .A2(net8),
    .A3(net35),
    .B1(_04676_),
    .X(_04915_));
 sky130_fd_sc_hd__and2_1 _15343_ (.A(net35),
    .B(net9),
    .X(_04916_));
 sky130_fd_sc_hd__nand2_1 _15344_ (.A(net34),
    .B(net11),
    .Y(_04917_));
 sky130_fd_sc_hd__nand4_2 _15345_ (.A(net64),
    .B(net34),
    .C(net10),
    .D(net11),
    .Y(_04918_));
 sky130_fd_sc_hd__a22o_2 _15346_ (.A1(net34),
    .A2(net10),
    .B1(net11),
    .B2(net64),
    .X(_04919_));
 sky130_fd_sc_hd__a22oi_2 _15347_ (.A1(net35),
    .A2(net9),
    .B1(_04918_),
    .B2(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__a22o_2 _15348_ (.A1(net35),
    .A2(net9),
    .B1(_04918_),
    .B2(_04919_),
    .X(_04922_));
 sky130_fd_sc_hd__o211a_1 _15349_ (.A1(_04673_),
    .A2(_04917_),
    .B1(_04916_),
    .C1(_04919_),
    .X(_04923_));
 sky130_fd_sc_hd__o2111ai_4 _15350_ (.A1(_04673_),
    .A2(_04917_),
    .B1(net35),
    .C1(net9),
    .D1(_04919_),
    .Y(_04924_));
 sky130_fd_sc_hd__o22ai_4 _15351_ (.A1(_04674_),
    .A2(_04914_),
    .B1(_04920_),
    .B2(_04923_),
    .Y(_04925_));
 sky130_fd_sc_hd__nand3_4 _15352_ (.A(_04915_),
    .B(_04922_),
    .C(_04924_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand2_1 _15353_ (.A(net6),
    .B(net38),
    .Y(_04927_));
 sky130_fd_sc_hd__a22oi_4 _15354_ (.A1(net37),
    .A2(net7),
    .B1(net8),
    .B2(net36),
    .Y(_04928_));
 sky130_fd_sc_hd__and4_1 _15355_ (.A(net36),
    .B(net37),
    .C(net7),
    .D(net8),
    .X(_04929_));
 sky130_fd_sc_hd__nand4_1 _15356_ (.A(net36),
    .B(net37),
    .C(net7),
    .D(net8),
    .Y(_04930_));
 sky130_fd_sc_hd__a211oi_2 _15357_ (.A1(net6),
    .A2(net38),
    .B1(_04928_),
    .C1(_04929_),
    .Y(_04931_));
 sky130_fd_sc_hd__a211o_1 _15358_ (.A1(net6),
    .A2(net38),
    .B1(_04928_),
    .C1(_04929_),
    .X(_04933_));
 sky130_fd_sc_hd__o211a_1 _15359_ (.A1(_04928_),
    .A2(_04929_),
    .B1(net6),
    .C1(net38),
    .X(_04934_));
 sky130_fd_sc_hd__o211ai_1 _15360_ (.A1(_04928_),
    .A2(_04929_),
    .B1(net6),
    .C1(net38),
    .Y(_04935_));
 sky130_fd_sc_hd__o2bb2a_1 _15361_ (.A1_N(net6),
    .A2_N(net38),
    .B1(_04928_),
    .B2(_04929_),
    .X(_04936_));
 sky130_fd_sc_hd__and4b_2 _15362_ (.A_N(_04928_),
    .B(_04930_),
    .C(net6),
    .D(net38),
    .X(_04937_));
 sky130_fd_sc_hd__nand2_1 _15363_ (.A(_04933_),
    .B(_04935_),
    .Y(_04938_));
 sky130_fd_sc_hd__and3_1 _15364_ (.A(_04925_),
    .B(_04926_),
    .C(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__o211ai_2 _15365_ (.A1(_04931_),
    .A2(_04934_),
    .B1(_04925_),
    .C1(_04926_),
    .Y(_04940_));
 sky130_fd_sc_hd__o2bb2ai_2 _15366_ (.A1_N(_04925_),
    .A2_N(_04926_),
    .B1(_04936_),
    .B2(_04937_),
    .Y(_04941_));
 sky130_fd_sc_hd__o211ai_4 _15367_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04925_),
    .C1(_04926_),
    .Y(_04942_));
 sky130_fd_sc_hd__o2bb2ai_2 _15368_ (.A1_N(_04925_),
    .A2_N(_04926_),
    .B1(_04931_),
    .B2(_04934_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand3_4 _15369_ (.A(_04944_),
    .B(_04913_),
    .C(_04942_),
    .Y(_04945_));
 sky130_fd_sc_hd__o21ai_1 _15370_ (.A1(_04604_),
    .A2(_04609_),
    .B1(_04941_),
    .Y(_04946_));
 sky130_fd_sc_hd__o211a_2 _15371_ (.A1(_04604_),
    .A2(_04609_),
    .B1(_04940_),
    .C1(_04941_),
    .X(_04947_));
 sky130_fd_sc_hd__o211ai_4 _15372_ (.A1(_04604_),
    .A2(_04609_),
    .B1(_04940_),
    .C1(_04941_),
    .Y(_04948_));
 sky130_fd_sc_hd__o21ai_4 _15373_ (.A1(_04693_),
    .A2(_04681_),
    .B1(_04684_),
    .Y(_04949_));
 sky130_fd_sc_hd__a21oi_4 _15374_ (.A1(_04945_),
    .A2(_04948_),
    .B1(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__a21o_1 _15375_ (.A1(_04945_),
    .A2(_04948_),
    .B1(_04949_),
    .X(_04951_));
 sky130_fd_sc_hd__a32oi_1 _15376_ (.A1(_04944_),
    .A2(_04913_),
    .A3(_04942_),
    .B1(_04697_),
    .B2(_04684_),
    .Y(_04952_));
 sky130_fd_sc_hd__a32o_1 _15377_ (.A1(_04944_),
    .A2(_04913_),
    .A3(_04942_),
    .B1(_04697_),
    .B2(_04684_),
    .X(_04953_));
 sky130_fd_sc_hd__and3_2 _15378_ (.A(_04945_),
    .B(_04948_),
    .C(_04949_),
    .X(_04955_));
 sky130_fd_sc_hd__a21oi_1 _15379_ (.A1(_04948_),
    .A2(_04952_),
    .B1(_04950_),
    .Y(_04956_));
 sky130_fd_sc_hd__o21ai_2 _15380_ (.A1(_04947_),
    .A2(_04953_),
    .B1(_04951_),
    .Y(_04957_));
 sky130_fd_sc_hd__o2111a_1 _15381_ (.A1(_04947_),
    .A2(_04953_),
    .B1(_04951_),
    .C1(_04911_),
    .D1(_04912_),
    .X(_04958_));
 sky130_fd_sc_hd__o2111ai_4 _15382_ (.A1(_04947_),
    .A2(_04953_),
    .B1(_04951_),
    .C1(_04911_),
    .D1(_04912_),
    .Y(_04959_));
 sky130_fd_sc_hd__o2bb2a_1 _15383_ (.A1_N(_04911_),
    .A2_N(_04912_),
    .B1(_04950_),
    .B2(_04955_),
    .X(_04960_));
 sky130_fd_sc_hd__o2bb2ai_2 _15384_ (.A1_N(_04911_),
    .A2_N(_04912_),
    .B1(_04950_),
    .B2(_04955_),
    .Y(_04961_));
 sky130_fd_sc_hd__a21o_1 _15385_ (.A1(_04911_),
    .A2(_04912_),
    .B1(_04957_),
    .X(_04962_));
 sky130_fd_sc_hd__o211ai_4 _15386_ (.A1(_04950_),
    .A2(_04955_),
    .B1(_04911_),
    .C1(_04912_),
    .Y(_04963_));
 sky130_fd_sc_hd__a2bb2oi_1 _15387_ (.A1_N(_04667_),
    .A2_N(_04825_),
    .B1(_04959_),
    .B2(_04961_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand3_4 _15388_ (.A(_04962_),
    .B(_04963_),
    .C(_04826_),
    .Y(_04966_));
 sky130_fd_sc_hd__a21oi_4 _15389_ (.A1(_04962_),
    .A2(_04963_),
    .B1(_04826_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand3_2 _15390_ (.A(_04827_),
    .B(_04959_),
    .C(_04961_),
    .Y(_04968_));
 sky130_fd_sc_hd__o311a_1 _15391_ (.A1(_01912_),
    .A2(_02010_),
    .A3(_04275_),
    .B1(_04279_),
    .C1(_04533_),
    .X(_04969_));
 sky130_fd_sc_hd__o21ai_1 _15392_ (.A1(_04518_),
    .A2(_04534_),
    .B1(_04533_),
    .Y(_04970_));
 sky130_fd_sc_hd__and3_1 _15393_ (.A(_04525_),
    .B(net41),
    .C(net2),
    .X(_04971_));
 sky130_fd_sc_hd__a31o_1 _15394_ (.A1(_04525_),
    .A2(net41),
    .A3(net2),
    .B1(_04523_),
    .X(_04972_));
 sky130_fd_sc_hd__o21ai_1 _15395_ (.A1(_04688_),
    .A2(_04685_),
    .B1(_04687_),
    .Y(_04973_));
 sky130_fd_sc_hd__o21a_1 _15396_ (.A1(_04688_),
    .A2(_04685_),
    .B1(_04687_),
    .X(_04974_));
 sky130_fd_sc_hd__nand2_1 _15397_ (.A(net3),
    .B(net41),
    .Y(_04975_));
 sky130_fd_sc_hd__a22oi_4 _15398_ (.A1(net5),
    .A2(net39),
    .B1(net40),
    .B2(net4),
    .Y(_04977_));
 sky130_fd_sc_hd__a22o_1 _15399_ (.A1(net5),
    .A2(net39),
    .B1(net40),
    .B2(net4),
    .X(_04978_));
 sky130_fd_sc_hd__and4_1 _15400_ (.A(net4),
    .B(net5),
    .C(net39),
    .D(net40),
    .X(_04979_));
 sky130_fd_sc_hd__nand4_2 _15401_ (.A(net4),
    .B(net5),
    .C(net39),
    .D(net40),
    .Y(_04980_));
 sky130_fd_sc_hd__o211ai_1 _15402_ (.A1(_01923_),
    .A2(_02010_),
    .B1(_04978_),
    .C1(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__o21bai_1 _15403_ (.A1(_04977_),
    .A2(_04979_),
    .B1_N(_04975_),
    .Y(_04982_));
 sky130_fd_sc_hd__o21ai_1 _15404_ (.A1(_04977_),
    .A2(_04979_),
    .B1(_04975_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand4_1 _15405_ (.A(_04978_),
    .B(_04980_),
    .C(net3),
    .D(net41),
    .Y(_04984_));
 sky130_fd_sc_hd__nand2_1 _15406_ (.A(_04983_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__and3_1 _15407_ (.A(_04983_),
    .B(_04984_),
    .C(_04973_),
    .X(_04986_));
 sky130_fd_sc_hd__nand3_1 _15408_ (.A(_04983_),
    .B(_04984_),
    .C(_04973_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand3_2 _15409_ (.A(_04974_),
    .B(_04981_),
    .C(_04982_),
    .Y(_04989_));
 sky130_fd_sc_hd__o21ai_2 _15410_ (.A1(_04523_),
    .A2(_04971_),
    .B1(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__o211a_1 _15411_ (.A1(_04523_),
    .A2(_04971_),
    .B1(_04988_),
    .C1(_04989_),
    .X(_04991_));
 sky130_fd_sc_hd__a21oi_2 _15412_ (.A1(_04988_),
    .A2(_04989_),
    .B1(_04972_),
    .Y(_04992_));
 sky130_fd_sc_hd__a21o_1 _15413_ (.A1(_04988_),
    .A2(_04989_),
    .B1(_04972_),
    .X(_04993_));
 sky130_fd_sc_hd__o211ai_4 _15414_ (.A1(_04986_),
    .A2(_04990_),
    .B1(_04970_),
    .C1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__o221a_1 _15415_ (.A1(_04518_),
    .A2(_04534_),
    .B1(_04991_),
    .B2(_04992_),
    .C1(_04533_),
    .X(_04995_));
 sky130_fd_sc_hd__o22ai_4 _15416_ (.A1(_04534_),
    .A2(_04969_),
    .B1(_04991_),
    .B2(_04992_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _15417_ (.A(net28),
    .B(net48),
    .Y(_04997_));
 sky130_fd_sc_hd__nand2_1 _15418_ (.A(net30),
    .B(net46),
    .Y(_04999_));
 sky130_fd_sc_hd__and4_2 _15419_ (.A(net29),
    .B(net30),
    .C(net46),
    .D(net47),
    .X(_05000_));
 sky130_fd_sc_hd__nand4_1 _15420_ (.A(net29),
    .B(net30),
    .C(net46),
    .D(net47),
    .Y(_05001_));
 sky130_fd_sc_hd__a22oi_1 _15421_ (.A1(net30),
    .A2(net46),
    .B1(net47),
    .B2(net29),
    .Y(_05002_));
 sky130_fd_sc_hd__nand3_2 _15422_ (.A(_04999_),
    .B(net47),
    .C(net29),
    .Y(_05003_));
 sky130_fd_sc_hd__nand3_2 _15423_ (.A(_04557_),
    .B(net46),
    .C(net30),
    .Y(_05004_));
 sky130_fd_sc_hd__a22oi_4 _15424_ (.A1(net28),
    .A2(net48),
    .B1(_05003_),
    .B2(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__and4_4 _15425_ (.A(_05003_),
    .B(_05004_),
    .C(net28),
    .D(net48),
    .X(_05006_));
 sky130_fd_sc_hd__a31o_1 _15426_ (.A1(_04546_),
    .A2(net45),
    .A3(net30),
    .B1(_04547_),
    .X(_05007_));
 sky130_fd_sc_hd__o31a_2 _15427_ (.A1(_01868_),
    .A2(_02054_),
    .A3(_04545_),
    .B1(_04549_),
    .X(_05008_));
 sky130_fd_sc_hd__nand2_1 _15428_ (.A(net31),
    .B(net45),
    .Y(_05010_));
 sky130_fd_sc_hd__and4_1 _15429_ (.A(net2),
    .B(net32),
    .C(net42),
    .D(net43),
    .X(_05011_));
 sky130_fd_sc_hd__nand4_2 _15430_ (.A(net2),
    .B(net32),
    .C(net42),
    .D(net43),
    .Y(_05012_));
 sky130_fd_sc_hd__a22oi_4 _15431_ (.A1(net2),
    .A2(net42),
    .B1(net43),
    .B2(net32),
    .Y(_05013_));
 sky130_fd_sc_hd__a22o_1 _15432_ (.A1(net2),
    .A2(net42),
    .B1(net43),
    .B2(net32),
    .X(_05014_));
 sky130_fd_sc_hd__o211ai_2 _15433_ (.A1(_01879_),
    .A2(_02054_),
    .B1(_05012_),
    .C1(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__a21o_1 _15434_ (.A1(_05012_),
    .A2(_05014_),
    .B1(_05010_),
    .X(_05016_));
 sky130_fd_sc_hd__o22ai_4 _15435_ (.A1(_01879_),
    .A2(_02054_),
    .B1(_05011_),
    .B2(_05013_),
    .Y(_05017_));
 sky130_fd_sc_hd__a41o_2 _15436_ (.A1(net2),
    .A2(net32),
    .A3(net42),
    .A4(net43),
    .B1(_05010_),
    .X(_05018_));
 sky130_fd_sc_hd__o21ai_2 _15437_ (.A1(_05013_),
    .A2(_05018_),
    .B1(_05017_),
    .Y(_05019_));
 sky130_fd_sc_hd__o211a_4 _15438_ (.A1(_05013_),
    .A2(_05018_),
    .B1(_05017_),
    .C1(_05007_),
    .X(_05021_));
 sky130_fd_sc_hd__o211ai_4 _15439_ (.A1(_05013_),
    .A2(_05018_),
    .B1(_05017_),
    .C1(_05007_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand3_4 _15440_ (.A(_05008_),
    .B(_05015_),
    .C(_05016_),
    .Y(_05023_));
 sky130_fd_sc_hd__a2bb2oi_1 _15441_ (.A1_N(_05005_),
    .A2_N(_05006_),
    .B1(_05022_),
    .B2(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__and4bb_1 _15442_ (.A_N(_05005_),
    .B_N(_05006_),
    .C(_05022_),
    .D(_05023_),
    .X(_05025_));
 sky130_fd_sc_hd__a2bb2oi_2 _15443_ (.A1_N(_05005_),
    .A2_N(_05006_),
    .B1(_05008_),
    .B2(_05019_),
    .Y(_05026_));
 sky130_fd_sc_hd__o21ai_4 _15444_ (.A1(_05005_),
    .A2(_05006_),
    .B1(_05023_),
    .Y(_05027_));
 sky130_fd_sc_hd__o211a_2 _15445_ (.A1(_05005_),
    .A2(_05006_),
    .B1(_05022_),
    .C1(_05023_),
    .X(_05028_));
 sky130_fd_sc_hd__a211oi_4 _15446_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_05005_),
    .C1(_05006_),
    .Y(_05029_));
 sky130_fd_sc_hd__a211o_1 _15447_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_05005_),
    .C1(_05006_),
    .X(_05030_));
 sky130_fd_sc_hd__o21ai_1 _15448_ (.A1(_05021_),
    .A2(_05027_),
    .B1(_05030_),
    .Y(_05032_));
 sky130_fd_sc_hd__o2bb2ai_4 _15449_ (.A1_N(_04994_),
    .A2_N(_04996_),
    .B1(_05028_),
    .B2(_05029_),
    .Y(_05033_));
 sky130_fd_sc_hd__o2111ai_4 _15450_ (.A1(_05021_),
    .A2(_05027_),
    .B1(_05030_),
    .C1(_04996_),
    .D1(_04994_),
    .Y(_05034_));
 sky130_fd_sc_hd__o211ai_4 _15451_ (.A1(_05028_),
    .A2(_05029_),
    .B1(_04994_),
    .C1(_04996_),
    .Y(_05035_));
 sky130_fd_sc_hd__o2bb2ai_2 _15452_ (.A1_N(_04994_),
    .A2_N(_04996_),
    .B1(_05024_),
    .B2(_05025_),
    .Y(_05036_));
 sky130_fd_sc_hd__a32oi_4 _15453_ (.A1(_04694_),
    .A2(_04695_),
    .A3(_04699_),
    .B1(_04704_),
    .B2(_04705_),
    .Y(_05037_));
 sky130_fd_sc_hd__a21oi_2 _15454_ (.A1(_04701_),
    .A2(_04706_),
    .B1(_04703_),
    .Y(_05038_));
 sky130_fd_sc_hd__a21oi_2 _15455_ (.A1(_05033_),
    .A2(_05034_),
    .B1(_05037_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand3_1 _15456_ (.A(_05035_),
    .B(_05036_),
    .C(_05038_),
    .Y(_05040_));
 sky130_fd_sc_hd__and3_2 _15457_ (.A(_05033_),
    .B(_05034_),
    .C(_05037_),
    .X(_05041_));
 sky130_fd_sc_hd__nand3_2 _15458_ (.A(_05033_),
    .B(_05034_),
    .C(_05037_),
    .Y(_05043_));
 sky130_fd_sc_hd__a31oi_4 _15459_ (.A1(_04543_),
    .A2(_04566_),
    .A3(_04568_),
    .B1(_04541_),
    .Y(_05044_));
 sky130_fd_sc_hd__a31o_1 _15460_ (.A1(_04543_),
    .A2(_04566_),
    .A3(_04568_),
    .B1(_04541_),
    .X(_05045_));
 sky130_fd_sc_hd__a21oi_2 _15461_ (.A1(_05040_),
    .A2(_05043_),
    .B1(_05044_),
    .Y(_05046_));
 sky130_fd_sc_hd__a22o_1 _15462_ (.A1(_04542_),
    .A2(_04571_),
    .B1(_05040_),
    .B2(_05043_),
    .X(_05047_));
 sky130_fd_sc_hd__a31oi_4 _15463_ (.A1(_05035_),
    .A2(_05036_),
    .A3(_05038_),
    .B1(_05045_),
    .Y(_05048_));
 sky130_fd_sc_hd__a31o_1 _15464_ (.A1(_05035_),
    .A2(_05036_),
    .A3(_05038_),
    .B1(_05045_),
    .X(_05049_));
 sky130_fd_sc_hd__and3_1 _15465_ (.A(_05040_),
    .B(_05043_),
    .C(_05044_),
    .X(_05050_));
 sky130_fd_sc_hd__o211a_1 _15466_ (.A1(_05039_),
    .A2(_05041_),
    .B1(_04542_),
    .C1(_04571_),
    .X(_05051_));
 sky130_fd_sc_hd__and3_1 _15467_ (.A(_05040_),
    .B(_05043_),
    .C(_05045_),
    .X(_05052_));
 sky130_fd_sc_hd__a21oi_4 _15468_ (.A1(_05043_),
    .A2(_05048_),
    .B1(_05046_),
    .Y(_05054_));
 sky130_fd_sc_hd__o21ai_2 _15469_ (.A1(_05041_),
    .A2(_05049_),
    .B1(_05047_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_1 _15470_ (.A(_04966_),
    .B(_05054_),
    .Y(_05056_));
 sky130_fd_sc_hd__o2bb2ai_1 _15471_ (.A1_N(_04966_),
    .A2_N(_04968_),
    .B1(_05046_),
    .B2(_05050_),
    .Y(_05057_));
 sky130_fd_sc_hd__o211ai_2 _15472_ (.A1(_05046_),
    .A2(_05050_),
    .B1(_04966_),
    .C1(_04968_),
    .Y(_05058_));
 sky130_fd_sc_hd__o2bb2ai_1 _15473_ (.A1_N(_04966_),
    .A2_N(_04968_),
    .B1(_05051_),
    .B2(_05052_),
    .Y(_05059_));
 sky130_fd_sc_hd__a32oi_4 _15474_ (.A1(_04587_),
    .A2(_04719_),
    .A3(_04720_),
    .B1(_04723_),
    .B2(_04586_),
    .Y(_05060_));
 sky130_fd_sc_hd__o2111ai_4 _15475_ (.A1(_04586_),
    .A2(_04721_),
    .B1(_04723_),
    .C1(_05058_),
    .D1(_05059_),
    .Y(_05061_));
 sky130_fd_sc_hd__o211ai_4 _15476_ (.A1(_04967_),
    .A2(_05056_),
    .B1(_05060_),
    .C1(_05057_),
    .Y(_05062_));
 sky130_fd_sc_hd__a2bb2oi_1 _15477_ (.A1_N(_04758_),
    .A2_N(_04762_),
    .B1(_04765_),
    .B2(_04761_),
    .Y(_05063_));
 sky130_fd_sc_hd__o2bb2ai_2 _15478_ (.A1_N(_04765_),
    .A2_N(_04761_),
    .B1(_04758_),
    .B2(_04762_),
    .Y(_05065_));
 sky130_fd_sc_hd__and3_1 _15479_ (.A(_04554_),
    .B(_04560_),
    .C(_04561_),
    .X(_05066_));
 sky130_fd_sc_hd__a31oi_2 _15480_ (.A1(_04554_),
    .A2(_04560_),
    .A3(_04561_),
    .B1(_04552_),
    .Y(_05067_));
 sky130_fd_sc_hd__o22a_1 _15481_ (.A1(_01769_),
    .A2(_02109_),
    .B1(_04251_),
    .B2(_04557_),
    .X(_05068_));
 sky130_fd_sc_hd__o22ai_1 _15482_ (.A1(_04251_),
    .A2(_04557_),
    .B1(_04555_),
    .B2(_04556_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_2 _15483_ (.A(net27),
    .B(net50),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2_2 _15484_ (.A(net27),
    .B(net49),
    .Y(_05071_));
 sky130_fd_sc_hd__and4_2 _15485_ (.A(net27),
    .B(net26),
    .C(net49),
    .D(net50),
    .X(_05072_));
 sky130_fd_sc_hd__nand4_1 _15486_ (.A(net27),
    .B(net26),
    .C(net49),
    .D(net50),
    .Y(_05073_));
 sky130_fd_sc_hd__a22oi_2 _15487_ (.A1(net27),
    .A2(net49),
    .B1(net50),
    .B2(net26),
    .Y(_05074_));
 sky130_fd_sc_hd__a22o_1 _15488_ (.A1(net27),
    .A2(net49),
    .B1(net50),
    .B2(net26),
    .X(_05076_));
 sky130_fd_sc_hd__a2bb2oi_2 _15489_ (.A1_N(_01802_),
    .A2_N(_02152_),
    .B1(_05073_),
    .B2(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__o22ai_1 _15490_ (.A1(_01802_),
    .A2(_02152_),
    .B1(_05072_),
    .B2(_05074_),
    .Y(_05078_));
 sky130_fd_sc_hd__o2111a_1 _15491_ (.A1(_04739_),
    .A2(_05070_),
    .B1(net23),
    .C1(net51),
    .D1(_05076_),
    .X(_05079_));
 sky130_fd_sc_hd__o2111ai_2 _15492_ (.A1(_04739_),
    .A2(_05070_),
    .B1(net23),
    .C1(net51),
    .D1(_05076_),
    .Y(_05080_));
 sky130_fd_sc_hd__o22ai_4 _15493_ (.A1(_04556_),
    .A2(_05068_),
    .B1(_05077_),
    .B2(_05079_),
    .Y(_05081_));
 sky130_fd_sc_hd__and3_2 _15494_ (.A(_05078_),
    .B(_05080_),
    .C(_05069_),
    .X(_05082_));
 sky130_fd_sc_hd__nand3_2 _15495_ (.A(_05078_),
    .B(_05080_),
    .C(_05069_),
    .Y(_05083_));
 sky130_fd_sc_hd__o32a_1 _15496_ (.A1(_01791_),
    .A2(_02120_),
    .A3(_04185_),
    .B1(_02152_),
    .B2(_01824_),
    .X(_05084_));
 sky130_fd_sc_hd__and3_1 _15497_ (.A(_04743_),
    .B(net51),
    .C(net12),
    .X(_05085_));
 sky130_fd_sc_hd__a31o_1 _15498_ (.A1(_04743_),
    .A2(net51),
    .A3(net12),
    .B1(_04740_),
    .X(_05087_));
 sky130_fd_sc_hd__a21oi_2 _15499_ (.A1(_05081_),
    .A2(_05083_),
    .B1(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__o2bb2ai_1 _15500_ (.A1_N(_05081_),
    .A2_N(_05083_),
    .B1(_05084_),
    .B2(_04742_),
    .Y(_05089_));
 sky130_fd_sc_hd__o21a_1 _15501_ (.A1(_04740_),
    .A2(_05085_),
    .B1(_05081_),
    .X(_05090_));
 sky130_fd_sc_hd__o21ai_4 _15502_ (.A1(_04740_),
    .A2(_05085_),
    .B1(_05081_),
    .Y(_05091_));
 sky130_fd_sc_hd__and3_1 _15503_ (.A(_05081_),
    .B(_05083_),
    .C(_05087_),
    .X(_05092_));
 sky130_fd_sc_hd__o211ai_1 _15504_ (.A1(_04740_),
    .A2(_05085_),
    .B1(_05083_),
    .C1(_05081_),
    .Y(_05093_));
 sky130_fd_sc_hd__o21ai_1 _15505_ (.A1(_05082_),
    .A2(_05091_),
    .B1(_05067_),
    .Y(_05094_));
 sky130_fd_sc_hd__o211a_1 _15506_ (.A1(_05082_),
    .A2(_05091_),
    .B1(_05067_),
    .C1(_05089_),
    .X(_05095_));
 sky130_fd_sc_hd__o211ai_2 _15507_ (.A1(_05082_),
    .A2(_05091_),
    .B1(_05067_),
    .C1(_05089_),
    .Y(_05096_));
 sky130_fd_sc_hd__a21oi_1 _15508_ (.A1(_05089_),
    .A2(_05093_),
    .B1(_05067_),
    .Y(_05098_));
 sky130_fd_sc_hd__o22ai_4 _15509_ (.A1(_04552_),
    .A2(_05066_),
    .B1(_05088_),
    .B2(_05092_),
    .Y(_05099_));
 sky130_fd_sc_hd__o31a_1 _15510_ (.A1(_04188_),
    .A2(_04732_),
    .A3(_04753_),
    .B1(_04752_),
    .X(_05100_));
 sky130_fd_sc_hd__a2bb2o_1 _15511_ (.A1_N(_04733_),
    .A2_N(_04753_),
    .B1(_04750_),
    .B2(_04748_),
    .X(_05101_));
 sky130_fd_sc_hd__o2111ai_4 _15512_ (.A1(_04753_),
    .A2(_04733_),
    .B1(_04752_),
    .C1(_05096_),
    .D1(_05099_),
    .Y(_05102_));
 sky130_fd_sc_hd__a22o_1 _15513_ (.A1(_04752_),
    .A2(_04755_),
    .B1(_05096_),
    .B2(_05099_),
    .X(_05103_));
 sky130_fd_sc_hd__o21ai_2 _15514_ (.A1(_05095_),
    .A2(_05098_),
    .B1(_05100_),
    .Y(_05104_));
 sky130_fd_sc_hd__o211ai_2 _15515_ (.A1(_05088_),
    .A2(_05094_),
    .B1(_05099_),
    .C1(_05101_),
    .Y(_05105_));
 sky130_fd_sc_hd__and3_1 _15516_ (.A(_05103_),
    .B(_05063_),
    .C(_05102_),
    .X(_05106_));
 sky130_fd_sc_hd__nand3_2 _15517_ (.A(_05103_),
    .B(_05063_),
    .C(_05102_),
    .Y(_05107_));
 sky130_fd_sc_hd__nand3_4 _15518_ (.A(_05065_),
    .B(_05104_),
    .C(_05105_),
    .Y(_05109_));
 sky130_fd_sc_hd__nand2_1 _15519_ (.A(net12),
    .B(net52),
    .Y(_05110_));
 sky130_fd_sc_hd__and4_4 _15520_ (.A(net12),
    .B(net1),
    .C(net52),
    .D(net53),
    .X(_05111_));
 sky130_fd_sc_hd__a22oi_4 _15521_ (.A1(net12),
    .A2(net52),
    .B1(net53),
    .B2(net1),
    .Y(_05112_));
 sky130_fd_sc_hd__a21oi_1 _15522_ (.A1(net1),
    .A2(net53),
    .B1(_05110_),
    .Y(_05113_));
 sky130_fd_sc_hd__and3_1 _15523_ (.A(_05110_),
    .B(net53),
    .C(net1),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_1 _15524_ (.A(_05111_),
    .B(_05112_),
    .Y(_05115_));
 sky130_fd_sc_hd__o2bb2ai_1 _15525_ (.A1_N(_05107_),
    .A2_N(_05109_),
    .B1(_05111_),
    .B2(_05112_),
    .Y(_05116_));
 sky130_fd_sc_hd__o211ai_2 _15526_ (.A1(_05113_),
    .A2(_05114_),
    .B1(_05107_),
    .C1(_05109_),
    .Y(_05117_));
 sky130_fd_sc_hd__o2bb2ai_2 _15527_ (.A1_N(_05107_),
    .A2_N(_05109_),
    .B1(_05113_),
    .B2(_05114_),
    .Y(_05118_));
 sky130_fd_sc_hd__o211ai_2 _15528_ (.A1(_05111_),
    .A2(_05112_),
    .B1(_05107_),
    .C1(_05109_),
    .Y(_05120_));
 sky130_fd_sc_hd__a21oi_2 _15529_ (.A1(_04577_),
    .A2(_04582_),
    .B1(_04578_),
    .Y(_05121_));
 sky130_fd_sc_hd__o21ai_2 _15530_ (.A1(_04576_),
    .A2(_04580_),
    .B1(_04579_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand3_1 _15531_ (.A(_05118_),
    .B(_05121_),
    .C(_05120_),
    .Y(_05123_));
 sky130_fd_sc_hd__and3_2 _15532_ (.A(_05116_),
    .B(_05117_),
    .C(_05122_),
    .X(_05124_));
 sky130_fd_sc_hd__nand3_2 _15533_ (.A(_05116_),
    .B(_05117_),
    .C(_05122_),
    .Y(_05125_));
 sky130_fd_sc_hd__a31o_1 _15534_ (.A1(_04772_),
    .A2(net52),
    .A3(net1),
    .B1(_04773_),
    .X(_05126_));
 sky130_fd_sc_hd__a31oi_2 _15535_ (.A1(_04772_),
    .A2(net52),
    .A3(net1),
    .B1(_04773_),
    .Y(_05127_));
 sky130_fd_sc_hd__a21oi_2 _15536_ (.A1(_05123_),
    .A2(_05125_),
    .B1(_05126_),
    .Y(_05128_));
 sky130_fd_sc_hd__a21o_1 _15537_ (.A1(_05123_),
    .A2(_05125_),
    .B1(_05126_),
    .X(_05129_));
 sky130_fd_sc_hd__a31oi_2 _15538_ (.A1(_05118_),
    .A2(_05120_),
    .A3(_05121_),
    .B1(_05127_),
    .Y(_05131_));
 sky130_fd_sc_hd__a31o_2 _15539_ (.A1(_05118_),
    .A2(_05120_),
    .A3(_05121_),
    .B1(_05127_),
    .X(_05132_));
 sky130_fd_sc_hd__and3_1 _15540_ (.A(_05123_),
    .B(_05125_),
    .C(_05126_),
    .X(_05133_));
 sky130_fd_sc_hd__o21ai_1 _15541_ (.A1(_05124_),
    .A2(_05132_),
    .B1(_05129_),
    .Y(_05134_));
 sky130_fd_sc_hd__o211ai_2 _15542_ (.A1(_05128_),
    .A2(_05133_),
    .B1(_05061_),
    .C1(_05062_),
    .Y(_05135_));
 sky130_fd_sc_hd__a21o_1 _15543_ (.A1(_05061_),
    .A2(_05062_),
    .B1(_05134_),
    .X(_05136_));
 sky130_fd_sc_hd__o2bb2ai_2 _15544_ (.A1_N(_05061_),
    .A2_N(_05062_),
    .B1(_05128_),
    .B2(_05133_),
    .Y(_05137_));
 sky130_fd_sc_hd__o211ai_2 _15545_ (.A1(_05124_),
    .A2(_05132_),
    .B1(_05129_),
    .C1(_05061_),
    .Y(_05138_));
 sky130_fd_sc_hd__o2111ai_4 _15546_ (.A1(_05124_),
    .A2(_05132_),
    .B1(_05129_),
    .C1(_05061_),
    .D1(_05062_),
    .Y(_05139_));
 sky130_fd_sc_hd__a22oi_4 _15547_ (.A1(_04731_),
    .A2(_04823_),
    .B1(_05137_),
    .B2(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__nand3_1 _15548_ (.A(_05136_),
    .B(_04824_),
    .C(_05135_),
    .Y(_05142_));
 sky130_fd_sc_hd__a22oi_1 _15549_ (.A1(_04730_),
    .A2(_04798_),
    .B1(_05135_),
    .B2(_05136_),
    .Y(_05143_));
 sky130_fd_sc_hd__nand4_4 _15550_ (.A(_04731_),
    .B(_04823_),
    .C(_05137_),
    .D(_05139_),
    .Y(_05144_));
 sky130_fd_sc_hd__nor2_1 _15551_ (.A(_04216_),
    .B(_04782_),
    .Y(_05145_));
 sky130_fd_sc_hd__a21oi_2 _15552_ (.A1(_04781_),
    .A2(_04216_),
    .B1(_04782_),
    .Y(_05146_));
 sky130_fd_sc_hd__a31oi_1 _15553_ (.A1(_05136_),
    .A2(_04824_),
    .A3(_05135_),
    .B1(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__nand2_1 _15554_ (.A(_05147_),
    .B(_05144_),
    .Y(_05148_));
 sky130_fd_sc_hd__o2bb2ai_1 _15555_ (.A1_N(_05142_),
    .A2_N(_05144_),
    .B1(_05145_),
    .B2(_04780_),
    .Y(_05149_));
 sky130_fd_sc_hd__o22ai_1 _15556_ (.A1(_04782_),
    .A2(_04787_),
    .B1(_05140_),
    .B2(_05143_),
    .Y(_05150_));
 sky130_fd_sc_hd__o2111ai_1 _15557_ (.A1(_04217_),
    .A2(_04780_),
    .B1(_04783_),
    .C1(_05142_),
    .D1(_05144_),
    .Y(_05151_));
 sky130_fd_sc_hd__nand2_1 _15558_ (.A(_05148_),
    .B(_05149_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21oi_1 _15559_ (.A1(_04511_),
    .A2(_04803_),
    .B1(_04800_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand3_1 _15560_ (.A(_05150_),
    .B(_05151_),
    .C(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21ai_1 _15561_ (.A1(_04800_),
    .A2(_04804_),
    .B1(_05149_),
    .Y(_05156_));
 sky130_fd_sc_hd__o211a_1 _15562_ (.A1(_04800_),
    .A2(_04804_),
    .B1(_05148_),
    .C1(_05149_),
    .X(_05157_));
 sky130_fd_sc_hd__o211ai_1 _15563_ (.A1(_04800_),
    .A2(_04804_),
    .B1(_05148_),
    .C1(_05149_),
    .Y(_05158_));
 sky130_fd_sc_hd__o2bb2ai_1 _15564_ (.A1_N(_05155_),
    .A2_N(_05158_),
    .B1(_04509_),
    .B2(_04811_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand3_1 _15565_ (.A(_05155_),
    .B(_04810_),
    .C(_04508_),
    .Y(_05160_));
 sky130_fd_sc_hd__o21a_1 _15566_ (.A1(_05157_),
    .A2(_05160_),
    .B1(_05159_),
    .X(_05161_));
 sky130_fd_sc_hd__a211o_1 _15567_ (.A1(_04499_),
    .A2(_04501_),
    .B1(_04813_),
    .C1(_04815_),
    .X(_05162_));
 sky130_fd_sc_hd__a21oi_1 _15568_ (.A1(_04499_),
    .A2(_04501_),
    .B1(_04817_),
    .Y(_05164_));
 sky130_fd_sc_hd__o31ai_4 _15569_ (.A1(_04503_),
    .A2(_04820_),
    .A3(_04507_),
    .B1(_05162_),
    .Y(_05165_));
 sky130_fd_sc_hd__xor2_1 _15570_ (.A(_05161_),
    .B(_05165_),
    .X(net85));
 sky130_fd_sc_hd__o21ai_1 _15571_ (.A1(_05146_),
    .A2(_05140_),
    .B1(_05144_),
    .Y(_05166_));
 sky130_fd_sc_hd__a31o_1 _15572_ (.A1(_05116_),
    .A2(_05117_),
    .A3(_05122_),
    .B1(_05131_),
    .X(_05167_));
 sky130_fd_sc_hd__inv_2 _15573_ (.A(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__o21ai_2 _15574_ (.A1(_05128_),
    .A2(_05133_),
    .B1(_05062_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_1 _15575_ (.A(_05062_),
    .B(_05138_),
    .Y(_05170_));
 sky130_fd_sc_hd__nand2_1 _15576_ (.A(_05061_),
    .B(_05169_),
    .Y(_05171_));
 sky130_fd_sc_hd__a31oi_4 _15577_ (.A1(_05033_),
    .A2(_05034_),
    .A3(_05037_),
    .B1(_05044_),
    .Y(_05172_));
 sky130_fd_sc_hd__o22ai_2 _15578_ (.A1(_05094_),
    .A2(_05088_),
    .B1(_05100_),
    .B2(_05098_),
    .Y(_05173_));
 sky130_fd_sc_hd__a21oi_2 _15579_ (.A1(_05099_),
    .A2(_05101_),
    .B1(_05095_),
    .Y(_05174_));
 sky130_fd_sc_hd__o41a_1 _15580_ (.A1(_04556_),
    .A2(_05068_),
    .A3(_05077_),
    .A4(_05079_),
    .B1(_05091_),
    .X(_05175_));
 sky130_fd_sc_hd__and3_1 _15581_ (.A(_05076_),
    .B(net51),
    .C(net23),
    .X(_05176_));
 sky130_fd_sc_hd__o32a_2 _15582_ (.A1(_01802_),
    .A2(_02152_),
    .A3(_05074_),
    .B1(_05070_),
    .B2(_04739_),
    .X(_05177_));
 sky130_fd_sc_hd__a21oi_2 _15583_ (.A1(_04557_),
    .A2(_04999_),
    .B1(_04997_),
    .Y(_05178_));
 sky130_fd_sc_hd__o21ai_2 _15584_ (.A1(_04997_),
    .A2(_05002_),
    .B1(_05001_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_2 _15585_ (.A(net28),
    .B(net50),
    .Y(_05180_));
 sky130_fd_sc_hd__and4_2 _15586_ (.A(net28),
    .B(net27),
    .C(net49),
    .D(net50),
    .X(_05181_));
 sky130_fd_sc_hd__nand2_2 _15587_ (.A(net28),
    .B(net49),
    .Y(_05182_));
 sky130_fd_sc_hd__o21a_1 _15588_ (.A1(_01748_),
    .A2(_02120_),
    .B1(_05070_),
    .X(_05184_));
 sky130_fd_sc_hd__a22o_2 _15589_ (.A1(net28),
    .A2(net49),
    .B1(net50),
    .B2(net27),
    .X(_05185_));
 sky130_fd_sc_hd__o2bb2ai_2 _15590_ (.A1_N(_05070_),
    .A2_N(_05182_),
    .B1(_05180_),
    .B2(_05071_),
    .Y(_05186_));
 sky130_fd_sc_hd__o221ai_4 _15591_ (.A1(_01791_),
    .A2(_02152_),
    .B1(_05071_),
    .B2(_05180_),
    .C1(_05185_),
    .Y(_05187_));
 sky130_fd_sc_hd__nand3_2 _15592_ (.A(_05186_),
    .B(net51),
    .C(net26),
    .Y(_05188_));
 sky130_fd_sc_hd__o2111ai_4 _15593_ (.A1(_05071_),
    .A2(_05180_),
    .B1(net26),
    .C1(net51),
    .D1(_05185_),
    .Y(_05189_));
 sky130_fd_sc_hd__o21ai_4 _15594_ (.A1(_01791_),
    .A2(_02152_),
    .B1(_05186_),
    .Y(_05190_));
 sky130_fd_sc_hd__a2bb2oi_4 _15595_ (.A1_N(_05000_),
    .A2_N(_05178_),
    .B1(_05187_),
    .B2(_05188_),
    .Y(_05191_));
 sky130_fd_sc_hd__o211ai_4 _15596_ (.A1(_05000_),
    .A2(_05178_),
    .B1(_05189_),
    .C1(_05190_),
    .Y(_05192_));
 sky130_fd_sc_hd__a21oi_4 _15597_ (.A1(_05189_),
    .A2(_05190_),
    .B1(_05179_),
    .Y(_05193_));
 sky130_fd_sc_hd__nand3b_2 _15598_ (.A_N(_05179_),
    .B(_05187_),
    .C(_05188_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21a_2 _15599_ (.A1(_05072_),
    .A2(_05176_),
    .B1(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__o21ai_1 _15600_ (.A1(_05072_),
    .A2(_05176_),
    .B1(_05195_),
    .Y(_05197_));
 sky130_fd_sc_hd__o21ai_1 _15601_ (.A1(_05191_),
    .A2(_05193_),
    .B1(_05177_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand3_4 _15602_ (.A(_05177_),
    .B(_05192_),
    .C(_05195_),
    .Y(_05199_));
 sky130_fd_sc_hd__o22ai_4 _15603_ (.A1(_05072_),
    .A2(_05176_),
    .B1(_05191_),
    .B2(_05193_),
    .Y(_05200_));
 sky130_fd_sc_hd__a2bb2oi_4 _15604_ (.A1_N(_05021_),
    .A2_N(_05026_),
    .B1(_05199_),
    .B2(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__o221ai_4 _15605_ (.A1(_05191_),
    .A2(_05197_),
    .B1(_05021_),
    .B2(_05026_),
    .C1(_05198_),
    .Y(_05202_));
 sky130_fd_sc_hd__o2111a_1 _15606_ (.A1(_05008_),
    .A2(_05019_),
    .B1(_05027_),
    .C1(_05199_),
    .D1(_05200_),
    .X(_05203_));
 sky130_fd_sc_hd__o2111ai_4 _15607_ (.A1(_05008_),
    .A2(_05019_),
    .B1(_05027_),
    .C1(_05199_),
    .D1(_05200_),
    .Y(_05204_));
 sky130_fd_sc_hd__o21a_1 _15608_ (.A1(_05082_),
    .A2(_05090_),
    .B1(_05204_),
    .X(_05206_));
 sky130_fd_sc_hd__o211ai_2 _15609_ (.A1(_05082_),
    .A2(_05090_),
    .B1(_05202_),
    .C1(_05204_),
    .Y(_05207_));
 sky130_fd_sc_hd__o21ai_2 _15610_ (.A1(_05201_),
    .A2(_05203_),
    .B1(_05175_),
    .Y(_05208_));
 sky130_fd_sc_hd__o22ai_4 _15611_ (.A1(_05082_),
    .A2(_05090_),
    .B1(_05201_),
    .B2(_05203_),
    .Y(_05209_));
 sky130_fd_sc_hd__nand4_2 _15612_ (.A(_05083_),
    .B(_05091_),
    .C(_05202_),
    .D(_05204_),
    .Y(_05210_));
 sky130_fd_sc_hd__nand3_4 _15613_ (.A(_05174_),
    .B(_05209_),
    .C(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__and3_2 _15614_ (.A(_05208_),
    .B(_05173_),
    .C(_05207_),
    .X(_05212_));
 sky130_fd_sc_hd__nand3_4 _15615_ (.A(_05208_),
    .B(_05173_),
    .C(_05207_),
    .Y(_05213_));
 sky130_fd_sc_hd__and4_1 _15616_ (.A(net23),
    .B(net12),
    .C(net52),
    .D(net53),
    .X(_05214_));
 sky130_fd_sc_hd__nand4_4 _15617_ (.A(net23),
    .B(net12),
    .C(net52),
    .D(net53),
    .Y(_05215_));
 sky130_fd_sc_hd__a22oi_1 _15618_ (.A1(net23),
    .A2(net52),
    .B1(net53),
    .B2(net12),
    .Y(_05217_));
 sky130_fd_sc_hd__or4bb_4 _15619_ (.A(_05217_),
    .B(_02207_),
    .C_N(net1),
    .D_N(_05215_),
    .X(_05218_));
 sky130_fd_sc_hd__a2bb2o_1 _15620_ (.A1_N(_05214_),
    .A2_N(_05217_),
    .B1(net1),
    .B2(net54),
    .X(_05219_));
 sky130_fd_sc_hd__and2_2 _15621_ (.A(_05218_),
    .B(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__nand2_1 _15622_ (.A(_05111_),
    .B(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__inv_2 _15623_ (.A(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__a21oi_2 _15624_ (.A1(_05218_),
    .A2(_05219_),
    .B1(_05111_),
    .Y(_05223_));
 sky130_fd_sc_hd__a41o_1 _15625_ (.A1(net12),
    .A2(net1),
    .A3(net52),
    .A4(net53),
    .B1(_05220_),
    .X(_05224_));
 sky130_fd_sc_hd__and4bb_1 _15626_ (.A_N(_05220_),
    .B_N(_05110_),
    .C(net53),
    .D(net1),
    .X(_05225_));
 sky130_fd_sc_hd__and3b_1 _15627_ (.A_N(_05111_),
    .B(_05218_),
    .C(_05219_),
    .X(_05226_));
 sky130_fd_sc_hd__nand2_1 _15628_ (.A(_05221_),
    .B(_05224_),
    .Y(_05228_));
 sky130_fd_sc_hd__o211ai_4 _15629_ (.A1(_05222_),
    .A2(_05223_),
    .B1(_05211_),
    .C1(_05213_),
    .Y(_05229_));
 sky130_fd_sc_hd__o2bb2ai_2 _15630_ (.A1_N(_05211_),
    .A2_N(_05213_),
    .B1(_05225_),
    .B2(_05226_),
    .Y(_05230_));
 sky130_fd_sc_hd__o2bb2ai_2 _15631_ (.A1_N(_05211_),
    .A2_N(_05213_),
    .B1(_05222_),
    .B2(_05223_),
    .Y(_05231_));
 sky130_fd_sc_hd__a31o_1 _15632_ (.A1(_05174_),
    .A2(_05209_),
    .A3(_05210_),
    .B1(_05228_),
    .X(_05232_));
 sky130_fd_sc_hd__o211a_1 _15633_ (.A1(_05039_),
    .A2(_05172_),
    .B1(_05229_),
    .C1(_05230_),
    .X(_05233_));
 sky130_fd_sc_hd__o211ai_4 _15634_ (.A1(_05039_),
    .A2(_05172_),
    .B1(_05229_),
    .C1(_05230_),
    .Y(_05234_));
 sky130_fd_sc_hd__o221a_1 _15635_ (.A1(_05041_),
    .A2(_05048_),
    .B1(_05212_),
    .B2(_05232_),
    .C1(_05231_),
    .X(_05235_));
 sky130_fd_sc_hd__o221ai_4 _15636_ (.A1(_05041_),
    .A2(_05048_),
    .B1(_05212_),
    .B2(_05232_),
    .C1(_05231_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_1 _15637_ (.A(_05234_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__o21a_1 _15638_ (.A1(_05111_),
    .A2(_05112_),
    .B1(_05109_),
    .X(_05239_));
 sky130_fd_sc_hd__a31o_1 _15639_ (.A1(_05063_),
    .A2(_05102_),
    .A3(_05103_),
    .B1(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__a32o_1 _15640_ (.A1(_05065_),
    .A2(_05104_),
    .A3(_05105_),
    .B1(_05107_),
    .B2(_05115_),
    .X(_05241_));
 sky130_fd_sc_hd__a21oi_2 _15641_ (.A1(_05234_),
    .A2(_05236_),
    .B1(_05240_),
    .Y(_05242_));
 sky130_fd_sc_hd__o21ai_1 _15642_ (.A1(_05106_),
    .A2(_05239_),
    .B1(_05236_),
    .Y(_05243_));
 sky130_fd_sc_hd__and3_1 _15643_ (.A(_05240_),
    .B(_05236_),
    .C(_05234_),
    .X(_05244_));
 sky130_fd_sc_hd__o311a_1 _15644_ (.A1(_05106_),
    .A2(_05111_),
    .A3(_05112_),
    .B1(_05237_),
    .C1(_05109_),
    .X(_05245_));
 sky130_fd_sc_hd__o2bb2ai_1 _15645_ (.A1_N(_05234_),
    .A2_N(_05236_),
    .B1(_05239_),
    .B2(_05106_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand2_1 _15646_ (.A(_05234_),
    .B(_05241_),
    .Y(_05247_));
 sky130_fd_sc_hd__and3_1 _15647_ (.A(_05234_),
    .B(_05236_),
    .C(_05241_),
    .X(_05248_));
 sky130_fd_sc_hd__o21ai_1 _15648_ (.A1(_05235_),
    .A2(_05247_),
    .B1(_05246_),
    .Y(_05250_));
 sky130_fd_sc_hd__o2bb2ai_2 _15649_ (.A1_N(_05237_),
    .A2_N(_05241_),
    .B1(_05243_),
    .B2(_05233_),
    .Y(_05251_));
 sky130_fd_sc_hd__o21ai_1 _15650_ (.A1(_05046_),
    .A2(_05050_),
    .B1(_04968_),
    .Y(_05252_));
 sky130_fd_sc_hd__a32oi_4 _15651_ (.A1(_04827_),
    .A2(_04959_),
    .A3(_04961_),
    .B1(_04966_),
    .B2(_05054_),
    .Y(_05253_));
 sky130_fd_sc_hd__o32ai_4 _15652_ (.A1(_04826_),
    .A2(_04958_),
    .A3(_04960_),
    .B1(_05055_),
    .B2(_04964_),
    .Y(_05254_));
 sky130_fd_sc_hd__o21ai_1 _15653_ (.A1(_04950_),
    .A2(_04955_),
    .B1(_04912_),
    .Y(_05255_));
 sky130_fd_sc_hd__a32oi_4 _15654_ (.A1(_04906_),
    .A2(_04907_),
    .A3(_04909_),
    .B1(_04912_),
    .B2(_04957_),
    .Y(_05256_));
 sky130_fd_sc_hd__a21boi_1 _15655_ (.A1(_04956_),
    .A2(_04911_),
    .B1_N(_04912_),
    .Y(_05257_));
 sky130_fd_sc_hd__o21ai_1 _15656_ (.A1(_04848_),
    .A2(_04851_),
    .B1(_04902_),
    .Y(_05258_));
 sky130_fd_sc_hd__o21ai_2 _15657_ (.A1(_04895_),
    .A2(_04898_),
    .B1(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__a31o_1 _15658_ (.A1(_04849_),
    .A2(_04852_),
    .A3(_04900_),
    .B1(_04901_),
    .X(_05261_));
 sky130_fd_sc_hd__o21a_1 _15659_ (.A1(_01835_),
    .A2(_02098_),
    .B1(_04879_),
    .X(_05262_));
 sky130_fd_sc_hd__o21ai_2 _15660_ (.A1(_04874_),
    .A2(_04875_),
    .B1(_04879_),
    .Y(_05263_));
 sky130_fd_sc_hd__o31a_1 _15661_ (.A1(_01835_),
    .A2(_02098_),
    .A3(_04875_),
    .B1(_04879_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_2 _15662_ (.A(net61),
    .B(net16),
    .Y(_05265_));
 sky130_fd_sc_hd__and4_1 _15663_ (.A(net61),
    .B(net62),
    .C(net15),
    .D(net16),
    .X(_05266_));
 sky130_fd_sc_hd__nand4_1 _15664_ (.A(net61),
    .B(net62),
    .C(net15),
    .D(net16),
    .Y(_05267_));
 sky130_fd_sc_hd__a22oi_4 _15665_ (.A1(net62),
    .A2(net15),
    .B1(net16),
    .B2(net61),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _15666_ (.A(_04831_),
    .B(_05265_),
    .Y(_05269_));
 sky130_fd_sc_hd__a2bb2oi_1 _15667_ (.A1_N(_01890_),
    .A2_N(_02065_),
    .B1(_05267_),
    .B2(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__o22ai_4 _15668_ (.A1(_01890_),
    .A2(_02065_),
    .B1(_05266_),
    .B2(_05268_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand3_2 _15669_ (.A(_05267_),
    .B(net14),
    .C(net63),
    .Y(_05273_));
 sky130_fd_sc_hd__a21oi_1 _15670_ (.A1(_04831_),
    .A2(_05265_),
    .B1(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__o21ai_2 _15671_ (.A1(_05268_),
    .A2(_05273_),
    .B1(_05272_),
    .Y(_05275_));
 sky130_fd_sc_hd__o22ai_4 _15672_ (.A1(_04875_),
    .A2(_05262_),
    .B1(_05270_),
    .B2(_05274_),
    .Y(_05276_));
 sky130_fd_sc_hd__o211a_2 _15673_ (.A1(_05268_),
    .A2(_05273_),
    .B1(_05263_),
    .C1(_05272_),
    .X(_05277_));
 sky130_fd_sc_hd__o211ai_4 _15674_ (.A1(_05268_),
    .A2(_05273_),
    .B1(_05263_),
    .C1(_05272_),
    .Y(_05278_));
 sky130_fd_sc_hd__o21a_1 _15675_ (.A1(_01890_),
    .A2(_02043_),
    .B1(_04834_),
    .X(_05279_));
 sky130_fd_sc_hd__or2_1 _15676_ (.A(_04830_),
    .B(_04835_),
    .X(_05280_));
 sky130_fd_sc_hd__a31o_1 _15677_ (.A1(_04836_),
    .A2(net13),
    .A3(net63),
    .B1(_04832_),
    .X(_05281_));
 sky130_fd_sc_hd__a21oi_1 _15678_ (.A1(_05276_),
    .A2(_05278_),
    .B1(_05281_),
    .Y(_05283_));
 sky130_fd_sc_hd__o2bb2ai_2 _15679_ (.A1_N(_05276_),
    .A2_N(_05278_),
    .B1(_05279_),
    .B2(_04835_),
    .Y(_05284_));
 sky130_fd_sc_hd__a22oi_4 _15680_ (.A1(_04834_),
    .A2(_05280_),
    .B1(_05275_),
    .B2(_05264_),
    .Y(_05285_));
 sky130_fd_sc_hd__nand2_1 _15681_ (.A(_05276_),
    .B(_05281_),
    .Y(_05286_));
 sky130_fd_sc_hd__o21ai_1 _15682_ (.A1(_05264_),
    .A2(_05275_),
    .B1(_05285_),
    .Y(_05287_));
 sky130_fd_sc_hd__a21oi_1 _15683_ (.A1(_05278_),
    .A2(_05285_),
    .B1(_05283_),
    .Y(_05288_));
 sky130_fd_sc_hd__o21ai_2 _15684_ (.A1(_05277_),
    .A2(_05286_),
    .B1(_05284_),
    .Y(_05289_));
 sky130_fd_sc_hd__o21ai_2 _15685_ (.A1(_04858_),
    .A2(_04859_),
    .B1(_04862_),
    .Y(_05290_));
 sky130_fd_sc_hd__o21a_1 _15686_ (.A1(_04858_),
    .A2(_04859_),
    .B1(_04862_),
    .X(_05291_));
 sky130_fd_sc_hd__nand2_1 _15687_ (.A(net55),
    .B(net20),
    .Y(_05292_));
 sky130_fd_sc_hd__nand2_2 _15688_ (.A(net33),
    .B(net22),
    .Y(_05294_));
 sky130_fd_sc_hd__a22oi_4 _15689_ (.A1(net44),
    .A2(net21),
    .B1(net22),
    .B2(net33),
    .Y(_05295_));
 sky130_fd_sc_hd__a22o_1 _15690_ (.A1(net44),
    .A2(net21),
    .B1(net22),
    .B2(net33),
    .X(_05296_));
 sky130_fd_sc_hd__and4_2 _15691_ (.A(net33),
    .B(net44),
    .C(net21),
    .D(net22),
    .X(_05297_));
 sky130_fd_sc_hd__nand4_2 _15692_ (.A(net33),
    .B(net44),
    .C(net21),
    .D(net22),
    .Y(_05298_));
 sky130_fd_sc_hd__o211ai_2 _15693_ (.A1(_01780_),
    .A2(_02163_),
    .B1(_05296_),
    .C1(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__o21bai_1 _15694_ (.A1(_05295_),
    .A2(_05297_),
    .B1_N(_05292_),
    .Y(_05300_));
 sky130_fd_sc_hd__o22a_4 _15695_ (.A1(_01780_),
    .A2(_02163_),
    .B1(_05295_),
    .B2(_05297_),
    .X(_05301_));
 sky130_fd_sc_hd__a22o_1 _15696_ (.A1(net55),
    .A2(net20),
    .B1(_05296_),
    .B2(_05298_),
    .X(_05302_));
 sky130_fd_sc_hd__nand4_2 _15697_ (.A(_05296_),
    .B(_05298_),
    .C(net55),
    .D(net20),
    .Y(_05303_));
 sky130_fd_sc_hd__nand3_4 _15698_ (.A(_05291_),
    .B(_05299_),
    .C(_05300_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_4 _15699_ (.A(_05290_),
    .B(_05303_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand3_2 _15700_ (.A(_05302_),
    .B(_05303_),
    .C(_05290_),
    .Y(_05307_));
 sky130_fd_sc_hd__o21ai_1 _15701_ (.A1(_05301_),
    .A2(_05306_),
    .B1(_05305_),
    .Y(_05308_));
 sky130_fd_sc_hd__nand2_1 _15702_ (.A(net60),
    .B(net17),
    .Y(_05309_));
 sky130_fd_sc_hd__a22oi_2 _15703_ (.A1(net59),
    .A2(net18),
    .B1(net19),
    .B2(net58),
    .Y(_05310_));
 sky130_fd_sc_hd__a22o_1 _15704_ (.A1(net59),
    .A2(net18),
    .B1(net19),
    .B2(net58),
    .X(_05311_));
 sky130_fd_sc_hd__and4_1 _15705_ (.A(net58),
    .B(net59),
    .C(net18),
    .D(net19),
    .X(_05312_));
 sky130_fd_sc_hd__nand4_2 _15706_ (.A(net58),
    .B(net59),
    .C(net18),
    .D(net19),
    .Y(_05313_));
 sky130_fd_sc_hd__and3_2 _15707_ (.A(_05309_),
    .B(_05311_),
    .C(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__nand3_1 _15708_ (.A(_05309_),
    .B(_05311_),
    .C(_05313_),
    .Y(_05316_));
 sky130_fd_sc_hd__o211a_2 _15709_ (.A1(_05310_),
    .A2(_05312_),
    .B1(net60),
    .C1(net17),
    .X(_05317_));
 sky130_fd_sc_hd__o21bai_1 _15710_ (.A1(_05310_),
    .A2(_05312_),
    .B1_N(_05309_),
    .Y(_05318_));
 sky130_fd_sc_hd__o2bb2a_1 _15711_ (.A1_N(net60),
    .A2_N(net17),
    .B1(_05310_),
    .B2(_05312_),
    .X(_05319_));
 sky130_fd_sc_hd__and4_1 _15712_ (.A(_05311_),
    .B(_05313_),
    .C(net60),
    .D(net17),
    .X(_05320_));
 sky130_fd_sc_hd__nor2_1 _15713_ (.A(_05314_),
    .B(_05317_),
    .Y(_05321_));
 sky130_fd_sc_hd__nand2_1 _15714_ (.A(_05316_),
    .B(_05318_),
    .Y(_05322_));
 sky130_fd_sc_hd__o21ai_1 _15715_ (.A1(_05314_),
    .A2(_05317_),
    .B1(_05305_),
    .Y(_05323_));
 sky130_fd_sc_hd__o221a_2 _15716_ (.A1(_05314_),
    .A2(_05317_),
    .B1(_05301_),
    .B2(_05306_),
    .C1(_05305_),
    .X(_05324_));
 sky130_fd_sc_hd__o221ai_4 _15717_ (.A1(_05314_),
    .A2(_05317_),
    .B1(_05301_),
    .B2(_05306_),
    .C1(_05305_),
    .Y(_05325_));
 sky130_fd_sc_hd__o2bb2ai_1 _15718_ (.A1_N(_05305_),
    .A2_N(_05307_),
    .B1(_05319_),
    .B2(_05320_),
    .Y(_05327_));
 sky130_fd_sc_hd__o221ai_4 _15719_ (.A1(_05301_),
    .A2(_05306_),
    .B1(_05319_),
    .B2(_05320_),
    .C1(_05305_),
    .Y(_05328_));
 sky130_fd_sc_hd__o2bb2ai_2 _15720_ (.A1_N(_05305_),
    .A2_N(_05307_),
    .B1(_05314_),
    .B2(_05317_),
    .Y(_05329_));
 sky130_fd_sc_hd__a32oi_2 _15721_ (.A1(_04857_),
    .A2(_04863_),
    .A3(_04864_),
    .B1(_04881_),
    .B2(_04883_),
    .Y(_05330_));
 sky130_fd_sc_hd__a21oi_2 _15722_ (.A1(_04870_),
    .A2(_04890_),
    .B1(_04872_),
    .Y(_05331_));
 sky130_fd_sc_hd__o22ai_2 _15723_ (.A1(_04865_),
    .A2(_04871_),
    .B1(_04889_),
    .B2(_04869_),
    .Y(_05332_));
 sky130_fd_sc_hd__nand3_4 _15724_ (.A(_05331_),
    .B(_05329_),
    .C(_05328_),
    .Y(_05333_));
 sky130_fd_sc_hd__o2bb2ai_2 _15725_ (.A1_N(_05321_),
    .A2_N(_05308_),
    .B1(_04872_),
    .B2(_05330_),
    .Y(_05334_));
 sky130_fd_sc_hd__nand3_4 _15726_ (.A(_05325_),
    .B(_05327_),
    .C(_05332_),
    .Y(_05335_));
 sky130_fd_sc_hd__o2111ai_4 _15727_ (.A1(_05286_),
    .A2(_05277_),
    .B1(_05284_),
    .C1(_05333_),
    .D1(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__a22o_2 _15728_ (.A1(_05284_),
    .A2(_05287_),
    .B1(_05333_),
    .B2(_05335_),
    .X(_05338_));
 sky130_fd_sc_hd__o211ai_2 _15729_ (.A1(_05324_),
    .A2(_05334_),
    .B1(_05333_),
    .C1(_05289_),
    .Y(_05339_));
 sky130_fd_sc_hd__a21o_1 _15730_ (.A1(_05333_),
    .A2(_05335_),
    .B1(_05289_),
    .X(_05340_));
 sky130_fd_sc_hd__o211ai_4 _15731_ (.A1(_04901_),
    .A2(_04904_),
    .B1(_05336_),
    .C1(_05338_),
    .Y(_05341_));
 sky130_fd_sc_hd__and3_1 _15732_ (.A(_05340_),
    .B(_05259_),
    .C(_05339_),
    .X(_05342_));
 sky130_fd_sc_hd__nand3_4 _15733_ (.A(_05340_),
    .B(_05259_),
    .C(_05339_),
    .Y(_05343_));
 sky130_fd_sc_hd__a21boi_2 _15734_ (.A1(_04841_),
    .A2(_04847_),
    .B1_N(_04845_),
    .Y(_05344_));
 sky130_fd_sc_hd__o21ai_4 _15735_ (.A1(_04839_),
    .A2(_04842_),
    .B1(_04850_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(net38),
    .B(net7),
    .Y(_05346_));
 sky130_fd_sc_hd__a22oi_4 _15737_ (.A1(net37),
    .A2(net8),
    .B1(net9),
    .B2(net36),
    .Y(_05347_));
 sky130_fd_sc_hd__and4_2 _15738_ (.A(net36),
    .B(net37),
    .C(net8),
    .D(net9),
    .X(_05349_));
 sky130_fd_sc_hd__nand4_1 _15739_ (.A(net36),
    .B(net37),
    .C(net8),
    .D(net9),
    .Y(_05350_));
 sky130_fd_sc_hd__a211o_2 _15740_ (.A1(net38),
    .A2(net7),
    .B1(_05347_),
    .C1(_05349_),
    .X(_05351_));
 sky130_fd_sc_hd__o211ai_4 _15741_ (.A1(_05347_),
    .A2(_05349_),
    .B1(net38),
    .C1(net7),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_2 _15742_ (.A(_05351_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__o2bb2ai_1 _15743_ (.A1_N(_04916_),
    .A2_N(_04919_),
    .B1(_04917_),
    .B2(_04673_),
    .Y(_05354_));
 sky130_fd_sc_hd__a21boi_2 _15744_ (.A1(_04919_),
    .A2(_04916_),
    .B1_N(_04918_),
    .Y(_05355_));
 sky130_fd_sc_hd__nand2_2 _15745_ (.A(net35),
    .B(net10),
    .Y(_05356_));
 sky130_fd_sc_hd__a22oi_4 _15746_ (.A1(net34),
    .A2(net11),
    .B1(net13),
    .B2(net64),
    .Y(_05357_));
 sky130_fd_sc_hd__a22o_1 _15747_ (.A1(net34),
    .A2(net11),
    .B1(net13),
    .B2(net64),
    .X(_05358_));
 sky130_fd_sc_hd__and4_1 _15748_ (.A(net64),
    .B(net34),
    .C(net11),
    .D(net13),
    .X(_05360_));
 sky130_fd_sc_hd__nand4_2 _15749_ (.A(net64),
    .B(net34),
    .C(net11),
    .D(net13),
    .Y(_05361_));
 sky130_fd_sc_hd__o211ai_2 _15750_ (.A1(_01934_),
    .A2(_02021_),
    .B1(_05358_),
    .C1(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__o21bai_2 _15751_ (.A1(_05357_),
    .A2(_05360_),
    .B1_N(_05356_),
    .Y(_05363_));
 sky130_fd_sc_hd__a41o_1 _15752_ (.A1(net64),
    .A2(net34),
    .A3(net11),
    .A4(net13),
    .B1(_05356_),
    .X(_05364_));
 sky130_fd_sc_hd__o21ai_1 _15753_ (.A1(_05357_),
    .A2(_05360_),
    .B1(_05356_),
    .Y(_05365_));
 sky130_fd_sc_hd__o211ai_4 _15754_ (.A1(_05357_),
    .A2(_05364_),
    .B1(_05354_),
    .C1(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__inv_2 _15755_ (.A(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand3_4 _15756_ (.A(_05355_),
    .B(_05362_),
    .C(_05363_),
    .Y(_05368_));
 sky130_fd_sc_hd__a22o_2 _15757_ (.A1(_05351_),
    .A2(_05352_),
    .B1(_05366_),
    .B2(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__nand4_4 _15758_ (.A(_05351_),
    .B(_05352_),
    .C(_05366_),
    .D(_05368_),
    .Y(_05371_));
 sky130_fd_sc_hd__a32o_1 _15759_ (.A1(_05355_),
    .A2(_05362_),
    .A3(_05363_),
    .B1(_05352_),
    .B2(_05351_),
    .X(_05372_));
 sky130_fd_sc_hd__nand3_2 _15760_ (.A(_05353_),
    .B(_05366_),
    .C(_05368_),
    .Y(_05373_));
 sky130_fd_sc_hd__a21o_2 _15761_ (.A1(_05366_),
    .A2(_05368_),
    .B1(_05353_),
    .X(_05374_));
 sky130_fd_sc_hd__o211a_1 _15762_ (.A1(_05367_),
    .A2(_05372_),
    .B1(_05374_),
    .C1(_05345_),
    .X(_05375_));
 sky130_fd_sc_hd__o211ai_4 _15763_ (.A1(_05367_),
    .A2(_05372_),
    .B1(_05374_),
    .C1(_05345_),
    .Y(_05376_));
 sky130_fd_sc_hd__and3_2 _15764_ (.A(_05344_),
    .B(_05369_),
    .C(_05371_),
    .X(_05377_));
 sky130_fd_sc_hd__nand4_4 _15765_ (.A(_04845_),
    .B(_04852_),
    .C(_05369_),
    .D(_05371_),
    .Y(_05378_));
 sky130_fd_sc_hd__a32oi_4 _15766_ (.A1(_04915_),
    .A2(_04922_),
    .A3(_04924_),
    .B1(_04925_),
    .B2(_04938_),
    .Y(_05379_));
 sky130_fd_sc_hd__a32o_2 _15767_ (.A1(_04915_),
    .A2(_04922_),
    .A3(_04924_),
    .B1(_04925_),
    .B2(_04938_),
    .X(_05380_));
 sky130_fd_sc_hd__and3_1 _15768_ (.A(_05376_),
    .B(_05378_),
    .C(_05379_),
    .X(_05382_));
 sky130_fd_sc_hd__a21oi_1 _15769_ (.A1(_05376_),
    .A2(_05378_),
    .B1(_05379_),
    .Y(_05383_));
 sky130_fd_sc_hd__a21oi_4 _15770_ (.A1(_05376_),
    .A2(_05378_),
    .B1(_05380_),
    .Y(_05384_));
 sky130_fd_sc_hd__a21o_1 _15771_ (.A1(_05376_),
    .A2(_05378_),
    .B1(_05380_),
    .X(_05385_));
 sky130_fd_sc_hd__a31oi_4 _15772_ (.A1(_05344_),
    .A2(_05369_),
    .A3(_05371_),
    .B1(_05379_),
    .Y(_05386_));
 sky130_fd_sc_hd__and3_2 _15773_ (.A(_05376_),
    .B(_05378_),
    .C(_05380_),
    .X(_05387_));
 sky130_fd_sc_hd__nand2_2 _15774_ (.A(_05386_),
    .B(_05376_),
    .Y(_05388_));
 sky130_fd_sc_hd__o2bb2ai_1 _15775_ (.A1_N(_05341_),
    .A2_N(_05343_),
    .B1(_05382_),
    .B2(_05383_),
    .Y(_05389_));
 sky130_fd_sc_hd__o211ai_2 _15776_ (.A1(_05384_),
    .A2(_05387_),
    .B1(_05341_),
    .C1(_05343_),
    .Y(_05390_));
 sky130_fd_sc_hd__o2bb2ai_4 _15777_ (.A1_N(_05341_),
    .A2_N(_05343_),
    .B1(_05384_),
    .B2(_05387_),
    .Y(_05391_));
 sky130_fd_sc_hd__o211a_1 _15778_ (.A1(_05382_),
    .A2(_05383_),
    .B1(_05341_),
    .C1(_05343_),
    .X(_05393_));
 sky130_fd_sc_hd__nand4_4 _15779_ (.A(_05341_),
    .B(_05343_),
    .C(_05385_),
    .D(_05388_),
    .Y(_05394_));
 sky130_fd_sc_hd__a22oi_4 _15780_ (.A1(_04911_),
    .A2(_05255_),
    .B1(_05391_),
    .B2(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand3_4 _15781_ (.A(_05257_),
    .B(_05389_),
    .C(_05390_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand2_1 _15782_ (.A(_05256_),
    .B(_05391_),
    .Y(_05397_));
 sky130_fd_sc_hd__and3_1 _15783_ (.A(_05256_),
    .B(_05391_),
    .C(_05394_),
    .X(_05398_));
 sky130_fd_sc_hd__nand3_4 _15784_ (.A(_05256_),
    .B(_05391_),
    .C(_05394_),
    .Y(_05399_));
 sky130_fd_sc_hd__o21ai_4 _15785_ (.A1(_04974_),
    .A2(_04985_),
    .B1(_04990_),
    .Y(_05400_));
 sky130_fd_sc_hd__o21ai_1 _15786_ (.A1(_04927_),
    .A2(_04928_),
    .B1(_04930_),
    .Y(_05401_));
 sky130_fd_sc_hd__o21a_1 _15787_ (.A1(_04927_),
    .A2(_04928_),
    .B1(_04930_),
    .X(_05402_));
 sky130_fd_sc_hd__nand2_1 _15788_ (.A(net4),
    .B(net41),
    .Y(_05404_));
 sky130_fd_sc_hd__a22oi_4 _15789_ (.A1(net6),
    .A2(net39),
    .B1(net40),
    .B2(net5),
    .Y(_05405_));
 sky130_fd_sc_hd__a22o_1 _15790_ (.A1(net6),
    .A2(net39),
    .B1(net40),
    .B2(net5),
    .X(_05406_));
 sky130_fd_sc_hd__and4_2 _15791_ (.A(net5),
    .B(net6),
    .C(net39),
    .D(net40),
    .X(_05407_));
 sky130_fd_sc_hd__nand4_4 _15792_ (.A(net5),
    .B(net6),
    .C(net39),
    .D(net40),
    .Y(_05408_));
 sky130_fd_sc_hd__o211ai_4 _15793_ (.A1(_01945_),
    .A2(_02010_),
    .B1(_05406_),
    .C1(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__o21bai_2 _15794_ (.A1(_05405_),
    .A2(_05407_),
    .B1_N(_05404_),
    .Y(_05410_));
 sky130_fd_sc_hd__o21ai_1 _15795_ (.A1(_05405_),
    .A2(_05407_),
    .B1(_05404_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand4_1 _15796_ (.A(_05406_),
    .B(_05408_),
    .C(net4),
    .D(net41),
    .Y(_05412_));
 sky130_fd_sc_hd__nand3_2 _15797_ (.A(_05402_),
    .B(_05409_),
    .C(_05410_),
    .Y(_05413_));
 sky130_fd_sc_hd__and3_2 _15798_ (.A(_05411_),
    .B(_05412_),
    .C(_05401_),
    .X(_05415_));
 sky130_fd_sc_hd__nand3_2 _15799_ (.A(_05411_),
    .B(_05412_),
    .C(_05401_),
    .Y(_05416_));
 sky130_fd_sc_hd__o21a_1 _15800_ (.A1(_01923_),
    .A2(_02010_),
    .B1(_04980_),
    .X(_05417_));
 sky130_fd_sc_hd__a31o_1 _15801_ (.A1(_04978_),
    .A2(net41),
    .A3(net3),
    .B1(_04979_),
    .X(_05418_));
 sky130_fd_sc_hd__o31a_1 _15802_ (.A1(_01923_),
    .A2(_02010_),
    .A3(_04977_),
    .B1(_04980_),
    .X(_05419_));
 sky130_fd_sc_hd__o2bb2ai_4 _15803_ (.A1_N(_05413_),
    .A2_N(_05416_),
    .B1(_05417_),
    .B2(_04977_),
    .Y(_05420_));
 sky130_fd_sc_hd__a31oi_4 _15804_ (.A1(_05402_),
    .A2(_05409_),
    .A3(_05410_),
    .B1(_05419_),
    .Y(_05421_));
 sky130_fd_sc_hd__a31o_1 _15805_ (.A1(_05402_),
    .A2(_05409_),
    .A3(_05410_),
    .B1(_05419_),
    .X(_05422_));
 sky130_fd_sc_hd__nand3_2 _15806_ (.A(_05413_),
    .B(_05416_),
    .C(_05418_),
    .Y(_05423_));
 sky130_fd_sc_hd__a21oi_4 _15807_ (.A1(_05420_),
    .A2(_05423_),
    .B1(_05400_),
    .Y(_05424_));
 sky130_fd_sc_hd__a21o_1 _15808_ (.A1(_05420_),
    .A2(_05423_),
    .B1(_05400_),
    .X(_05426_));
 sky130_fd_sc_hd__o211a_2 _15809_ (.A1(_05415_),
    .A2(_05422_),
    .B1(_05420_),
    .C1(_05400_),
    .X(_05427_));
 sky130_fd_sc_hd__o211ai_4 _15810_ (.A1(_05415_),
    .A2(_05422_),
    .B1(_05420_),
    .C1(_05400_),
    .Y(_05428_));
 sky130_fd_sc_hd__o21ai_1 _15811_ (.A1(_01879_),
    .A2(_02054_),
    .B1(_05012_),
    .Y(_05429_));
 sky130_fd_sc_hd__o21a_1 _15812_ (.A1(_05010_),
    .A2(_05013_),
    .B1(_05012_),
    .X(_05430_));
 sky130_fd_sc_hd__nand2_1 _15813_ (.A(net32),
    .B(net45),
    .Y(_05431_));
 sky130_fd_sc_hd__nand2_1 _15814_ (.A(net3),
    .B(net42),
    .Y(_05432_));
 sky130_fd_sc_hd__a22oi_4 _15815_ (.A1(net3),
    .A2(net42),
    .B1(net43),
    .B2(net2),
    .Y(_05433_));
 sky130_fd_sc_hd__a22o_1 _15816_ (.A1(net3),
    .A2(net42),
    .B1(net43),
    .B2(net2),
    .X(_05434_));
 sky130_fd_sc_hd__and4_1 _15817_ (.A(net2),
    .B(net3),
    .C(net42),
    .D(net43),
    .X(_05435_));
 sky130_fd_sc_hd__nand4_2 _15818_ (.A(net2),
    .B(net3),
    .C(net42),
    .D(net43),
    .Y(_05437_));
 sky130_fd_sc_hd__o211ai_1 _15819_ (.A1(_01912_),
    .A2(_02054_),
    .B1(_05434_),
    .C1(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__o21bai_1 _15820_ (.A1(_05433_),
    .A2(_05435_),
    .B1_N(_05431_),
    .Y(_05439_));
 sky130_fd_sc_hd__o22a_2 _15821_ (.A1(_01912_),
    .A2(_02054_),
    .B1(_05433_),
    .B2(_05435_),
    .X(_05440_));
 sky130_fd_sc_hd__a41o_1 _15822_ (.A1(net2),
    .A2(net3),
    .A3(net42),
    .A4(net43),
    .B1(_05431_),
    .X(_05441_));
 sky130_fd_sc_hd__nand3_2 _15823_ (.A(_05430_),
    .B(_05438_),
    .C(_05439_),
    .Y(_05442_));
 sky130_fd_sc_hd__o211ai_4 _15824_ (.A1(_05433_),
    .A2(_05441_),
    .B1(_05014_),
    .C1(_05429_),
    .Y(_05443_));
 sky130_fd_sc_hd__o21ai_1 _15825_ (.A1(_05440_),
    .A2(_05443_),
    .B1(_05442_),
    .Y(_05444_));
 sky130_fd_sc_hd__nand2_1 _15826_ (.A(net29),
    .B(net48),
    .Y(_05445_));
 sky130_fd_sc_hd__a22oi_4 _15827_ (.A1(net31),
    .A2(net46),
    .B1(net47),
    .B2(net30),
    .Y(_05446_));
 sky130_fd_sc_hd__a22o_1 _15828_ (.A1(net31),
    .A2(net46),
    .B1(net47),
    .B2(net30),
    .X(_05448_));
 sky130_fd_sc_hd__and4_1 _15829_ (.A(net30),
    .B(net31),
    .C(net46),
    .D(net47),
    .X(_05449_));
 sky130_fd_sc_hd__nand4_2 _15830_ (.A(net30),
    .B(net31),
    .C(net46),
    .D(net47),
    .Y(_05450_));
 sky130_fd_sc_hd__a22oi_2 _15831_ (.A1(net29),
    .A2(net48),
    .B1(_05448_),
    .B2(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__nor3_2 _15832_ (.A(_05445_),
    .B(_05446_),
    .C(_05449_),
    .Y(_05452_));
 sky130_fd_sc_hd__nor2_2 _15833_ (.A(_05451_),
    .B(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__o21ai_2 _15834_ (.A1(_05451_),
    .A2(_05452_),
    .B1(_05444_),
    .Y(_05454_));
 sky130_fd_sc_hd__o211ai_4 _15835_ (.A1(_05440_),
    .A2(_05443_),
    .B1(_05453_),
    .C1(_05442_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand2_2 _15836_ (.A(_05454_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__o21ai_1 _15837_ (.A1(_05424_),
    .A2(_05427_),
    .B1(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__and4_1 _15838_ (.A(_05426_),
    .B(_05428_),
    .C(_05454_),
    .D(_05455_),
    .X(_05459_));
 sky130_fd_sc_hd__nand4_2 _15839_ (.A(_05426_),
    .B(_05428_),
    .C(_05454_),
    .D(_05455_),
    .Y(_05460_));
 sky130_fd_sc_hd__o21bai_4 _15840_ (.A1(_05424_),
    .A2(_05427_),
    .B1_N(_05456_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand3_2 _15841_ (.A(_05426_),
    .B(_05428_),
    .C(_05456_),
    .Y(_05462_));
 sky130_fd_sc_hd__a21oi_4 _15842_ (.A1(_04945_),
    .A2(_04949_),
    .B1(_04947_),
    .Y(_05463_));
 sky130_fd_sc_hd__o2bb2ai_2 _15843_ (.A1_N(_04945_),
    .A2_N(_04949_),
    .B1(_04946_),
    .B2(_04939_),
    .Y(_05464_));
 sky130_fd_sc_hd__nand3_4 _15844_ (.A(_05461_),
    .B(_05463_),
    .C(_05462_),
    .Y(_05465_));
 sky130_fd_sc_hd__inv_2 _15845_ (.A(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__nand3_4 _15846_ (.A(_05457_),
    .B(_05460_),
    .C(_05464_),
    .Y(_05467_));
 sky130_fd_sc_hd__nand2_1 _15847_ (.A(_05465_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__o41a_1 _15848_ (.A1(_04534_),
    .A2(_04969_),
    .A3(_04991_),
    .A4(_04992_),
    .B1(_05032_),
    .X(_05470_));
 sky130_fd_sc_hd__o21a_2 _15849_ (.A1(_04995_),
    .A2(_05032_),
    .B1(_04994_),
    .X(_05471_));
 sky130_fd_sc_hd__nor2_1 _15850_ (.A(_05468_),
    .B(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand3b_2 _15851_ (.A_N(_05471_),
    .B(_05467_),
    .C(_05465_),
    .Y(_05473_));
 sky130_fd_sc_hd__o311a_1 _15852_ (.A1(_04995_),
    .A2(_05028_),
    .A3(_05029_),
    .B1(_05468_),
    .C1(_04994_),
    .X(_05474_));
 sky130_fd_sc_hd__o2bb2ai_2 _15853_ (.A1_N(_05465_),
    .A2_N(_05467_),
    .B1(_05470_),
    .B2(_04995_),
    .Y(_05475_));
 sky130_fd_sc_hd__a21oi_2 _15854_ (.A1(_05465_),
    .A2(_05467_),
    .B1(_05471_),
    .Y(_05476_));
 sky130_fd_sc_hd__and3_1 _15855_ (.A(_05465_),
    .B(_05467_),
    .C(_05471_),
    .X(_05477_));
 sky130_fd_sc_hd__nand2_2 _15856_ (.A(_05473_),
    .B(_05475_),
    .Y(_05478_));
 sky130_fd_sc_hd__o211ai_2 _15857_ (.A1(_05393_),
    .A2(_05397_),
    .B1(_05478_),
    .C1(_05396_),
    .Y(_05479_));
 sky130_fd_sc_hd__o2bb2ai_2 _15858_ (.A1_N(_05396_),
    .A2_N(_05399_),
    .B1(_05476_),
    .B2(_05477_),
    .Y(_05481_));
 sky130_fd_sc_hd__o2bb2ai_4 _15859_ (.A1_N(_05396_),
    .A2_N(_05399_),
    .B1(_05472_),
    .B2(_05474_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21ai_1 _15860_ (.A1(_05476_),
    .A2(_05477_),
    .B1(_05396_),
    .Y(_05483_));
 sky130_fd_sc_hd__o211ai_4 _15861_ (.A1(_05476_),
    .A2(_05477_),
    .B1(_05396_),
    .C1(_05399_),
    .Y(_05484_));
 sky130_fd_sc_hd__a22oi_4 _15862_ (.A1(_04966_),
    .A2(_05252_),
    .B1(_05482_),
    .B2(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__nand3_2 _15863_ (.A(_05253_),
    .B(_05479_),
    .C(_05481_),
    .Y(_05486_));
 sky130_fd_sc_hd__o211a_2 _15864_ (.A1(_05483_),
    .A2(_05398_),
    .B1(_05254_),
    .C1(_05482_),
    .X(_05487_));
 sky130_fd_sc_hd__o2111ai_4 _15865_ (.A1(_04967_),
    .A2(_05054_),
    .B1(_05482_),
    .C1(_05484_),
    .D1(_04966_),
    .Y(_05488_));
 sky130_fd_sc_hd__o22ai_2 _15866_ (.A1(_05242_),
    .A2(_05244_),
    .B1(_05485_),
    .B2(_05487_),
    .Y(_05489_));
 sky130_fd_sc_hd__nand3_1 _15867_ (.A(_05488_),
    .B(_05250_),
    .C(_05486_),
    .Y(_05490_));
 sky130_fd_sc_hd__a31oi_2 _15868_ (.A1(_05253_),
    .A2(_05479_),
    .A3(_05481_),
    .B1(_05250_),
    .Y(_05492_));
 sky130_fd_sc_hd__o211ai_4 _15869_ (.A1(_05242_),
    .A2(_05244_),
    .B1(_05486_),
    .C1(_05488_),
    .Y(_05493_));
 sky130_fd_sc_hd__o22ai_4 _15870_ (.A1(_05245_),
    .A2(_05248_),
    .B1(_05485_),
    .B2(_05487_),
    .Y(_05494_));
 sky130_fd_sc_hd__a22oi_2 _15871_ (.A1(_05062_),
    .A2(_05138_),
    .B1(_05489_),
    .B2(_05490_),
    .Y(_05495_));
 sky130_fd_sc_hd__nand4_2 _15872_ (.A(_05061_),
    .B(_05169_),
    .C(_05493_),
    .D(_05494_),
    .Y(_05496_));
 sky130_fd_sc_hd__a22oi_4 _15873_ (.A1(_05061_),
    .A2(_05169_),
    .B1(_05493_),
    .B2(_05494_),
    .Y(_05497_));
 sky130_fd_sc_hd__nand3_1 _15874_ (.A(_05171_),
    .B(_05489_),
    .C(_05490_),
    .Y(_05498_));
 sky130_fd_sc_hd__nand2_1 _15875_ (.A(_05496_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__nand3_1 _15876_ (.A(_05496_),
    .B(_05498_),
    .C(_05168_),
    .Y(_05500_));
 sky130_fd_sc_hd__o22ai_2 _15877_ (.A1(_05124_),
    .A2(_05131_),
    .B1(_05495_),
    .B2(_05497_),
    .Y(_05501_));
 sky130_fd_sc_hd__o211ai_2 _15878_ (.A1(_05124_),
    .A2(_05131_),
    .B1(_05496_),
    .C1(_05498_),
    .Y(_05503_));
 sky130_fd_sc_hd__o21bai_1 _15879_ (.A1(_05495_),
    .A2(_05497_),
    .B1_N(_05167_),
    .Y(_05504_));
 sky130_fd_sc_hd__a2bb2oi_1 _15880_ (.A1_N(_05143_),
    .A2_N(_05147_),
    .B1(_05168_),
    .B2(_05499_),
    .Y(_05505_));
 sky130_fd_sc_hd__nand3_2 _15881_ (.A(_05504_),
    .B(_05166_),
    .C(_05503_),
    .Y(_05506_));
 sky130_fd_sc_hd__o2111ai_4 _15882_ (.A1(_05146_),
    .A2(_05140_),
    .B1(_05144_),
    .C1(_05500_),
    .D1(_05501_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_1 _15883_ (.A(_05506_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__nand4b_1 _15884_ (.A_N(_05156_),
    .B(_05506_),
    .C(_05507_),
    .D(_05148_),
    .Y(_05509_));
 sky130_fd_sc_hd__o2bb2ai_1 _15885_ (.A1_N(_05506_),
    .A2_N(_05507_),
    .B1(_05153_),
    .B2(_05154_),
    .Y(_05510_));
 sky130_fd_sc_hd__and2_1 _15886_ (.A(_05509_),
    .B(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__o2bb2a_1 _15887_ (.A1_N(_05161_),
    .A2_N(_05165_),
    .B1(_05157_),
    .B2(_05160_),
    .X(_05512_));
 sky130_fd_sc_hd__o2111a_2 _15888_ (.A1(_05157_),
    .A2(_05160_),
    .B1(_05509_),
    .C1(_05510_),
    .D1(_05159_),
    .X(_05514_));
 sky130_fd_sc_hd__xnor2_1 _15889_ (.A(_05511_),
    .B(_05512_),
    .Y(net86));
 sky130_fd_sc_hd__a31oi_1 _15890_ (.A1(_05170_),
    .A2(_05493_),
    .A3(_05494_),
    .B1(_05167_),
    .Y(_05515_));
 sky130_fd_sc_hd__o21ai_1 _15891_ (.A1(_05168_),
    .A2(_05497_),
    .B1(_05496_),
    .Y(_05516_));
 sky130_fd_sc_hd__a31o_1 _15892_ (.A1(_05125_),
    .A2(_05132_),
    .A3(_05496_),
    .B1(_05497_),
    .X(_05517_));
 sky130_fd_sc_hd__a32oi_4 _15893_ (.A1(_05254_),
    .A2(_05482_),
    .A3(_05484_),
    .B1(_05486_),
    .B2(_05251_),
    .Y(_05518_));
 sky130_fd_sc_hd__nand2_4 _15894_ (.A(net12),
    .B(net54),
    .Y(_05519_));
 sky130_fd_sc_hd__nand2_1 _15895_ (.A(net26),
    .B(net53),
    .Y(_05520_));
 sky130_fd_sc_hd__and4_1 _15896_ (.A(net26),
    .B(net23),
    .C(net52),
    .D(net53),
    .X(_05521_));
 sky130_fd_sc_hd__nand4_2 _15897_ (.A(net26),
    .B(net23),
    .C(net52),
    .D(net53),
    .Y(_05522_));
 sky130_fd_sc_hd__a22oi_4 _15898_ (.A1(net26),
    .A2(net52),
    .B1(net53),
    .B2(net23),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_1 _15899_ (.A1(_05521_),
    .A2(_05524_),
    .B1(_05519_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand4b_1 _15900_ (.A_N(_05524_),
    .B(net54),
    .C(net12),
    .D(_05522_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_2 _15901_ (.A(_05525_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21oi_2 _15902_ (.A1(_05215_),
    .A2(_05218_),
    .B1(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__a21o_1 _15903_ (.A1(_05215_),
    .A2(_05218_),
    .B1(_05527_),
    .X(_05529_));
 sky130_fd_sc_hd__nand3_1 _15904_ (.A(_05527_),
    .B(_05218_),
    .C(_05215_),
    .Y(_05530_));
 sky130_fd_sc_hd__a22o_2 _15905_ (.A1(net1),
    .A2(net56),
    .B1(_05529_),
    .B2(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__nand4_4 _15906_ (.A(_05529_),
    .B(_05530_),
    .C(net1),
    .D(net56),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _15907_ (.A(_05531_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__a22oi_4 _15908_ (.A1(_05111_),
    .A2(_05220_),
    .B1(_05531_),
    .B2(_05532_),
    .Y(_05535_));
 sky130_fd_sc_hd__inv_2 _15909_ (.A(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__and3_2 _15910_ (.A(_05222_),
    .B(_05531_),
    .C(_05532_),
    .X(_05537_));
 sky130_fd_sc_hd__nand4_4 _15911_ (.A(_05531_),
    .B(_05532_),
    .C(_05111_),
    .D(_05220_),
    .Y(_05538_));
 sky130_fd_sc_hd__nand2_1 _15912_ (.A(_05202_),
    .B(_05175_),
    .Y(_05539_));
 sky130_fd_sc_hd__nand2_1 _15913_ (.A(_05204_),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__o2bb2ai_4 _15914_ (.A1_N(_05442_),
    .A2_N(_05453_),
    .B1(_05443_),
    .B2(_05440_),
    .Y(_05541_));
 sky130_fd_sc_hd__o32a_1 _15915_ (.A1(_01769_),
    .A2(_02120_),
    .A3(_05180_),
    .B1(_02152_),
    .B2(_01791_),
    .X(_05542_));
 sky130_fd_sc_hd__and3_1 _15916_ (.A(_05185_),
    .B(net51),
    .C(net26),
    .X(_05543_));
 sky130_fd_sc_hd__a31o_1 _15917_ (.A1(_05185_),
    .A2(net51),
    .A3(net26),
    .B1(_05181_),
    .X(_05544_));
 sky130_fd_sc_hd__nor2_1 _15918_ (.A(_05445_),
    .B(_05446_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21ai_2 _15919_ (.A1(_05445_),
    .A2(_05446_),
    .B1(_05450_),
    .Y(_05547_));
 sky130_fd_sc_hd__o21a_1 _15920_ (.A1(_05445_),
    .A2(_05446_),
    .B1(_05450_),
    .X(_05548_));
 sky130_fd_sc_hd__nor2_1 _15921_ (.A(_01769_),
    .B(_02152_),
    .Y(_05549_));
 sky130_fd_sc_hd__a22oi_4 _15922_ (.A1(net29),
    .A2(net49),
    .B1(net50),
    .B2(net28),
    .Y(_05550_));
 sky130_fd_sc_hd__a22o_2 _15923_ (.A1(net29),
    .A2(net49),
    .B1(net50),
    .B2(net28),
    .X(_05551_));
 sky130_fd_sc_hd__nand2_4 _15924_ (.A(net29),
    .B(net50),
    .Y(_05552_));
 sky130_fd_sc_hd__and4_1 _15925_ (.A(net28),
    .B(net29),
    .C(net49),
    .D(net50),
    .X(_05553_));
 sky130_fd_sc_hd__o221ai_4 _15926_ (.A1(_01769_),
    .A2(_02152_),
    .B1(_05182_),
    .B2(_05552_),
    .C1(_05551_),
    .Y(_05554_));
 sky130_fd_sc_hd__o21ai_2 _15927_ (.A1(_05550_),
    .A2(_05553_),
    .B1(_05549_),
    .Y(_05555_));
 sky130_fd_sc_hd__o2111ai_4 _15928_ (.A1(_05182_),
    .A2(_05552_),
    .B1(net27),
    .C1(net51),
    .D1(_05551_),
    .Y(_05557_));
 sky130_fd_sc_hd__o22ai_4 _15929_ (.A1(_01769_),
    .A2(_02152_),
    .B1(_05550_),
    .B2(_05553_),
    .Y(_05558_));
 sky130_fd_sc_hd__a2bb2oi_4 _15930_ (.A1_N(_05449_),
    .A2_N(_05546_),
    .B1(_05554_),
    .B2(_05555_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand3_4 _15931_ (.A(_05558_),
    .B(_05547_),
    .C(_05557_),
    .Y(_05560_));
 sky130_fd_sc_hd__a21oi_2 _15932_ (.A1(_05557_),
    .A2(_05558_),
    .B1(_05547_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand3_4 _15933_ (.A(_05548_),
    .B(_05554_),
    .C(_05555_),
    .Y(_05562_));
 sky130_fd_sc_hd__o21ai_2 _15934_ (.A1(_05181_),
    .A2(_05543_),
    .B1(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__o211a_2 _15935_ (.A1(_05181_),
    .A2(_05543_),
    .B1(_05560_),
    .C1(_05562_),
    .X(_05564_));
 sky130_fd_sc_hd__o211ai_4 _15936_ (.A1(_05181_),
    .A2(_05543_),
    .B1(_05560_),
    .C1(_05562_),
    .Y(_05565_));
 sky130_fd_sc_hd__a21oi_1 _15937_ (.A1(_05560_),
    .A2(_05562_),
    .B1(_05544_),
    .Y(_05566_));
 sky130_fd_sc_hd__o22ai_4 _15938_ (.A1(_05184_),
    .A2(_05542_),
    .B1(_05559_),
    .B2(_05561_),
    .Y(_05568_));
 sky130_fd_sc_hd__a21oi_4 _15939_ (.A1(_05565_),
    .A2(_05568_),
    .B1(_05541_),
    .Y(_05569_));
 sky130_fd_sc_hd__o21bai_4 _15940_ (.A1(_05564_),
    .A2(_05566_),
    .B1_N(_05541_),
    .Y(_05570_));
 sky130_fd_sc_hd__nand2_1 _15941_ (.A(_05541_),
    .B(_05568_),
    .Y(_05571_));
 sky130_fd_sc_hd__o211a_2 _15942_ (.A1(_05563_),
    .A2(_05559_),
    .B1(_05541_),
    .C1(_05568_),
    .X(_05572_));
 sky130_fd_sc_hd__o211ai_4 _15943_ (.A1(_05563_),
    .A2(_05559_),
    .B1(_05541_),
    .C1(_05568_),
    .Y(_05573_));
 sky130_fd_sc_hd__o311a_1 _15944_ (.A1(_01802_),
    .A2(_05074_),
    .A3(_02152_),
    .B1(_05073_),
    .C1(_05192_),
    .X(_05574_));
 sky130_fd_sc_hd__o31a_1 _15945_ (.A1(_05072_),
    .A2(_05176_),
    .A3(_05191_),
    .B1(_05195_),
    .X(_05575_));
 sky130_fd_sc_hd__o21a_1 _15946_ (.A1(_05177_),
    .A2(_05193_),
    .B1(_05192_),
    .X(_05576_));
 sky130_fd_sc_hd__o2bb2ai_2 _15947_ (.A1_N(_05570_),
    .A2_N(_05573_),
    .B1(_05574_),
    .B2(_05193_),
    .Y(_05577_));
 sky130_fd_sc_hd__o21ai_4 _15948_ (.A1(_05191_),
    .A2(_05196_),
    .B1(_05570_),
    .Y(_05579_));
 sky130_fd_sc_hd__o221ai_4 _15949_ (.A1(_05191_),
    .A2(_05196_),
    .B1(_05564_),
    .B2(_05571_),
    .C1(_05570_),
    .Y(_05580_));
 sky130_fd_sc_hd__o22ai_4 _15950_ (.A1(_05191_),
    .A2(_05196_),
    .B1(_05569_),
    .B2(_05572_),
    .Y(_05581_));
 sky130_fd_sc_hd__o2111ai_4 _15951_ (.A1(_05193_),
    .A2(_05177_),
    .B1(_05192_),
    .C1(_05570_),
    .D1(_05573_),
    .Y(_05582_));
 sky130_fd_sc_hd__a22oi_4 _15952_ (.A1(_05204_),
    .A2(_05539_),
    .B1(_05577_),
    .B2(_05580_),
    .Y(_05583_));
 sky130_fd_sc_hd__nand3_2 _15953_ (.A(_05540_),
    .B(_05581_),
    .C(_05582_),
    .Y(_05584_));
 sky130_fd_sc_hd__a21oi_4 _15954_ (.A1(_05581_),
    .A2(_05582_),
    .B1(_05540_),
    .Y(_05585_));
 sky130_fd_sc_hd__o221ai_4 _15955_ (.A1(_05572_),
    .A2(_05579_),
    .B1(_05201_),
    .B2(_05206_),
    .C1(_05577_),
    .Y(_05586_));
 sky130_fd_sc_hd__o22ai_4 _15956_ (.A1(_05535_),
    .A2(_05537_),
    .B1(_05583_),
    .B2(_05585_),
    .Y(_05587_));
 sky130_fd_sc_hd__and3_1 _15957_ (.A(_05536_),
    .B(_05538_),
    .C(_05584_),
    .X(_05588_));
 sky130_fd_sc_hd__nand3_2 _15958_ (.A(_05536_),
    .B(_05538_),
    .C(_05584_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand4_4 _15959_ (.A(_05536_),
    .B(_05538_),
    .C(_05584_),
    .D(_05586_),
    .Y(_05591_));
 sky130_fd_sc_hd__o211a_1 _15960_ (.A1(_04995_),
    .A2(_05032_),
    .B1(_05467_),
    .C1(_04994_),
    .X(_05592_));
 sky130_fd_sc_hd__a32oi_4 _15961_ (.A1(_05461_),
    .A2(_05462_),
    .A3(_05463_),
    .B1(_05467_),
    .B2(_05471_),
    .Y(_05593_));
 sky130_fd_sc_hd__a21oi_4 _15962_ (.A1(_05587_),
    .A2(_05591_),
    .B1(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__o2bb2ai_2 _15963_ (.A1_N(_05587_),
    .A2_N(_05591_),
    .B1(_05592_),
    .B2(_05466_),
    .Y(_05595_));
 sky130_fd_sc_hd__o211a_2 _15964_ (.A1(_05585_),
    .A2(_05590_),
    .B1(_05593_),
    .C1(_05587_),
    .X(_05596_));
 sky130_fd_sc_hd__o211ai_4 _15965_ (.A1(_05585_),
    .A2(_05590_),
    .B1(_05593_),
    .C1(_05587_),
    .Y(_05597_));
 sky130_fd_sc_hd__a31o_1 _15966_ (.A1(_05211_),
    .A2(_05221_),
    .A3(_05224_),
    .B1(_05212_),
    .X(_05598_));
 sky130_fd_sc_hd__a32o_2 _15967_ (.A1(_05174_),
    .A2(_05209_),
    .A3(_05210_),
    .B1(_05213_),
    .B2(_05228_),
    .X(_05599_));
 sky130_fd_sc_hd__a21oi_1 _15968_ (.A1(_05595_),
    .A2(_05597_),
    .B1(_05598_),
    .Y(_05601_));
 sky130_fd_sc_hd__o21ai_4 _15969_ (.A1(_05594_),
    .A2(_05596_),
    .B1(_05599_),
    .Y(_05602_));
 sky130_fd_sc_hd__o311a_1 _15970_ (.A1(_05212_),
    .A2(_05225_),
    .A3(_05226_),
    .B1(_05595_),
    .C1(_05211_),
    .X(_05603_));
 sky130_fd_sc_hd__nand2_1 _15971_ (.A(_05595_),
    .B(_05598_),
    .Y(_05604_));
 sky130_fd_sc_hd__and3_1 _15972_ (.A(_05595_),
    .B(_05597_),
    .C(_05598_),
    .X(_05605_));
 sky130_fd_sc_hd__nand3_2 _15973_ (.A(_05595_),
    .B(_05597_),
    .C(_05598_),
    .Y(_05606_));
 sky130_fd_sc_hd__a21oi_1 _15974_ (.A1(_05595_),
    .A2(_05597_),
    .B1(_05599_),
    .Y(_05607_));
 sky130_fd_sc_hd__and3_1 _15975_ (.A(_05595_),
    .B(_05597_),
    .C(_05599_),
    .X(_05608_));
 sky130_fd_sc_hd__o21ai_1 _15976_ (.A1(_05596_),
    .A2(_05604_),
    .B1(_05602_),
    .Y(_05609_));
 sky130_fd_sc_hd__a32oi_4 _15977_ (.A1(_05256_),
    .A2(_05391_),
    .A3(_05394_),
    .B1(_05473_),
    .B2(_05475_),
    .Y(_05610_));
 sky130_fd_sc_hd__nand2_1 _15978_ (.A(_05399_),
    .B(_05478_),
    .Y(_05612_));
 sky130_fd_sc_hd__o22ai_4 _15979_ (.A1(_05393_),
    .A2(_05397_),
    .B1(_05478_),
    .B2(_05395_),
    .Y(_05613_));
 sky130_fd_sc_hd__a32oi_4 _15980_ (.A1(_05261_),
    .A2(_05336_),
    .A3(_05338_),
    .B1(_05385_),
    .B2(_05388_),
    .Y(_05614_));
 sky130_fd_sc_hd__o21ai_4 _15981_ (.A1(_05384_),
    .A2(_05387_),
    .B1(_05341_),
    .Y(_05615_));
 sky130_fd_sc_hd__a31o_2 _15982_ (.A1(_05269_),
    .A2(net14),
    .A3(net63),
    .B1(_05266_),
    .X(_05616_));
 sky130_fd_sc_hd__o21ai_2 _15983_ (.A1(_05309_),
    .A2(_05310_),
    .B1(_05313_),
    .Y(_05617_));
 sky130_fd_sc_hd__nand2_1 _15984_ (.A(net63),
    .B(net15),
    .Y(_05618_));
 sky130_fd_sc_hd__a22oi_4 _15985_ (.A1(net62),
    .A2(net16),
    .B1(net17),
    .B2(net61),
    .Y(_05619_));
 sky130_fd_sc_hd__a22o_1 _15986_ (.A1(net62),
    .A2(net16),
    .B1(net17),
    .B2(net61),
    .X(_05620_));
 sky130_fd_sc_hd__nand2_2 _15987_ (.A(net62),
    .B(net17),
    .Y(_05621_));
 sky130_fd_sc_hd__and4_1 _15988_ (.A(net61),
    .B(net62),
    .C(net16),
    .D(net17),
    .X(_05623_));
 sky130_fd_sc_hd__o221ai_4 _15989_ (.A1(_01890_),
    .A2(_02076_),
    .B1(_05265_),
    .B2(_05621_),
    .C1(_05620_),
    .Y(_05624_));
 sky130_fd_sc_hd__o21bai_1 _15990_ (.A1(_05619_),
    .A2(_05623_),
    .B1_N(_05618_),
    .Y(_05625_));
 sky130_fd_sc_hd__o21ai_2 _15991_ (.A1(_05619_),
    .A2(_05623_),
    .B1(_05618_),
    .Y(_05626_));
 sky130_fd_sc_hd__a41o_1 _15992_ (.A1(net61),
    .A2(net62),
    .A3(net16),
    .A4(net17),
    .B1(_05618_),
    .X(_05627_));
 sky130_fd_sc_hd__o211a_2 _15993_ (.A1(_05619_),
    .A2(_05627_),
    .B1(_05617_),
    .C1(_05626_),
    .X(_05628_));
 sky130_fd_sc_hd__o211ai_4 _15994_ (.A1(_05619_),
    .A2(_05627_),
    .B1(_05617_),
    .C1(_05626_),
    .Y(_05629_));
 sky130_fd_sc_hd__nand3b_4 _15995_ (.A_N(_05617_),
    .B(_05624_),
    .C(_05625_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_2 _15996_ (.A(_05630_),
    .B(_05616_),
    .Y(_05631_));
 sky130_fd_sc_hd__and3_2 _15997_ (.A(_05630_),
    .B(_05616_),
    .C(_05629_),
    .X(_05632_));
 sky130_fd_sc_hd__a21oi_4 _15998_ (.A1(_05629_),
    .A2(_05630_),
    .B1(_05616_),
    .Y(_05634_));
 sky130_fd_sc_hd__a21o_1 _15999_ (.A1(_05629_),
    .A2(_05630_),
    .B1(_05616_),
    .X(_05635_));
 sky130_fd_sc_hd__o21ai_2 _16000_ (.A1(_05628_),
    .A2(_05631_),
    .B1(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__nor2_1 _16001_ (.A(_05292_),
    .B(_05295_),
    .Y(_05637_));
 sky130_fd_sc_hd__o21a_2 _16002_ (.A1(_05292_),
    .A2(_05295_),
    .B1(_05298_),
    .X(_05638_));
 sky130_fd_sc_hd__nand2_4 _16003_ (.A(net55),
    .B(net21),
    .Y(_05639_));
 sky130_fd_sc_hd__a22oi_4 _16004_ (.A1(net44),
    .A2(net22),
    .B1(net24),
    .B2(net33),
    .Y(_05640_));
 sky130_fd_sc_hd__a22o_1 _16005_ (.A1(net44),
    .A2(net22),
    .B1(net24),
    .B2(net33),
    .X(_05641_));
 sky130_fd_sc_hd__nand2_2 _16006_ (.A(net44),
    .B(net24),
    .Y(_05642_));
 sky130_fd_sc_hd__and4_2 _16007_ (.A(net33),
    .B(net44),
    .C(net22),
    .D(net24),
    .X(_05643_));
 sky130_fd_sc_hd__o221ai_4 _16008_ (.A1(_01780_),
    .A2(_02185_),
    .B1(_05294_),
    .B2(_05642_),
    .C1(_05641_),
    .Y(_05645_));
 sky130_fd_sc_hd__o21bai_1 _16009_ (.A1(_05640_),
    .A2(_05643_),
    .B1_N(_05639_),
    .Y(_05646_));
 sky130_fd_sc_hd__o21ai_4 _16010_ (.A1(_05640_),
    .A2(_05643_),
    .B1(_05639_),
    .Y(_05647_));
 sky130_fd_sc_hd__a41o_2 _16011_ (.A1(net33),
    .A2(net44),
    .A3(net22),
    .A4(net24),
    .B1(_05639_),
    .X(_05648_));
 sky130_fd_sc_hd__o21ai_4 _16012_ (.A1(_05640_),
    .A2(_05648_),
    .B1(_05647_),
    .Y(_05649_));
 sky130_fd_sc_hd__nand3_4 _16013_ (.A(_05638_),
    .B(_05645_),
    .C(_05646_),
    .Y(_05650_));
 sky130_fd_sc_hd__o221a_4 _16014_ (.A1(_05640_),
    .A2(_05648_),
    .B1(_05297_),
    .B2(_05637_),
    .C1(_05647_),
    .X(_05651_));
 sky130_fd_sc_hd__o221ai_4 _16015_ (.A1(_05640_),
    .A2(_05648_),
    .B1(_05297_),
    .B2(_05637_),
    .C1(_05647_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(net60),
    .B(net18),
    .Y(_05653_));
 sky130_fd_sc_hd__a22oi_2 _16017_ (.A1(net59),
    .A2(net19),
    .B1(net20),
    .B2(net58),
    .Y(_05654_));
 sky130_fd_sc_hd__a22o_1 _16018_ (.A1(net59),
    .A2(net19),
    .B1(net20),
    .B2(net58),
    .X(_05656_));
 sky130_fd_sc_hd__nand2_1 _16019_ (.A(net59),
    .B(net20),
    .Y(_05657_));
 sky130_fd_sc_hd__and4_1 _16020_ (.A(net58),
    .B(net59),
    .C(net19),
    .D(net20),
    .X(_05658_));
 sky130_fd_sc_hd__nand4_4 _16021_ (.A(net58),
    .B(net59),
    .C(net19),
    .D(net20),
    .Y(_05659_));
 sky130_fd_sc_hd__and3_2 _16022_ (.A(_05653_),
    .B(_05656_),
    .C(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__o211ai_4 _16023_ (.A1(_01835_),
    .A2(_02131_),
    .B1(_05656_),
    .C1(_05659_),
    .Y(_05661_));
 sky130_fd_sc_hd__o211a_2 _16024_ (.A1(_05654_),
    .A2(_05658_),
    .B1(net60),
    .C1(net18),
    .X(_05662_));
 sky130_fd_sc_hd__a21o_2 _16025_ (.A1(_05656_),
    .A2(_05659_),
    .B1(_05653_),
    .X(_05663_));
 sky130_fd_sc_hd__o22a_1 _16026_ (.A1(_01835_),
    .A2(_02131_),
    .B1(_05654_),
    .B2(_05658_),
    .X(_05664_));
 sky130_fd_sc_hd__and4_1 _16027_ (.A(_05656_),
    .B(_05659_),
    .C(net60),
    .D(net18),
    .X(_05665_));
 sky130_fd_sc_hd__nand2_1 _16028_ (.A(_05661_),
    .B(_05663_),
    .Y(_05667_));
 sky130_fd_sc_hd__o2bb2ai_4 _16029_ (.A1_N(_05650_),
    .A2_N(_05652_),
    .B1(_05660_),
    .B2(_05662_),
    .Y(_05668_));
 sky130_fd_sc_hd__nand4_4 _16030_ (.A(_05650_),
    .B(_05652_),
    .C(_05661_),
    .D(_05663_),
    .Y(_05669_));
 sky130_fd_sc_hd__o2bb2ai_2 _16031_ (.A1_N(_05650_),
    .A2_N(_05652_),
    .B1(_05664_),
    .B2(_05665_),
    .Y(_05670_));
 sky130_fd_sc_hd__a22oi_4 _16032_ (.A1(_05661_),
    .A2(_05663_),
    .B1(_05649_),
    .B2(_05638_),
    .Y(_05671_));
 sky130_fd_sc_hd__o21ai_2 _16033_ (.A1(_05660_),
    .A2(_05662_),
    .B1(_05650_),
    .Y(_05672_));
 sky130_fd_sc_hd__o211ai_2 _16034_ (.A1(_05660_),
    .A2(_05662_),
    .B1(_05650_),
    .C1(_05652_),
    .Y(_05673_));
 sky130_fd_sc_hd__a2bb2oi_2 _16035_ (.A1_N(_05301_),
    .A2_N(_05306_),
    .B1(_05322_),
    .B2(_05305_),
    .Y(_05674_));
 sky130_fd_sc_hd__o2bb2ai_4 _16036_ (.A1_N(_05305_),
    .A2_N(_05322_),
    .B1(_05306_),
    .B2(_05301_),
    .Y(_05675_));
 sky130_fd_sc_hd__a22oi_2 _16037_ (.A1(_05307_),
    .A2(_05323_),
    .B1(_05668_),
    .B2(_05669_),
    .Y(_05676_));
 sky130_fd_sc_hd__o211ai_4 _16038_ (.A1(_05651_),
    .A2(_05672_),
    .B1(_05675_),
    .C1(_05670_),
    .Y(_05678_));
 sky130_fd_sc_hd__a21oi_4 _16039_ (.A1(_05670_),
    .A2(_05673_),
    .B1(_05675_),
    .Y(_05679_));
 sky130_fd_sc_hd__nand3_2 _16040_ (.A(_05668_),
    .B(_05674_),
    .C(_05669_),
    .Y(_05680_));
 sky130_fd_sc_hd__o21a_1 _16041_ (.A1(_05632_),
    .A2(_05634_),
    .B1(_05678_),
    .X(_05681_));
 sky130_fd_sc_hd__a32oi_4 _16042_ (.A1(_05668_),
    .A2(_05674_),
    .A3(_05669_),
    .B1(_05636_),
    .B2(_05678_),
    .Y(_05682_));
 sky130_fd_sc_hd__a21o_1 _16043_ (.A1(_05678_),
    .A2(_05680_),
    .B1(_05636_),
    .X(_05683_));
 sky130_fd_sc_hd__o211ai_4 _16044_ (.A1(_05632_),
    .A2(_05634_),
    .B1(_05678_),
    .C1(_05680_),
    .Y(_05684_));
 sky130_fd_sc_hd__o22ai_4 _16045_ (.A1(_05632_),
    .A2(_05634_),
    .B1(_05676_),
    .B2(_05679_),
    .Y(_05685_));
 sky130_fd_sc_hd__o2111ai_4 _16046_ (.A1(_05628_),
    .A2(_05631_),
    .B1(_05635_),
    .C1(_05678_),
    .D1(_05680_),
    .Y(_05686_));
 sky130_fd_sc_hd__a32oi_4 _16047_ (.A1(_05328_),
    .A2(_05329_),
    .A3(_05331_),
    .B1(_05335_),
    .B2(_05289_),
    .Y(_05687_));
 sky130_fd_sc_hd__a2bb2oi_4 _16048_ (.A1_N(_05324_),
    .A2_N(_05334_),
    .B1(_05333_),
    .B2(_05288_),
    .Y(_05689_));
 sky130_fd_sc_hd__and3_1 _16049_ (.A(_05685_),
    .B(_05687_),
    .C(_05686_),
    .X(_05690_));
 sky130_fd_sc_hd__nand3_4 _16050_ (.A(_05685_),
    .B(_05687_),
    .C(_05686_),
    .Y(_05691_));
 sky130_fd_sc_hd__nand3_4 _16051_ (.A(_05683_),
    .B(_05684_),
    .C(_05689_),
    .Y(_05692_));
 sky130_fd_sc_hd__a21boi_4 _16052_ (.A1(_05276_),
    .A2(_05281_),
    .B1_N(_05278_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_4 _16053_ (.A1(_05356_),
    .A2(_05357_),
    .B1(_05361_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_2 _16054_ (.A(net35),
    .B(net11),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_1 _16055_ (.A(net34),
    .B(net14),
    .Y(_05696_));
 sky130_fd_sc_hd__and4_1 _16056_ (.A(net64),
    .B(net34),
    .C(net13),
    .D(net14),
    .X(_05697_));
 sky130_fd_sc_hd__nand4_2 _16057_ (.A(net64),
    .B(net34),
    .C(net13),
    .D(net14),
    .Y(_05698_));
 sky130_fd_sc_hd__a22oi_4 _16058_ (.A1(net34),
    .A2(net13),
    .B1(net14),
    .B2(net64),
    .Y(_05700_));
 sky130_fd_sc_hd__a22o_1 _16059_ (.A1(net34),
    .A2(net13),
    .B1(net14),
    .B2(net64),
    .X(_05701_));
 sky130_fd_sc_hd__o211ai_2 _16060_ (.A1(_01934_),
    .A2(_02032_),
    .B1(_05698_),
    .C1(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__o21bai_2 _16061_ (.A1(_05697_),
    .A2(_05700_),
    .B1_N(_05695_),
    .Y(_05703_));
 sky130_fd_sc_hd__o22a_2 _16062_ (.A1(_01934_),
    .A2(_02032_),
    .B1(_05697_),
    .B2(_05700_),
    .X(_05704_));
 sky130_fd_sc_hd__o21ai_1 _16063_ (.A1(_05697_),
    .A2(_05700_),
    .B1(_05695_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand4_2 _16064_ (.A(_05701_),
    .B(net11),
    .C(net35),
    .D(_05698_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand2_2 _16065_ (.A(_05694_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand3_2 _16066_ (.A(_05705_),
    .B(_05706_),
    .C(_05694_),
    .Y(_05708_));
 sky130_fd_sc_hd__a21oi_2 _16067_ (.A1(_05705_),
    .A2(_05706_),
    .B1(_05694_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand3b_4 _16068_ (.A_N(_05694_),
    .B(_05702_),
    .C(_05703_),
    .Y(_05711_));
 sky130_fd_sc_hd__nand2_1 _16069_ (.A(net38),
    .B(net8),
    .Y(_05712_));
 sky130_fd_sc_hd__a22oi_2 _16070_ (.A1(net37),
    .A2(net9),
    .B1(net10),
    .B2(net36),
    .Y(_05713_));
 sky130_fd_sc_hd__a22o_1 _16071_ (.A1(net37),
    .A2(net9),
    .B1(net10),
    .B2(net36),
    .X(_05714_));
 sky130_fd_sc_hd__nand2_2 _16072_ (.A(net37),
    .B(net10),
    .Y(_05715_));
 sky130_fd_sc_hd__and4_1 _16073_ (.A(net36),
    .B(net37),
    .C(net9),
    .D(net10),
    .X(_05716_));
 sky130_fd_sc_hd__nand4_2 _16074_ (.A(net36),
    .B(net37),
    .C(net9),
    .D(net10),
    .Y(_05717_));
 sky130_fd_sc_hd__and3_1 _16075_ (.A(_05712_),
    .B(_05714_),
    .C(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nand3_1 _16076_ (.A(_05712_),
    .B(_05714_),
    .C(_05717_),
    .Y(_05719_));
 sky130_fd_sc_hd__o211a_1 _16077_ (.A1(_05713_),
    .A2(_05716_),
    .B1(net38),
    .C1(net8),
    .X(_05720_));
 sky130_fd_sc_hd__a21o_1 _16078_ (.A1(_05714_),
    .A2(_05717_),
    .B1(_05712_),
    .X(_05722_));
 sky130_fd_sc_hd__o2bb2a_1 _16079_ (.A1_N(net38),
    .A2_N(net8),
    .B1(_05713_),
    .B2(_05716_),
    .X(_05723_));
 sky130_fd_sc_hd__and4_1 _16080_ (.A(_05714_),
    .B(_05717_),
    .C(net38),
    .D(net8),
    .X(_05724_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(_05719_),
    .B(_05722_),
    .Y(_05725_));
 sky130_fd_sc_hd__o221ai_4 _16082_ (.A1(_05704_),
    .A2(_05707_),
    .B1(_05723_),
    .B2(_05724_),
    .C1(_05711_),
    .Y(_05726_));
 sky130_fd_sc_hd__o2bb2ai_4 _16083_ (.A1_N(_05708_),
    .A2_N(_05711_),
    .B1(_05718_),
    .B2(_05720_),
    .Y(_05727_));
 sky130_fd_sc_hd__o2bb2ai_2 _16084_ (.A1_N(_05708_),
    .A2_N(_05711_),
    .B1(_05723_),
    .B2(_05724_),
    .Y(_05728_));
 sky130_fd_sc_hd__o21ai_2 _16085_ (.A1(_05704_),
    .A2(_05707_),
    .B1(_05725_),
    .Y(_05729_));
 sky130_fd_sc_hd__nand3_2 _16086_ (.A(_05727_),
    .B(_05693_),
    .C(_05726_),
    .Y(_05730_));
 sky130_fd_sc_hd__o221a_2 _16087_ (.A1(_05709_),
    .A2(_05729_),
    .B1(_05277_),
    .B2(_05285_),
    .C1(_05728_),
    .X(_05731_));
 sky130_fd_sc_hd__o221ai_4 _16088_ (.A1(_05709_),
    .A2(_05729_),
    .B1(_05277_),
    .B2(_05285_),
    .C1(_05728_),
    .Y(_05733_));
 sky130_fd_sc_hd__a21oi_4 _16089_ (.A1(_05353_),
    .A2(_05368_),
    .B1(_05367_),
    .Y(_05734_));
 sky130_fd_sc_hd__a21oi_2 _16090_ (.A1(_05730_),
    .A2(_05733_),
    .B1(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__a22o_1 _16091_ (.A1(_05366_),
    .A2(_05373_),
    .B1(_05730_),
    .B2(_05733_),
    .X(_05736_));
 sky130_fd_sc_hd__and3_1 _16092_ (.A(_05730_),
    .B(_05733_),
    .C(_05734_),
    .X(_05737_));
 sky130_fd_sc_hd__nand4_2 _16093_ (.A(_05366_),
    .B(_05373_),
    .C(_05730_),
    .D(_05733_),
    .Y(_05738_));
 sky130_fd_sc_hd__a221oi_2 _16094_ (.A1(_05353_),
    .A2(_05368_),
    .B1(_05730_),
    .B2(_05733_),
    .C1(_05367_),
    .Y(_05739_));
 sky130_fd_sc_hd__a31oi_4 _16095_ (.A1(_05693_),
    .A2(_05726_),
    .A3(_05727_),
    .B1(_05734_),
    .Y(_05740_));
 sky130_fd_sc_hd__a311oi_2 _16096_ (.A1(_05693_),
    .A2(_05726_),
    .A3(_05727_),
    .B1(_05731_),
    .C1(_05734_),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(_05736_),
    .B(_05738_),
    .Y(_05742_));
 sky130_fd_sc_hd__a32oi_4 _16098_ (.A1(_05683_),
    .A2(_05684_),
    .A3(_05689_),
    .B1(_05736_),
    .B2(_05738_),
    .Y(_05744_));
 sky130_fd_sc_hd__o211a_4 _16099_ (.A1(_05735_),
    .A2(_05737_),
    .B1(_05691_),
    .C1(_05692_),
    .X(_05745_));
 sky130_fd_sc_hd__o211ai_4 _16100_ (.A1(_05735_),
    .A2(_05737_),
    .B1(_05691_),
    .C1(_05692_),
    .Y(_05746_));
 sky130_fd_sc_hd__a21oi_1 _16101_ (.A1(_05691_),
    .A2(_05692_),
    .B1(_05742_),
    .Y(_05747_));
 sky130_fd_sc_hd__o2bb2ai_4 _16102_ (.A1_N(_05691_),
    .A2_N(_05692_),
    .B1(_05739_),
    .B2(_05741_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand3_4 _16103_ (.A(_05343_),
    .B(_05615_),
    .C(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__nand4_4 _16104_ (.A(_05343_),
    .B(_05615_),
    .C(_05746_),
    .D(_05748_),
    .Y(_05750_));
 sky130_fd_sc_hd__a22oi_4 _16105_ (.A1(_05343_),
    .A2(_05615_),
    .B1(_05746_),
    .B2(_05748_),
    .Y(_05751_));
 sky130_fd_sc_hd__o22ai_4 _16106_ (.A1(_05342_),
    .A2(_05614_),
    .B1(_05745_),
    .B2(_05747_),
    .Y(_05752_));
 sky130_fd_sc_hd__a31oi_4 _16107_ (.A1(_05345_),
    .A2(_05373_),
    .A3(_05374_),
    .B1(_05380_),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2_1 _16108_ (.A(net30),
    .B(net48),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(net32),
    .B(net47),
    .Y(_05756_));
 sky130_fd_sc_hd__nand4_4 _16110_ (.A(net31),
    .B(net32),
    .C(net46),
    .D(net47),
    .Y(_05757_));
 sky130_fd_sc_hd__a22oi_1 _16111_ (.A1(net32),
    .A2(net46),
    .B1(net47),
    .B2(net31),
    .Y(_05758_));
 sky130_fd_sc_hd__a22o_1 _16112_ (.A1(net32),
    .A2(net46),
    .B1(net47),
    .B2(net31),
    .X(_05759_));
 sky130_fd_sc_hd__a22o_1 _16113_ (.A1(net30),
    .A2(net48),
    .B1(_05757_),
    .B2(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__nand4_2 _16114_ (.A(_05759_),
    .B(net48),
    .C(net30),
    .D(_05757_),
    .Y(_05761_));
 sky130_fd_sc_hd__nand2_2 _16115_ (.A(_05760_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__o21ai_4 _16116_ (.A1(_05431_),
    .A2(_05433_),
    .B1(_05437_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2_4 _16117_ (.A(net4),
    .B(net43),
    .Y(_05764_));
 sky130_fd_sc_hd__and4_1 _16118_ (.A(net3),
    .B(net4),
    .C(net42),
    .D(net43),
    .X(_05766_));
 sky130_fd_sc_hd__nand4_1 _16119_ (.A(net3),
    .B(net4),
    .C(net42),
    .D(net43),
    .Y(_05767_));
 sky130_fd_sc_hd__a22o_2 _16120_ (.A1(net4),
    .A2(net42),
    .B1(net43),
    .B2(net3),
    .X(_05768_));
 sky130_fd_sc_hd__a22oi_1 _16121_ (.A1(net2),
    .A2(net45),
    .B1(_05767_),
    .B2(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__o2bb2ai_2 _16122_ (.A1_N(_05767_),
    .A2_N(_05768_),
    .B1(_01901_),
    .B2(_02054_),
    .Y(_05770_));
 sky130_fd_sc_hd__o2111a_1 _16123_ (.A1(_05432_),
    .A2(_05764_),
    .B1(net2),
    .C1(net45),
    .D1(_05768_),
    .X(_05771_));
 sky130_fd_sc_hd__o2111ai_4 _16124_ (.A1(_05432_),
    .A2(_05764_),
    .B1(net2),
    .C1(net45),
    .D1(_05768_),
    .Y(_05772_));
 sky130_fd_sc_hd__nand3_4 _16125_ (.A(_05770_),
    .B(_05772_),
    .C(_05763_),
    .Y(_05773_));
 sky130_fd_sc_hd__a21oi_1 _16126_ (.A1(_05770_),
    .A2(_05772_),
    .B1(_05763_),
    .Y(_05774_));
 sky130_fd_sc_hd__o21bai_2 _16127_ (.A1(_05769_),
    .A2(_05771_),
    .B1_N(_05763_),
    .Y(_05775_));
 sky130_fd_sc_hd__a21oi_2 _16128_ (.A1(_05773_),
    .A2(_05775_),
    .B1(_05762_),
    .Y(_05777_));
 sky130_fd_sc_hd__and3_1 _16129_ (.A(_05775_),
    .B(_05762_),
    .C(_05773_),
    .X(_05778_));
 sky130_fd_sc_hd__nand4_2 _16130_ (.A(_05760_),
    .B(_05761_),
    .C(_05773_),
    .D(_05775_),
    .Y(_05779_));
 sky130_fd_sc_hd__a22o_1 _16131_ (.A1(_05760_),
    .A2(_05761_),
    .B1(_05773_),
    .B2(_05775_),
    .X(_05780_));
 sky130_fd_sc_hd__a21boi_1 _16132_ (.A1(_05413_),
    .A2(_05418_),
    .B1_N(_05416_),
    .Y(_05781_));
 sky130_fd_sc_hd__o21a_1 _16133_ (.A1(_01945_),
    .A2(_02010_),
    .B1(_05408_),
    .X(_05782_));
 sky130_fd_sc_hd__and3_1 _16134_ (.A(_05406_),
    .B(net41),
    .C(net4),
    .X(_05783_));
 sky130_fd_sc_hd__a31o_1 _16135_ (.A1(_05406_),
    .A2(net41),
    .A3(net4),
    .B1(_05407_),
    .X(_05784_));
 sky130_fd_sc_hd__o31a_1 _16136_ (.A1(_01945_),
    .A2(_02010_),
    .A3(_05405_),
    .B1(_05408_),
    .X(_05785_));
 sky130_fd_sc_hd__a21boi_1 _16137_ (.A1(net38),
    .A2(net7),
    .B1_N(_05350_),
    .Y(_05786_));
 sky130_fd_sc_hd__nor2_1 _16138_ (.A(_05346_),
    .B(_05347_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21a_1 _16139_ (.A1(_05346_),
    .A2(_05347_),
    .B1(_05350_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _16140_ (.A(net5),
    .B(net41),
    .Y(_05790_));
 sky130_fd_sc_hd__a22oi_4 _16141_ (.A1(net7),
    .A2(net39),
    .B1(net40),
    .B2(net6),
    .Y(_05791_));
 sky130_fd_sc_hd__a22o_1 _16142_ (.A1(net7),
    .A2(net39),
    .B1(net40),
    .B2(net6),
    .X(_05792_));
 sky130_fd_sc_hd__nand2_2 _16143_ (.A(net7),
    .B(net40),
    .Y(_05793_));
 sky130_fd_sc_hd__and4_2 _16144_ (.A(net6),
    .B(net7),
    .C(net39),
    .D(net40),
    .X(_05794_));
 sky130_fd_sc_hd__nand4_2 _16145_ (.A(net6),
    .B(net7),
    .C(net39),
    .D(net40),
    .Y(_05795_));
 sky130_fd_sc_hd__o211ai_2 _16146_ (.A1(_01956_),
    .A2(_02010_),
    .B1(_05792_),
    .C1(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__o21bai_2 _16147_ (.A1(_05791_),
    .A2(_05794_),
    .B1_N(_05790_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand4_2 _16148_ (.A(_05792_),
    .B(_05795_),
    .C(net5),
    .D(net41),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ai_2 _16149_ (.A1(_05791_),
    .A2(_05794_),
    .B1(_05790_),
    .Y(_05800_));
 sky130_fd_sc_hd__a2bb2oi_2 _16150_ (.A1_N(_05349_),
    .A2_N(_05788_),
    .B1(_05796_),
    .B2(_05797_),
    .Y(_05801_));
 sky130_fd_sc_hd__o211ai_4 _16151_ (.A1(_05349_),
    .A2(_05788_),
    .B1(_05799_),
    .C1(_05800_),
    .Y(_05802_));
 sky130_fd_sc_hd__a2bb2oi_2 _16152_ (.A1_N(_05347_),
    .A2_N(_05786_),
    .B1(_05799_),
    .B2(_05800_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand3_2 _16153_ (.A(_05789_),
    .B(_05796_),
    .C(_05797_),
    .Y(_05804_));
 sky130_fd_sc_hd__o211ai_2 _16154_ (.A1(_05407_),
    .A2(_05783_),
    .B1(_05802_),
    .C1(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__o22ai_2 _16155_ (.A1(_05405_),
    .A2(_05782_),
    .B1(_05801_),
    .B2(_05803_),
    .Y(_05806_));
 sky130_fd_sc_hd__o2111ai_4 _16156_ (.A1(_05404_),
    .A2(_05405_),
    .B1(_05408_),
    .C1(_05802_),
    .D1(_05804_),
    .Y(_05807_));
 sky130_fd_sc_hd__o22ai_2 _16157_ (.A1(_05407_),
    .A2(_05783_),
    .B1(_05801_),
    .B2(_05803_),
    .Y(_05808_));
 sky130_fd_sc_hd__o211a_1 _16158_ (.A1(_05415_),
    .A2(_05421_),
    .B1(_05805_),
    .C1(_05806_),
    .X(_05810_));
 sky130_fd_sc_hd__o211ai_4 _16159_ (.A1(_05415_),
    .A2(_05421_),
    .B1(_05805_),
    .C1(_05806_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand3_4 _16160_ (.A(_05808_),
    .B(_05781_),
    .C(_05807_),
    .Y(_05812_));
 sky130_fd_sc_hd__o21a_1 _16161_ (.A1(_05777_),
    .A2(_05778_),
    .B1(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__o211a_1 _16162_ (.A1(_05777_),
    .A2(_05778_),
    .B1(_05811_),
    .C1(_05812_),
    .X(_05814_));
 sky130_fd_sc_hd__o211ai_4 _16163_ (.A1(_05777_),
    .A2(_05778_),
    .B1(_05811_),
    .C1(_05812_),
    .Y(_05815_));
 sky130_fd_sc_hd__a22oi_2 _16164_ (.A1(_05779_),
    .A2(_05780_),
    .B1(_05811_),
    .B2(_05812_),
    .Y(_05816_));
 sky130_fd_sc_hd__a22o_1 _16165_ (.A1(_05779_),
    .A2(_05780_),
    .B1(_05811_),
    .B2(_05812_),
    .X(_05817_));
 sky130_fd_sc_hd__a2bb2oi_2 _16166_ (.A1_N(_05377_),
    .A2_N(_05753_),
    .B1(_05815_),
    .B2(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__o22ai_4 _16167_ (.A1(_05377_),
    .A2(_05753_),
    .B1(_05814_),
    .B2(_05816_),
    .Y(_05819_));
 sky130_fd_sc_hd__o211a_1 _16168_ (.A1(_05375_),
    .A2(_05386_),
    .B1(_05815_),
    .C1(_05817_),
    .X(_05821_));
 sky130_fd_sc_hd__o211ai_4 _16169_ (.A1(_05375_),
    .A2(_05386_),
    .B1(_05815_),
    .C1(_05817_),
    .Y(_05822_));
 sky130_fd_sc_hd__a21oi_1 _16170_ (.A1(_05454_),
    .A2(_05455_),
    .B1(_05427_),
    .Y(_05823_));
 sky130_fd_sc_hd__o21ai_1 _16171_ (.A1(_05424_),
    .A2(_05456_),
    .B1(_05428_),
    .Y(_05824_));
 sky130_fd_sc_hd__o21ai_2 _16172_ (.A1(_05427_),
    .A2(_05459_),
    .B1(_05819_),
    .Y(_05825_));
 sky130_fd_sc_hd__and3_2 _16173_ (.A(_05819_),
    .B(_05822_),
    .C(_05824_),
    .X(_05826_));
 sky130_fd_sc_hd__o22a_2 _16174_ (.A1(_05818_),
    .A2(_05821_),
    .B1(_05823_),
    .B2(_05424_),
    .X(_05827_));
 sky130_fd_sc_hd__o2bb2ai_1 _16175_ (.A1_N(_05819_),
    .A2_N(_05822_),
    .B1(_05823_),
    .B2(_05424_),
    .Y(_05828_));
 sky130_fd_sc_hd__o211a_1 _16176_ (.A1(_05424_),
    .A2(_05823_),
    .B1(_05822_),
    .C1(_05819_),
    .X(_05829_));
 sky130_fd_sc_hd__o2111ai_1 _16177_ (.A1(_05424_),
    .A2(_05456_),
    .B1(_05819_),
    .C1(_05822_),
    .D1(_05428_),
    .Y(_05830_));
 sky130_fd_sc_hd__o22a_2 _16178_ (.A1(_05427_),
    .A2(_05459_),
    .B1(_05818_),
    .B2(_05821_),
    .X(_05832_));
 sky130_fd_sc_hd__o22ai_1 _16179_ (.A1(_05427_),
    .A2(_05459_),
    .B1(_05818_),
    .B2(_05821_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_1 _16180_ (.A(_05830_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__o21ai_1 _16181_ (.A1(_05821_),
    .A2(_05825_),
    .B1(_05828_),
    .Y(_05835_));
 sky130_fd_sc_hd__o221ai_4 _16182_ (.A1(_05826_),
    .A2(_05827_),
    .B1(_05745_),
    .B2(_05749_),
    .C1(_05752_),
    .Y(_05836_));
 sky130_fd_sc_hd__o2bb2ai_1 _16183_ (.A1_N(_05750_),
    .A2_N(_05752_),
    .B1(_05829_),
    .B2(_05832_),
    .Y(_05837_));
 sky130_fd_sc_hd__o2bb2ai_4 _16184_ (.A1_N(_05750_),
    .A2_N(_05752_),
    .B1(_05826_),
    .B2(_05827_),
    .Y(_05838_));
 sky130_fd_sc_hd__o21ai_2 _16185_ (.A1(_05829_),
    .A2(_05832_),
    .B1(_05750_),
    .Y(_05839_));
 sky130_fd_sc_hd__o211ai_4 _16186_ (.A1(_05829_),
    .A2(_05832_),
    .B1(_05750_),
    .C1(_05752_),
    .Y(_05840_));
 sky130_fd_sc_hd__a22oi_4 _16187_ (.A1(_05396_),
    .A2(_05612_),
    .B1(_05838_),
    .B2(_05840_),
    .Y(_05841_));
 sky130_fd_sc_hd__o211ai_4 _16188_ (.A1(_05395_),
    .A2(_05610_),
    .B1(_05836_),
    .C1(_05837_),
    .Y(_05843_));
 sky130_fd_sc_hd__o211a_2 _16189_ (.A1(_05751_),
    .A2(_05839_),
    .B1(_05613_),
    .C1(_05838_),
    .X(_05844_));
 sky130_fd_sc_hd__o211ai_4 _16190_ (.A1(_05751_),
    .A2(_05839_),
    .B1(_05613_),
    .C1(_05838_),
    .Y(_05845_));
 sky130_fd_sc_hd__nand3_2 _16191_ (.A(_05609_),
    .B(_05843_),
    .C(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__o22ai_4 _16192_ (.A1(_05607_),
    .A2(_05608_),
    .B1(_05841_),
    .B2(_05844_),
    .Y(_05847_));
 sky130_fd_sc_hd__o211ai_2 _16193_ (.A1(_05604_),
    .A2(_05596_),
    .B1(_05602_),
    .C1(_05843_),
    .Y(_05848_));
 sky130_fd_sc_hd__nand4_1 _16194_ (.A(_05602_),
    .B(_05606_),
    .C(_05843_),
    .D(_05845_),
    .Y(_05849_));
 sky130_fd_sc_hd__o22ai_2 _16195_ (.A1(_05601_),
    .A2(_05605_),
    .B1(_05841_),
    .B2(_05844_),
    .Y(_05850_));
 sky130_fd_sc_hd__o221a_2 _16196_ (.A1(_05844_),
    .A2(_05848_),
    .B1(_05487_),
    .B2(_05492_),
    .C1(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__o211ai_2 _16197_ (.A1(_05487_),
    .A2(_05492_),
    .B1(_05849_),
    .C1(_05850_),
    .Y(_05852_));
 sky130_fd_sc_hd__nand3_1 _16198_ (.A(_05847_),
    .B(_05518_),
    .C(_05846_),
    .Y(_05854_));
 sky130_fd_sc_hd__a21o_1 _16199_ (.A1(_05234_),
    .A2(_05241_),
    .B1(_05235_),
    .X(_05855_));
 sky130_fd_sc_hd__inv_2 _16200_ (.A(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__o2111ai_1 _16201_ (.A1(_05233_),
    .A2(_05240_),
    .B1(_05852_),
    .C1(_05854_),
    .D1(_05236_),
    .Y(_05857_));
 sky130_fd_sc_hd__a22o_1 _16202_ (.A1(_05236_),
    .A2(_05247_),
    .B1(_05852_),
    .B2(_05854_),
    .X(_05858_));
 sky130_fd_sc_hd__a22o_1 _16203_ (.A1(_05234_),
    .A2(_05243_),
    .B1(_05852_),
    .B2(_05854_),
    .X(_05859_));
 sky130_fd_sc_hd__a31oi_4 _16204_ (.A1(_05847_),
    .A2(_05518_),
    .A3(_05846_),
    .B1(_05856_),
    .Y(_05860_));
 sky130_fd_sc_hd__a31o_1 _16205_ (.A1(_05847_),
    .A2(_05518_),
    .A3(_05846_),
    .B1(_05856_),
    .X(_05861_));
 sky130_fd_sc_hd__o21ai_1 _16206_ (.A1(_05851_),
    .A2(_05861_),
    .B1(_05859_),
    .Y(_05862_));
 sky130_fd_sc_hd__o211ai_1 _16207_ (.A1(_05497_),
    .A2(_05515_),
    .B1(_05857_),
    .C1(_05858_),
    .Y(_05863_));
 sky130_fd_sc_hd__o211ai_4 _16208_ (.A1(_05851_),
    .A2(_05861_),
    .B1(_05859_),
    .C1(_05516_),
    .Y(_05865_));
 sky130_fd_sc_hd__inv_2 _16209_ (.A(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__a22oi_1 _16210_ (.A1(_05505_),
    .A2(_05503_),
    .B1(_05865_),
    .B2(_05863_),
    .Y(_05867_));
 sky130_fd_sc_hd__a21oi_1 _16211_ (.A1(_05862_),
    .A2(_05517_),
    .B1(_05506_),
    .Y(_05868_));
 sky130_fd_sc_hd__and4_1 _16212_ (.A(_05503_),
    .B(_05865_),
    .C(_05505_),
    .D(_05863_),
    .X(_05869_));
 sky130_fd_sc_hd__a21oi_2 _16213_ (.A1(_05868_),
    .A2(_05865_),
    .B1(_05867_),
    .Y(_05870_));
 sky130_fd_sc_hd__a21oi_1 _16214_ (.A1(_05158_),
    .A2(_05160_),
    .B1(_05508_),
    .Y(_05871_));
 sky130_fd_sc_hd__a31o_1 _16215_ (.A1(_05165_),
    .A2(_05511_),
    .A3(_05161_),
    .B1(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__xor2_1 _16216_ (.A(_05870_),
    .B(_05872_),
    .X(net88));
 sky130_fd_sc_hd__a32o_1 _16217_ (.A1(_05518_),
    .A2(_05846_),
    .A3(_05847_),
    .B1(_05852_),
    .B2(_05856_),
    .X(_05873_));
 sky130_fd_sc_hd__and3_1 _16218_ (.A(_05213_),
    .B(_05232_),
    .C(_05597_),
    .X(_05875_));
 sky130_fd_sc_hd__a31o_1 _16219_ (.A1(_05587_),
    .A2(_05591_),
    .A3(_05593_),
    .B1(_05603_),
    .X(_05876_));
 sky130_fd_sc_hd__a31o_1 _16220_ (.A1(_05213_),
    .A2(_05232_),
    .A3(_05597_),
    .B1(_05594_),
    .X(_05877_));
 sky130_fd_sc_hd__a32oi_4 _16221_ (.A1(_05613_),
    .A2(_05838_),
    .A3(_05840_),
    .B1(_05606_),
    .B2(_05602_),
    .Y(_05878_));
 sky130_fd_sc_hd__a31o_1 _16222_ (.A1(_05602_),
    .A2(_05606_),
    .A3(_05843_),
    .B1(_05844_),
    .X(_05879_));
 sky130_fd_sc_hd__o31a_2 _16223_ (.A1(_05535_),
    .A2(_05537_),
    .A3(_05583_),
    .B1(_05586_),
    .X(_05880_));
 sky130_fd_sc_hd__o211a_1 _16224_ (.A1(_05424_),
    .A2(_05456_),
    .B1(_05822_),
    .C1(_05428_),
    .X(_05881_));
 sky130_fd_sc_hd__a21o_2 _16225_ (.A1(_05819_),
    .A2(_05824_),
    .B1(_05821_),
    .X(_05882_));
 sky130_fd_sc_hd__a22o_1 _16226_ (.A1(net23),
    .A2(net54),
    .B1(net56),
    .B2(net12),
    .X(_05883_));
 sky130_fd_sc_hd__nand2_2 _16227_ (.A(net23),
    .B(net56),
    .Y(_05884_));
 sky130_fd_sc_hd__nand4_1 _16228_ (.A(net23),
    .B(net12),
    .C(net54),
    .D(net56),
    .Y(_05886_));
 sky130_fd_sc_hd__a22o_1 _16229_ (.A1(_01846_),
    .A2(net57),
    .B1(_05883_),
    .B2(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__o2111ai_4 _16230_ (.A1(_05519_),
    .A2(_05884_),
    .B1(net57),
    .C1(_05883_),
    .D1(_01846_),
    .Y(_05888_));
 sky130_fd_sc_hd__nand2_1 _16231_ (.A(_05887_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__o21ai_4 _16232_ (.A1(_05519_),
    .A2(_05524_),
    .B1(_05522_),
    .Y(_05890_));
 sky130_fd_sc_hd__a22oi_4 _16233_ (.A1(net28),
    .A2(net51),
    .B1(net52),
    .B2(net27),
    .Y(_05891_));
 sky130_fd_sc_hd__and4_1 _16234_ (.A(net28),
    .B(net27),
    .C(net51),
    .D(net52),
    .X(_05892_));
 sky130_fd_sc_hd__nand4_1 _16235_ (.A(net28),
    .B(net27),
    .C(net51),
    .D(net52),
    .Y(_05893_));
 sky130_fd_sc_hd__o21ai_2 _16236_ (.A1(_05891_),
    .A2(_05892_),
    .B1(_05520_),
    .Y(_05894_));
 sky130_fd_sc_hd__a41o_1 _16237_ (.A1(net28),
    .A2(net27),
    .A3(net51),
    .A4(net52),
    .B1(_05520_),
    .X(_05895_));
 sky130_fd_sc_hd__nand4b_1 _16238_ (.A_N(_05891_),
    .B(_05893_),
    .C(net26),
    .D(net53),
    .Y(_05897_));
 sky130_fd_sc_hd__a21oi_2 _16239_ (.A1(_05894_),
    .A2(_05897_),
    .B1(_05890_),
    .Y(_05898_));
 sky130_fd_sc_hd__a21o_1 _16240_ (.A1(_05894_),
    .A2(_05897_),
    .B1(_05890_),
    .X(_05899_));
 sky130_fd_sc_hd__o211a_1 _16241_ (.A1(_05891_),
    .A2(_05895_),
    .B1(_05890_),
    .C1(_05894_),
    .X(_05900_));
 sky130_fd_sc_hd__o211ai_4 _16242_ (.A1(_05891_),
    .A2(_05895_),
    .B1(_05890_),
    .C1(_05894_),
    .Y(_05901_));
 sky130_fd_sc_hd__nand4_4 _16243_ (.A(_05887_),
    .B(_05888_),
    .C(_05899_),
    .D(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__o2bb2a_1 _16244_ (.A1_N(_05887_),
    .A2_N(_05888_),
    .B1(_05898_),
    .B2(_05900_),
    .X(_05903_));
 sky130_fd_sc_hd__o21ai_2 _16245_ (.A1(_05898_),
    .A2(_05900_),
    .B1(_05889_),
    .Y(_05904_));
 sky130_fd_sc_hd__a311oi_4 _16246_ (.A1(_05527_),
    .A2(_05218_),
    .A3(_05215_),
    .B1(_01846_),
    .C1(_02229_),
    .Y(_05905_));
 sky130_fd_sc_hd__a211o_2 _16247_ (.A1(_05902_),
    .A2(_05904_),
    .B1(_05905_),
    .C1(_05528_),
    .X(_05906_));
 sky130_fd_sc_hd__o21ai_2 _16248_ (.A1(_05528_),
    .A2(_05905_),
    .B1(_05902_),
    .Y(_05908_));
 sky130_fd_sc_hd__o211a_1 _16249_ (.A1(_05528_),
    .A2(_05905_),
    .B1(_05904_),
    .C1(_05902_),
    .X(_05909_));
 sky130_fd_sc_hd__o211ai_4 _16250_ (.A1(_05528_),
    .A2(_05905_),
    .B1(_05904_),
    .C1(_05902_),
    .Y(_05910_));
 sky130_fd_sc_hd__o21ai_1 _16251_ (.A1(_05903_),
    .A2(_05908_),
    .B1(_05906_),
    .Y(_05911_));
 sky130_fd_sc_hd__o21ai_1 _16252_ (.A1(_05755_),
    .A2(_05758_),
    .B1(_05757_),
    .Y(_05912_));
 sky130_fd_sc_hd__o21a_1 _16253_ (.A1(_05755_),
    .A2(_05758_),
    .B1(_05757_),
    .X(_05913_));
 sky130_fd_sc_hd__a22oi_4 _16254_ (.A1(net31),
    .A2(net48),
    .B1(net49),
    .B2(net30),
    .Y(_05914_));
 sky130_fd_sc_hd__a22o_1 _16255_ (.A1(net31),
    .A2(net48),
    .B1(net49),
    .B2(net30),
    .X(_05915_));
 sky130_fd_sc_hd__and4_1 _16256_ (.A(net30),
    .B(net31),
    .C(net48),
    .D(net49),
    .X(_05916_));
 sky130_fd_sc_hd__nand4_2 _16257_ (.A(net30),
    .B(net31),
    .C(net48),
    .D(net49),
    .Y(_05917_));
 sky130_fd_sc_hd__nand3_1 _16258_ (.A(_05552_),
    .B(_05915_),
    .C(_05917_),
    .Y(_05919_));
 sky130_fd_sc_hd__o21bai_2 _16259_ (.A1(_05914_),
    .A2(_05916_),
    .B1_N(_05552_),
    .Y(_05920_));
 sky130_fd_sc_hd__a22o_1 _16260_ (.A1(net29),
    .A2(net50),
    .B1(_05915_),
    .B2(_05917_),
    .X(_05921_));
 sky130_fd_sc_hd__nand4_1 _16261_ (.A(_05915_),
    .B(_05917_),
    .C(net29),
    .D(net50),
    .Y(_05922_));
 sky130_fd_sc_hd__nand3_4 _16262_ (.A(_05913_),
    .B(_05919_),
    .C(_05920_),
    .Y(_05923_));
 sky130_fd_sc_hd__and3_2 _16263_ (.A(_05921_),
    .B(_05922_),
    .C(_05912_),
    .X(_05924_));
 sky130_fd_sc_hd__nand3_2 _16264_ (.A(_05921_),
    .B(_05922_),
    .C(_05912_),
    .Y(_05925_));
 sky130_fd_sc_hd__o32a_1 _16265_ (.A1(_01748_),
    .A2(_02120_),
    .A3(_05552_),
    .B1(_02152_),
    .B2(_01769_),
    .X(_05926_));
 sky130_fd_sc_hd__a31o_1 _16266_ (.A1(_05551_),
    .A2(net51),
    .A3(net27),
    .B1(_05553_),
    .X(_05927_));
 sky130_fd_sc_hd__o2bb2ai_4 _16267_ (.A1_N(_05923_),
    .A2_N(_05925_),
    .B1(_05926_),
    .B2(_05550_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _16268_ (.A(_05923_),
    .B(_05927_),
    .Y(_05930_));
 sky130_fd_sc_hd__and3_1 _16269_ (.A(_05923_),
    .B(_05925_),
    .C(_05927_),
    .X(_05931_));
 sky130_fd_sc_hd__nand3_1 _16270_ (.A(_05923_),
    .B(_05925_),
    .C(_05927_),
    .Y(_05932_));
 sky130_fd_sc_hd__o21ai_4 _16271_ (.A1(_05762_),
    .A2(_05774_),
    .B1(_05773_),
    .Y(_05933_));
 sky130_fd_sc_hd__a21oi_2 _16272_ (.A1(_05928_),
    .A2(_05932_),
    .B1(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__a21o_1 _16273_ (.A1(_05928_),
    .A2(_05932_),
    .B1(_05933_),
    .X(_05935_));
 sky130_fd_sc_hd__o211a_1 _16274_ (.A1(_05930_),
    .A2(_05924_),
    .B1(_05928_),
    .C1(_05933_),
    .X(_05936_));
 sky130_fd_sc_hd__o211ai_4 _16275_ (.A1(_05930_),
    .A2(_05924_),
    .B1(_05928_),
    .C1(_05933_),
    .Y(_05937_));
 sky130_fd_sc_hd__o31a_2 _16276_ (.A1(_05184_),
    .A2(_05542_),
    .A3(_05561_),
    .B1(_05560_),
    .X(_05938_));
 sky130_fd_sc_hd__a32o_1 _16277_ (.A1(_05547_),
    .A2(_05557_),
    .A3(_05558_),
    .B1(_05562_),
    .B2(_05544_),
    .X(_05939_));
 sky130_fd_sc_hd__o21ai_2 _16278_ (.A1(_05934_),
    .A2(_05936_),
    .B1(_05938_),
    .Y(_05941_));
 sky130_fd_sc_hd__nand3_2 _16279_ (.A(_05935_),
    .B(_05937_),
    .C(_05939_),
    .Y(_05942_));
 sky130_fd_sc_hd__o2bb2ai_2 _16280_ (.A1_N(_05560_),
    .A2_N(_05563_),
    .B1(_05934_),
    .B2(_05936_),
    .Y(_05943_));
 sky130_fd_sc_hd__nand3_2 _16281_ (.A(_05935_),
    .B(_05937_),
    .C(_05938_),
    .Y(_05944_));
 sky130_fd_sc_hd__a31oi_2 _16282_ (.A1(_05541_),
    .A2(_05565_),
    .A3(_05568_),
    .B1(_05575_),
    .Y(_05945_));
 sky130_fd_sc_hd__o22ai_2 _16283_ (.A1(_05564_),
    .A2(_05571_),
    .B1(_05576_),
    .B2(_05569_),
    .Y(_05946_));
 sky130_fd_sc_hd__and3_1 _16284_ (.A(_05941_),
    .B(_05946_),
    .C(_05942_),
    .X(_05947_));
 sky130_fd_sc_hd__nand3_4 _16285_ (.A(_05941_),
    .B(_05946_),
    .C(_05942_),
    .Y(_05948_));
 sky130_fd_sc_hd__o211ai_4 _16286_ (.A1(_05569_),
    .A2(_05945_),
    .B1(_05944_),
    .C1(_05943_),
    .Y(_05949_));
 sky130_fd_sc_hd__a41oi_4 _16287_ (.A1(_05573_),
    .A2(_05579_),
    .A3(_05943_),
    .A4(_05944_),
    .B1(_05911_),
    .Y(_05950_));
 sky130_fd_sc_hd__o2111a_2 _16288_ (.A1(_05908_),
    .A2(_05903_),
    .B1(_05906_),
    .C1(_05948_),
    .D1(_05949_),
    .X(_05952_));
 sky130_fd_sc_hd__nand2_2 _16289_ (.A(_05950_),
    .B(_05948_),
    .Y(_05953_));
 sky130_fd_sc_hd__a22oi_4 _16290_ (.A1(_05906_),
    .A2(_05910_),
    .B1(_05948_),
    .B2(_05949_),
    .Y(_05954_));
 sky130_fd_sc_hd__a22o_2 _16291_ (.A1(_05906_),
    .A2(_05910_),
    .B1(_05948_),
    .B2(_05949_),
    .X(_05955_));
 sky130_fd_sc_hd__a221oi_4 _16292_ (.A1(_05950_),
    .A2(_05948_),
    .B1(_05825_),
    .B2(_05822_),
    .C1(_05954_),
    .Y(_05956_));
 sky130_fd_sc_hd__nand3_4 _16293_ (.A(_05882_),
    .B(_05953_),
    .C(_05955_),
    .Y(_05957_));
 sky130_fd_sc_hd__a21oi_4 _16294_ (.A1(_05953_),
    .A2(_05955_),
    .B1(_05882_),
    .Y(_05958_));
 sky130_fd_sc_hd__o22ai_4 _16295_ (.A1(_05818_),
    .A2(_05881_),
    .B1(_05952_),
    .B2(_05954_),
    .Y(_05959_));
 sky130_fd_sc_hd__o21ai_1 _16296_ (.A1(_05585_),
    .A2(_05588_),
    .B1(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__inv_2 _16297_ (.A(_05960_),
    .Y(_05961_));
 sky130_fd_sc_hd__o211a_1 _16298_ (.A1(_05585_),
    .A2(_05588_),
    .B1(_05957_),
    .C1(_05959_),
    .X(_05963_));
 sky130_fd_sc_hd__a21boi_1 _16299_ (.A1(_05957_),
    .A2(_05959_),
    .B1_N(_05880_),
    .Y(_05964_));
 sky130_fd_sc_hd__o21ai_1 _16300_ (.A1(_05956_),
    .A2(_05958_),
    .B1(_05880_),
    .Y(_05965_));
 sky130_fd_sc_hd__a21oi_1 _16301_ (.A1(_05957_),
    .A2(_05959_),
    .B1(_05880_),
    .Y(_05966_));
 sky130_fd_sc_hd__o22ai_4 _16302_ (.A1(_05585_),
    .A2(_05588_),
    .B1(_05956_),
    .B2(_05958_),
    .Y(_05967_));
 sky130_fd_sc_hd__and3_1 _16303_ (.A(_05957_),
    .B(_05959_),
    .C(_05880_),
    .X(_05968_));
 sky130_fd_sc_hd__nand3_2 _16304_ (.A(_05959_),
    .B(_05880_),
    .C(_05957_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2_1 _16305_ (.A(_05967_),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__o21ai_1 _16306_ (.A1(_05956_),
    .A2(_05960_),
    .B1(_05965_),
    .Y(_05971_));
 sky130_fd_sc_hd__a32oi_4 _16307_ (.A1(_05685_),
    .A2(_05687_),
    .A3(_05686_),
    .B1(_05742_),
    .B2(_05692_),
    .Y(_05972_));
 sky130_fd_sc_hd__o21ai_2 _16308_ (.A1(_05653_),
    .A2(_05654_),
    .B1(_05659_),
    .Y(_05974_));
 sky130_fd_sc_hd__a22oi_4 _16309_ (.A1(net61),
    .A2(net18),
    .B1(net19),
    .B2(net60),
    .Y(_05975_));
 sky130_fd_sc_hd__a22o_1 _16310_ (.A1(net61),
    .A2(net18),
    .B1(net19),
    .B2(net60),
    .X(_05976_));
 sky130_fd_sc_hd__and4_2 _16311_ (.A(net60),
    .B(net61),
    .C(net18),
    .D(net19),
    .X(_05977_));
 sky130_fd_sc_hd__nand4_1 _16312_ (.A(net60),
    .B(net61),
    .C(net18),
    .D(net19),
    .Y(_05978_));
 sky130_fd_sc_hd__nand3_1 _16313_ (.A(_05621_),
    .B(_05976_),
    .C(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21bai_2 _16314_ (.A1(_05975_),
    .A2(_05977_),
    .B1_N(_05621_),
    .Y(_05980_));
 sky130_fd_sc_hd__o21ai_1 _16315_ (.A1(_05975_),
    .A2(_05977_),
    .B1(_05621_),
    .Y(_05981_));
 sky130_fd_sc_hd__nand4_1 _16316_ (.A(_05976_),
    .B(_05978_),
    .C(net62),
    .D(net17),
    .Y(_05982_));
 sky130_fd_sc_hd__a21oi_1 _16317_ (.A1(_05981_),
    .A2(_05982_),
    .B1(_05974_),
    .Y(_05983_));
 sky130_fd_sc_hd__nand3b_4 _16318_ (.A_N(_05974_),
    .B(_05979_),
    .C(_05980_),
    .Y(_05985_));
 sky130_fd_sc_hd__nand3_2 _16319_ (.A(_05981_),
    .B(_05982_),
    .C(_05974_),
    .Y(_05986_));
 sky130_fd_sc_hd__a31o_1 _16320_ (.A1(_05620_),
    .A2(net15),
    .A3(net63),
    .B1(_05623_),
    .X(_05987_));
 sky130_fd_sc_hd__o32a_2 _16321_ (.A1(_01890_),
    .A2(_02076_),
    .A3(_05619_),
    .B1(_05621_),
    .B2(_05265_),
    .X(_05988_));
 sky130_fd_sc_hd__a21oi_2 _16322_ (.A1(_05985_),
    .A2(_05986_),
    .B1(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__a21o_1 _16323_ (.A1(_05985_),
    .A2(_05986_),
    .B1(_05988_),
    .X(_05990_));
 sky130_fd_sc_hd__and3_1 _16324_ (.A(_05985_),
    .B(_05986_),
    .C(_05988_),
    .X(_05991_));
 sky130_fd_sc_hd__nand3_2 _16325_ (.A(_05985_),
    .B(_05986_),
    .C(_05988_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand2_2 _16326_ (.A(_05990_),
    .B(_05992_),
    .Y(_05993_));
 sky130_fd_sc_hd__a21oi_1 _16327_ (.A1(_05650_),
    .A2(_05667_),
    .B1(_05651_),
    .Y(_05994_));
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(net58),
    .B(net22),
    .Y(_05996_));
 sky130_fd_sc_hd__nand4_4 _16329_ (.A(net55),
    .B(net58),
    .C(net21),
    .D(net22),
    .Y(_05997_));
 sky130_fd_sc_hd__a22oi_4 _16330_ (.A1(net58),
    .A2(net21),
    .B1(net22),
    .B2(net55),
    .Y(_05998_));
 sky130_fd_sc_hd__a22o_2 _16331_ (.A1(net58),
    .A2(net21),
    .B1(net22),
    .B2(net55),
    .X(_05999_));
 sky130_fd_sc_hd__o221a_2 _16332_ (.A1(_01813_),
    .A2(_02163_),
    .B1(_05639_),
    .B2(_05996_),
    .C1(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__a21oi_2 _16333_ (.A1(_05997_),
    .A2(_05999_),
    .B1(_05657_),
    .Y(_06001_));
 sky130_fd_sc_hd__a22oi_4 _16334_ (.A1(net59),
    .A2(net20),
    .B1(_05997_),
    .B2(_05999_),
    .Y(_06002_));
 sky130_fd_sc_hd__o2bb2ai_1 _16335_ (.A1_N(_05997_),
    .A2_N(_05999_),
    .B1(_01813_),
    .B2(_02163_),
    .Y(_06003_));
 sky130_fd_sc_hd__a41o_1 _16336_ (.A1(net55),
    .A2(net58),
    .A3(net21),
    .A4(net22),
    .B1(_05657_),
    .X(_06004_));
 sky130_fd_sc_hd__and4_1 _16337_ (.A(_05999_),
    .B(net20),
    .C(net59),
    .D(_05997_),
    .X(_06005_));
 sky130_fd_sc_hd__o21ai_2 _16338_ (.A1(_05998_),
    .A2(_06004_),
    .B1(_06003_),
    .Y(_06007_));
 sky130_fd_sc_hd__o21ai_1 _16339_ (.A1(_05294_),
    .A2(_05642_),
    .B1(_05639_),
    .Y(_06008_));
 sky130_fd_sc_hd__nor2_1 _16340_ (.A(_05639_),
    .B(_05640_),
    .Y(_06009_));
 sky130_fd_sc_hd__o22ai_2 _16341_ (.A1(_05294_),
    .A2(_05642_),
    .B1(_05639_),
    .B2(_05640_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2_2 _16342_ (.A(net33),
    .B(net25),
    .Y(_06011_));
 sky130_fd_sc_hd__a21oi_2 _16343_ (.A1(net33),
    .A2(net25),
    .B1(net57),
    .Y(_06012_));
 sky130_fd_sc_hd__a21o_1 _16344_ (.A1(net33),
    .A2(net25),
    .B1(net57),
    .X(_06013_));
 sky130_fd_sc_hd__and3_2 _16345_ (.A(net33),
    .B(net57),
    .C(net25),
    .X(_06014_));
 sky130_fd_sc_hd__nand3_2 _16346_ (.A(net33),
    .B(net57),
    .C(net25),
    .Y(_06015_));
 sky130_fd_sc_hd__o22ai_4 _16347_ (.A1(_01759_),
    .A2(_02218_),
    .B1(_06012_),
    .B2(_06014_),
    .Y(_06016_));
 sky130_fd_sc_hd__a21oi_2 _16348_ (.A1(_02240_),
    .A2(_06011_),
    .B1(_05642_),
    .Y(_06018_));
 sky130_fd_sc_hd__nand4_4 _16349_ (.A(_06013_),
    .B(_06015_),
    .C(net44),
    .D(net24),
    .Y(_06019_));
 sky130_fd_sc_hd__o211ai_2 _16350_ (.A1(_01759_),
    .A2(_02218_),
    .B1(_06013_),
    .C1(_06015_),
    .Y(_06020_));
 sky130_fd_sc_hd__o21bai_1 _16351_ (.A1(_06012_),
    .A2(_06014_),
    .B1_N(_05642_),
    .Y(_06021_));
 sky130_fd_sc_hd__a22oi_4 _16352_ (.A1(_05641_),
    .A2(_06008_),
    .B1(_06016_),
    .B2(_06019_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand3b_2 _16353_ (.A_N(_06010_),
    .B(_06020_),
    .C(_06021_),
    .Y(_06023_));
 sky130_fd_sc_hd__a2bb2oi_2 _16354_ (.A1_N(_05643_),
    .A2_N(_06009_),
    .B1(_06020_),
    .B2(_06021_),
    .Y(_06024_));
 sky130_fd_sc_hd__nand3_4 _16355_ (.A(_06016_),
    .B(_06019_),
    .C(_06010_),
    .Y(_06025_));
 sky130_fd_sc_hd__o21ai_2 _16356_ (.A1(_06000_),
    .A2(_06001_),
    .B1(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__o21ai_2 _16357_ (.A1(_06022_),
    .A2(_06024_),
    .B1(_06007_),
    .Y(_06027_));
 sky130_fd_sc_hd__o211ai_4 _16358_ (.A1(_06002_),
    .A2(_06005_),
    .B1(_06023_),
    .C1(_06025_),
    .Y(_06029_));
 sky130_fd_sc_hd__o22ai_4 _16359_ (.A1(_06000_),
    .A2(_06001_),
    .B1(_06022_),
    .B2(_06024_),
    .Y(_06030_));
 sky130_fd_sc_hd__o221a_4 _16360_ (.A1(_06022_),
    .A2(_06026_),
    .B1(_05651_),
    .B2(_05671_),
    .C1(_06027_),
    .X(_06031_));
 sky130_fd_sc_hd__o221ai_4 _16361_ (.A1(_06022_),
    .A2(_06026_),
    .B1(_05651_),
    .B2(_05671_),
    .C1(_06027_),
    .Y(_06032_));
 sky130_fd_sc_hd__o2111ai_4 _16362_ (.A1(_05638_),
    .A2(_05649_),
    .B1(_05672_),
    .C1(_06029_),
    .D1(_06030_),
    .Y(_06033_));
 sky130_fd_sc_hd__a32oi_4 _16363_ (.A1(_05994_),
    .A2(_06029_),
    .A3(_06030_),
    .B1(_05992_),
    .B2(_05990_),
    .Y(_06034_));
 sky130_fd_sc_hd__o21ai_2 _16364_ (.A1(_05989_),
    .A2(_05991_),
    .B1(_06033_),
    .Y(_06035_));
 sky130_fd_sc_hd__o211a_2 _16365_ (.A1(_05989_),
    .A2(_05991_),
    .B1(_06032_),
    .C1(_06033_),
    .X(_06036_));
 sky130_fd_sc_hd__o211ai_2 _16366_ (.A1(_05989_),
    .A2(_05991_),
    .B1(_06032_),
    .C1(_06033_),
    .Y(_06037_));
 sky130_fd_sc_hd__a21oi_2 _16367_ (.A1(_06032_),
    .A2(_06033_),
    .B1(_05993_),
    .Y(_06038_));
 sky130_fd_sc_hd__a21o_2 _16368_ (.A1(_06032_),
    .A2(_06033_),
    .B1(_05993_),
    .X(_06040_));
 sky130_fd_sc_hd__nand2_1 _16369_ (.A(_06040_),
    .B(_05682_),
    .Y(_06041_));
 sky130_fd_sc_hd__and3_1 _16370_ (.A(_06040_),
    .B(_05682_),
    .C(_06037_),
    .X(_06042_));
 sky130_fd_sc_hd__o211ai_4 _16371_ (.A1(_06031_),
    .A2(_06035_),
    .B1(_05682_),
    .C1(_06040_),
    .Y(_06043_));
 sky130_fd_sc_hd__o22a_2 _16372_ (.A1(_05679_),
    .A2(_05681_),
    .B1(_06036_),
    .B2(_06038_),
    .X(_06044_));
 sky130_fd_sc_hd__o22ai_4 _16373_ (.A1(_05679_),
    .A2(_05681_),
    .B1(_06036_),
    .B2(_06038_),
    .Y(_06045_));
 sky130_fd_sc_hd__a21oi_2 _16374_ (.A1(_05630_),
    .A2(_05616_),
    .B1(_05628_),
    .Y(_06046_));
 sky130_fd_sc_hd__a21o_2 _16375_ (.A1(_05616_),
    .A2(_05630_),
    .B1(_05628_),
    .X(_06047_));
 sky130_fd_sc_hd__o21ai_2 _16376_ (.A1(_05695_),
    .A2(_05700_),
    .B1(_05698_),
    .Y(_06048_));
 sky130_fd_sc_hd__a22oi_1 _16377_ (.A1(net64),
    .A2(net15),
    .B1(net16),
    .B2(net63),
    .Y(_06049_));
 sky130_fd_sc_hd__a22o_1 _16378_ (.A1(net64),
    .A2(net15),
    .B1(net16),
    .B2(net63),
    .X(_06051_));
 sky130_fd_sc_hd__and4_1 _16379_ (.A(net63),
    .B(net64),
    .C(net15),
    .D(net16),
    .X(_06052_));
 sky130_fd_sc_hd__nand4_2 _16380_ (.A(net63),
    .B(net64),
    .C(net15),
    .D(net16),
    .Y(_06053_));
 sky130_fd_sc_hd__nand3_1 _16381_ (.A(_05696_),
    .B(_06051_),
    .C(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__a21o_1 _16382_ (.A1(_06051_),
    .A2(_06053_),
    .B1(_05696_),
    .X(_06055_));
 sky130_fd_sc_hd__a22o_1 _16383_ (.A1(net34),
    .A2(net14),
    .B1(_06051_),
    .B2(_06053_),
    .X(_06056_));
 sky130_fd_sc_hd__nand4_2 _16384_ (.A(_06051_),
    .B(_06053_),
    .C(net34),
    .D(net14),
    .Y(_06057_));
 sky130_fd_sc_hd__nand3_4 _16385_ (.A(_06056_),
    .B(_06057_),
    .C(_06048_),
    .Y(_06058_));
 sky130_fd_sc_hd__a21oi_1 _16386_ (.A1(_06056_),
    .A2(_06057_),
    .B1(_06048_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand3b_4 _16387_ (.A_N(_06048_),
    .B(_06054_),
    .C(_06055_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _16388_ (.A(net35),
    .B(net13),
    .Y(_06062_));
 sky130_fd_sc_hd__nand2_1 _16389_ (.A(net36),
    .B(net11),
    .Y(_06063_));
 sky130_fd_sc_hd__a22oi_4 _16390_ (.A1(net36),
    .A2(net11),
    .B1(net13),
    .B2(net35),
    .Y(_06064_));
 sky130_fd_sc_hd__nand2_1 _16391_ (.A(net36),
    .B(net13),
    .Y(_06065_));
 sky130_fd_sc_hd__and4_4 _16392_ (.A(net35),
    .B(net36),
    .C(net11),
    .D(net13),
    .X(_06066_));
 sky130_fd_sc_hd__a211oi_4 _16393_ (.A1(net37),
    .A2(net10),
    .B1(_06064_),
    .C1(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__a211o_1 _16394_ (.A1(net37),
    .A2(net10),
    .B1(_06064_),
    .C1(_06066_),
    .X(_06068_));
 sky130_fd_sc_hd__o211a_2 _16395_ (.A1(_06064_),
    .A2(_06066_),
    .B1(net37),
    .C1(net10),
    .X(_06069_));
 sky130_fd_sc_hd__o211ai_1 _16396_ (.A1(_06064_),
    .A2(_06066_),
    .B1(net37),
    .C1(net10),
    .Y(_06070_));
 sky130_fd_sc_hd__o2bb2a_1 _16397_ (.A1_N(net37),
    .A2_N(net10),
    .B1(_06064_),
    .B2(_06066_),
    .X(_06071_));
 sky130_fd_sc_hd__nor3_2 _16398_ (.A(_05715_),
    .B(_06064_),
    .C(_06066_),
    .Y(_06073_));
 sky130_fd_sc_hd__o211ai_4 _16399_ (.A1(_06071_),
    .A2(_06073_),
    .B1(_06058_),
    .C1(_06060_),
    .Y(_06074_));
 sky130_fd_sc_hd__o2bb2ai_2 _16400_ (.A1_N(_06058_),
    .A2_N(_06060_),
    .B1(_06067_),
    .B2(_06069_),
    .Y(_06075_));
 sky130_fd_sc_hd__o2bb2ai_2 _16401_ (.A1_N(_06058_),
    .A2_N(_06060_),
    .B1(_06071_),
    .B2(_06073_),
    .Y(_06076_));
 sky130_fd_sc_hd__o211ai_4 _16402_ (.A1(_06067_),
    .A2(_06069_),
    .B1(_06058_),
    .C1(_06060_),
    .Y(_06077_));
 sky130_fd_sc_hd__and3_1 _16403_ (.A(_06075_),
    .B(_06046_),
    .C(_06074_),
    .X(_06078_));
 sky130_fd_sc_hd__nand4_2 _16404_ (.A(_05629_),
    .B(_05631_),
    .C(_06074_),
    .D(_06075_),
    .Y(_06079_));
 sky130_fd_sc_hd__and3_1 _16405_ (.A(_06047_),
    .B(_06076_),
    .C(_06077_),
    .X(_06080_));
 sky130_fd_sc_hd__nand3_2 _16406_ (.A(_06047_),
    .B(_06076_),
    .C(_06077_),
    .Y(_06081_));
 sky130_fd_sc_hd__a2bb2o_2 _16407_ (.A1_N(_05707_),
    .A2_N(_05704_),
    .B1(_05725_),
    .B2(_05711_),
    .X(_06082_));
 sky130_fd_sc_hd__a31o_2 _16408_ (.A1(_05708_),
    .A2(_05719_),
    .A3(_05722_),
    .B1(_05709_),
    .X(_06084_));
 sky130_fd_sc_hd__a31oi_4 _16409_ (.A1(_06075_),
    .A2(_06046_),
    .A3(_06074_),
    .B1(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__a31o_1 _16410_ (.A1(_06046_),
    .A2(_06074_),
    .A3(_06075_),
    .B1(_06084_),
    .X(_06086_));
 sky130_fd_sc_hd__and3_1 _16411_ (.A(_06079_),
    .B(_06081_),
    .C(_06082_),
    .X(_06087_));
 sky130_fd_sc_hd__a21oi_1 _16412_ (.A1(_06079_),
    .A2(_06081_),
    .B1(_06082_),
    .Y(_06088_));
 sky130_fd_sc_hd__a21o_1 _16413_ (.A1(_06079_),
    .A2(_06081_),
    .B1(_06082_),
    .X(_06089_));
 sky130_fd_sc_hd__a21oi_2 _16414_ (.A1(_06079_),
    .A2(_06081_),
    .B1(_06084_),
    .Y(_06090_));
 sky130_fd_sc_hd__and3_2 _16415_ (.A(_06079_),
    .B(_06081_),
    .C(_06084_),
    .X(_06091_));
 sky130_fd_sc_hd__o21ai_2 _16416_ (.A1(_06080_),
    .A2(_06086_),
    .B1(_06089_),
    .Y(_06092_));
 sky130_fd_sc_hd__nand3_1 _16417_ (.A(_06043_),
    .B(_06045_),
    .C(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__o2bb2ai_1 _16418_ (.A1_N(_06043_),
    .A2_N(_06045_),
    .B1(_06090_),
    .B2(_06091_),
    .Y(_06095_));
 sky130_fd_sc_hd__o2bb2ai_2 _16419_ (.A1_N(_06043_),
    .A2_N(_06045_),
    .B1(_06087_),
    .B2(_06088_),
    .Y(_06096_));
 sky130_fd_sc_hd__o21ai_1 _16420_ (.A1(_06090_),
    .A2(_06091_),
    .B1(_06045_),
    .Y(_06097_));
 sky130_fd_sc_hd__o211a_1 _16421_ (.A1(_06090_),
    .A2(_06091_),
    .B1(_06043_),
    .C1(_06045_),
    .X(_06098_));
 sky130_fd_sc_hd__nand3_4 _16422_ (.A(_06095_),
    .B(_05972_),
    .C(_06093_),
    .Y(_06099_));
 sky130_fd_sc_hd__o21ai_2 _16423_ (.A1(_05690_),
    .A2(_05744_),
    .B1(_06096_),
    .Y(_06100_));
 sky130_fd_sc_hd__o221ai_4 _16424_ (.A1(_05690_),
    .A2(_05744_),
    .B1(_06042_),
    .B2(_06097_),
    .C1(_06096_),
    .Y(_06101_));
 sky130_fd_sc_hd__o21ai_1 _16425_ (.A1(_05712_),
    .A2(_05713_),
    .B1(_05717_),
    .Y(_06102_));
 sky130_fd_sc_hd__o21a_1 _16426_ (.A1(_05712_),
    .A2(_05713_),
    .B1(_05717_),
    .X(_06103_));
 sky130_fd_sc_hd__a22oi_4 _16427_ (.A1(net39),
    .A2(net8),
    .B1(net9),
    .B2(net38),
    .Y(_06104_));
 sky130_fd_sc_hd__a22o_1 _16428_ (.A1(net39),
    .A2(net8),
    .B1(net9),
    .B2(net38),
    .X(_06106_));
 sky130_fd_sc_hd__and4_4 _16429_ (.A(net38),
    .B(net39),
    .C(net8),
    .D(net9),
    .X(_06107_));
 sky130_fd_sc_hd__nand4_4 _16430_ (.A(net38),
    .B(net39),
    .C(net8),
    .D(net9),
    .Y(_06108_));
 sky130_fd_sc_hd__nand3_1 _16431_ (.A(_05793_),
    .B(_06106_),
    .C(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__o21bai_2 _16432_ (.A1(_06104_),
    .A2(_06107_),
    .B1_N(_05793_),
    .Y(_06110_));
 sky130_fd_sc_hd__o21ai_1 _16433_ (.A1(_06104_),
    .A2(_06107_),
    .B1(_05793_),
    .Y(_06111_));
 sky130_fd_sc_hd__nand4_1 _16434_ (.A(_06106_),
    .B(_06108_),
    .C(net7),
    .D(net40),
    .Y(_06112_));
 sky130_fd_sc_hd__a21oi_1 _16435_ (.A1(_06111_),
    .A2(_06112_),
    .B1(_06102_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand3_4 _16436_ (.A(_06103_),
    .B(_06109_),
    .C(_06110_),
    .Y(_06114_));
 sky130_fd_sc_hd__nand3_2 _16437_ (.A(_06111_),
    .B(_06112_),
    .C(_06102_),
    .Y(_06115_));
 sky130_fd_sc_hd__and3_1 _16438_ (.A(_05792_),
    .B(net41),
    .C(net5),
    .X(_06117_));
 sky130_fd_sc_hd__a31o_1 _16439_ (.A1(_05792_),
    .A2(net41),
    .A3(net5),
    .B1(_05794_),
    .X(_06118_));
 sky130_fd_sc_hd__o31a_1 _16440_ (.A1(_01956_),
    .A2(_02010_),
    .A3(_05791_),
    .B1(_05795_),
    .X(_06119_));
 sky130_fd_sc_hd__a21o_1 _16441_ (.A1(_06114_),
    .A2(_06115_),
    .B1(_06118_),
    .X(_06120_));
 sky130_fd_sc_hd__o211ai_2 _16442_ (.A1(_05794_),
    .A2(_06117_),
    .B1(_06115_),
    .C1(_06114_),
    .Y(_06121_));
 sky130_fd_sc_hd__o2111ai_1 _16443_ (.A1(_05790_),
    .A2(_05791_),
    .B1(_05795_),
    .C1(_06114_),
    .D1(_06115_),
    .Y(_06122_));
 sky130_fd_sc_hd__o2bb2ai_1 _16444_ (.A1_N(_06114_),
    .A2_N(_06115_),
    .B1(_06117_),
    .B2(_05794_),
    .Y(_06123_));
 sky130_fd_sc_hd__o21ai_2 _16445_ (.A1(_05785_),
    .A2(_05803_),
    .B1(_05802_),
    .Y(_06124_));
 sky130_fd_sc_hd__a21oi_1 _16446_ (.A1(_05804_),
    .A2(_05784_),
    .B1(_05801_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand3_2 _16447_ (.A(_06122_),
    .B(_06123_),
    .C(_06125_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand3_4 _16448_ (.A(_06120_),
    .B(_06124_),
    .C(_06121_),
    .Y(_06128_));
 sky130_fd_sc_hd__a31o_1 _16449_ (.A1(_05768_),
    .A2(net45),
    .A3(net2),
    .B1(_05766_),
    .X(_06129_));
 sky130_fd_sc_hd__a31oi_1 _16450_ (.A1(_05768_),
    .A2(net45),
    .A3(net2),
    .B1(_05766_),
    .Y(_06130_));
 sky130_fd_sc_hd__a22oi_4 _16451_ (.A1(net6),
    .A2(net41),
    .B1(net42),
    .B2(net5),
    .Y(_06131_));
 sky130_fd_sc_hd__a22o_2 _16452_ (.A1(net6),
    .A2(net41),
    .B1(net42),
    .B2(net5),
    .X(_06132_));
 sky130_fd_sc_hd__and4_1 _16453_ (.A(net5),
    .B(net6),
    .C(net41),
    .D(net42),
    .X(_06133_));
 sky130_fd_sc_hd__nand4_4 _16454_ (.A(net5),
    .B(net6),
    .C(net41),
    .D(net42),
    .Y(_06134_));
 sky130_fd_sc_hd__nand3_1 _16455_ (.A(_05764_),
    .B(_06132_),
    .C(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__a21o_1 _16456_ (.A1(_06132_),
    .A2(_06134_),
    .B1(_05764_),
    .X(_06136_));
 sky130_fd_sc_hd__a22o_1 _16457_ (.A1(net4),
    .A2(net43),
    .B1(_06132_),
    .B2(_06134_),
    .X(_06137_));
 sky130_fd_sc_hd__nand4_2 _16458_ (.A(_06132_),
    .B(_06134_),
    .C(net4),
    .D(net43),
    .Y(_06139_));
 sky130_fd_sc_hd__nand3_2 _16459_ (.A(_06130_),
    .B(_06135_),
    .C(_06136_),
    .Y(_06140_));
 sky130_fd_sc_hd__nand3_4 _16460_ (.A(_06129_),
    .B(_06137_),
    .C(_06139_),
    .Y(_06141_));
 sky130_fd_sc_hd__nand2_2 _16461_ (.A(net3),
    .B(net46),
    .Y(_06142_));
 sky130_fd_sc_hd__and4_2 _16462_ (.A(net2),
    .B(net3),
    .C(net45),
    .D(net46),
    .X(_06143_));
 sky130_fd_sc_hd__nand4_1 _16463_ (.A(net2),
    .B(net3),
    .C(net45),
    .D(net46),
    .Y(_06144_));
 sky130_fd_sc_hd__a22oi_2 _16464_ (.A1(net3),
    .A2(net45),
    .B1(net46),
    .B2(net2),
    .Y(_06145_));
 sky130_fd_sc_hd__a22o_1 _16465_ (.A1(net3),
    .A2(net45),
    .B1(net46),
    .B2(net2),
    .X(_06146_));
 sky130_fd_sc_hd__o311a_1 _16466_ (.A1(_01901_),
    .A2(_02054_),
    .A3(_06142_),
    .B1(_06146_),
    .C1(_05756_),
    .X(_06147_));
 sky130_fd_sc_hd__o211a_1 _16467_ (.A1(_06143_),
    .A2(_06145_),
    .B1(net32),
    .C1(net47),
    .X(_06148_));
 sky130_fd_sc_hd__a22oi_1 _16468_ (.A1(net32),
    .A2(net47),
    .B1(_06144_),
    .B2(_06146_),
    .Y(_06150_));
 sky130_fd_sc_hd__and3_1 _16469_ (.A(_06144_),
    .B(net47),
    .C(net32),
    .X(_06151_));
 sky130_fd_sc_hd__a21oi_2 _16470_ (.A1(_06151_),
    .A2(_06146_),
    .B1(_06150_),
    .Y(_06152_));
 sky130_fd_sc_hd__o21ai_2 _16471_ (.A1(_06147_),
    .A2(_06148_),
    .B1(_06140_),
    .Y(_06153_));
 sky130_fd_sc_hd__and3_1 _16472_ (.A(_06140_),
    .B(_06141_),
    .C(_06152_),
    .X(_06154_));
 sky130_fd_sc_hd__a21oi_2 _16473_ (.A1(_06140_),
    .A2(_06141_),
    .B1(_06152_),
    .Y(_06155_));
 sky130_fd_sc_hd__nand3b_1 _16474_ (.A_N(_06152_),
    .B(_06141_),
    .C(_06140_),
    .Y(_06156_));
 sky130_fd_sc_hd__o2bb2ai_1 _16475_ (.A1_N(_06140_),
    .A2_N(_06141_),
    .B1(_06147_),
    .B2(_06148_),
    .Y(_06157_));
 sky130_fd_sc_hd__nand2_1 _16476_ (.A(_06156_),
    .B(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__o2bb2ai_4 _16477_ (.A1_N(_06126_),
    .A2_N(_06128_),
    .B1(_06154_),
    .B2(_06155_),
    .Y(_06159_));
 sky130_fd_sc_hd__nand3_4 _16478_ (.A(_06158_),
    .B(_06128_),
    .C(_06126_),
    .Y(_06161_));
 sky130_fd_sc_hd__a32oi_4 _16479_ (.A1(_05693_),
    .A2(_05726_),
    .A3(_05727_),
    .B1(_05733_),
    .B2(_05734_),
    .Y(_06162_));
 sky130_fd_sc_hd__a21oi_4 _16480_ (.A1(_06159_),
    .A2(_06161_),
    .B1(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__a21o_1 _16481_ (.A1(_06159_),
    .A2(_06161_),
    .B1(_06162_),
    .X(_06164_));
 sky130_fd_sc_hd__o211a_1 _16482_ (.A1(_05731_),
    .A2(_05740_),
    .B1(_06159_),
    .C1(_06161_),
    .X(_06165_));
 sky130_fd_sc_hd__o211ai_4 _16483_ (.A1(_05731_),
    .A2(_05740_),
    .B1(_06159_),
    .C1(_06161_),
    .Y(_06166_));
 sky130_fd_sc_hd__nor2_2 _16484_ (.A(_05810_),
    .B(_05813_),
    .Y(_06167_));
 sky130_fd_sc_hd__o211a_1 _16485_ (.A1(_05810_),
    .A2(_05813_),
    .B1(_06164_),
    .C1(_06166_),
    .X(_06168_));
 sky130_fd_sc_hd__o21a_1 _16486_ (.A1(_06163_),
    .A2(_06165_),
    .B1(_06167_),
    .X(_06169_));
 sky130_fd_sc_hd__and3_1 _16487_ (.A(_06164_),
    .B(_06166_),
    .C(_06167_),
    .X(_06170_));
 sky130_fd_sc_hd__nand3_1 _16488_ (.A(_06164_),
    .B(_06166_),
    .C(_06167_),
    .Y(_06172_));
 sky130_fd_sc_hd__o22a_1 _16489_ (.A1(_05810_),
    .A2(_05813_),
    .B1(_06163_),
    .B2(_06165_),
    .X(_06173_));
 sky130_fd_sc_hd__o22ai_1 _16490_ (.A1(_05810_),
    .A2(_05813_),
    .B1(_06163_),
    .B2(_06165_),
    .Y(_06174_));
 sky130_fd_sc_hd__nand2_2 _16491_ (.A(_06172_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__o211ai_4 _16492_ (.A1(_06168_),
    .A2(_06169_),
    .B1(_06099_),
    .C1(_06101_),
    .Y(_06176_));
 sky130_fd_sc_hd__o2bb2ai_2 _16493_ (.A1_N(_06099_),
    .A2_N(_06101_),
    .B1(_06170_),
    .B2(_06173_),
    .Y(_06177_));
 sky130_fd_sc_hd__a21oi_1 _16494_ (.A1(_06099_),
    .A2(_06101_),
    .B1(_06175_),
    .Y(_06178_));
 sky130_fd_sc_hd__o2bb2ai_2 _16495_ (.A1_N(_06099_),
    .A2_N(_06101_),
    .B1(_06168_),
    .B2(_06169_),
    .Y(_06179_));
 sky130_fd_sc_hd__o211ai_4 _16496_ (.A1(_06170_),
    .A2(_06173_),
    .B1(_06099_),
    .C1(_06101_),
    .Y(_06180_));
 sky130_fd_sc_hd__a2bb2oi_2 _16497_ (.A1_N(_05745_),
    .A2_N(_05749_),
    .B1(_05834_),
    .B2(_05752_),
    .Y(_06181_));
 sky130_fd_sc_hd__o22ai_4 _16498_ (.A1(_05745_),
    .A2(_05749_),
    .B1(_05835_),
    .B2(_05751_),
    .Y(_06183_));
 sky130_fd_sc_hd__a21oi_1 _16499_ (.A1(_06179_),
    .A2(_06180_),
    .B1(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand3_2 _16500_ (.A(_06181_),
    .B(_06177_),
    .C(_06176_),
    .Y(_06185_));
 sky130_fd_sc_hd__nor2_1 _16501_ (.A(_06178_),
    .B(_06181_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand3_4 _16502_ (.A(_06179_),
    .B(_06180_),
    .C(_06183_),
    .Y(_06187_));
 sky130_fd_sc_hd__a32oi_4 _16503_ (.A1(_06181_),
    .A2(_06177_),
    .A3(_06176_),
    .B1(_05967_),
    .B2(_05969_),
    .Y(_06188_));
 sky130_fd_sc_hd__a32o_1 _16504_ (.A1(_06181_),
    .A2(_06177_),
    .A3(_06176_),
    .B1(_05967_),
    .B2(_05969_),
    .X(_06189_));
 sky130_fd_sc_hd__o211a_1 _16505_ (.A1(_05966_),
    .A2(_05968_),
    .B1(_06185_),
    .C1(_06187_),
    .X(_06190_));
 sky130_fd_sc_hd__nand2_1 _16506_ (.A(_06188_),
    .B(_06187_),
    .Y(_06191_));
 sky130_fd_sc_hd__a2bb2oi_4 _16507_ (.A1_N(_05963_),
    .A2_N(_05964_),
    .B1(_06185_),
    .B2(_06187_),
    .Y(_06192_));
 sky130_fd_sc_hd__a21o_1 _16508_ (.A1(_06185_),
    .A2(_06187_),
    .B1(_05970_),
    .X(_06194_));
 sky130_fd_sc_hd__a21oi_1 _16509_ (.A1(_06187_),
    .A2(_06188_),
    .B1(_06192_),
    .Y(_06195_));
 sky130_fd_sc_hd__a221oi_4 _16510_ (.A1(_06188_),
    .A2(_06187_),
    .B1(_05848_),
    .B2(_05845_),
    .C1(_06192_),
    .Y(_06196_));
 sky130_fd_sc_hd__nand3_2 _16511_ (.A(_05879_),
    .B(_06191_),
    .C(_06194_),
    .Y(_06197_));
 sky130_fd_sc_hd__a2bb2oi_2 _16512_ (.A1_N(_05841_),
    .A2_N(_05878_),
    .B1(_06191_),
    .B2(_06194_),
    .Y(_06198_));
 sky130_fd_sc_hd__o22ai_4 _16513_ (.A1(_05841_),
    .A2(_05878_),
    .B1(_06190_),
    .B2(_06192_),
    .Y(_06199_));
 sky130_fd_sc_hd__o22ai_2 _16514_ (.A1(_05596_),
    .A2(_05603_),
    .B1(_05879_),
    .B2(_06195_),
    .Y(_06200_));
 sky130_fd_sc_hd__o22ai_2 _16515_ (.A1(_05594_),
    .A2(_05875_),
    .B1(_06196_),
    .B2(_06198_),
    .Y(_06201_));
 sky130_fd_sc_hd__o22ai_2 _16516_ (.A1(_05596_),
    .A2(_05603_),
    .B1(_06196_),
    .B2(_06198_),
    .Y(_06202_));
 sky130_fd_sc_hd__o2111ai_4 _16517_ (.A1(_05599_),
    .A2(_05594_),
    .B1(_05597_),
    .C1(_06197_),
    .D1(_06199_),
    .Y(_06203_));
 sky130_fd_sc_hd__o221a_1 _16518_ (.A1(_05851_),
    .A2(_05860_),
    .B1(_06196_),
    .B2(_06200_),
    .C1(_06201_),
    .X(_06205_));
 sky130_fd_sc_hd__o221ai_4 _16519_ (.A1(_05851_),
    .A2(_05860_),
    .B1(_06196_),
    .B2(_06200_),
    .C1(_06201_),
    .Y(_06206_));
 sky130_fd_sc_hd__nand3_2 _16520_ (.A(_05873_),
    .B(_06202_),
    .C(_06203_),
    .Y(_06207_));
 sky130_fd_sc_hd__a31oi_2 _16521_ (.A1(_05873_),
    .A2(_06202_),
    .A3(_06203_),
    .B1(_05538_),
    .Y(_06208_));
 sky130_fd_sc_hd__and3_1 _16522_ (.A(_06206_),
    .B(_06207_),
    .C(_05537_),
    .X(_06209_));
 sky130_fd_sc_hd__nand3_1 _16523_ (.A(_06207_),
    .B(_05537_),
    .C(_06206_),
    .Y(_06210_));
 sky130_fd_sc_hd__o2bb2ai_2 _16524_ (.A1_N(_06206_),
    .A2_N(_06207_),
    .B1(_05221_),
    .B2(_05533_),
    .Y(_06211_));
 sky130_fd_sc_hd__o2bb2ai_1 _16525_ (.A1_N(_06210_),
    .A2_N(_06211_),
    .B1(_05517_),
    .B2(_05862_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_1 _16526_ (.A(_06211_),
    .B(_05866_),
    .Y(_06213_));
 sky130_fd_sc_hd__nand3_1 _16527_ (.A(_06211_),
    .B(_05866_),
    .C(_06210_),
    .Y(_06214_));
 sky130_fd_sc_hd__o21a_1 _16528_ (.A1(_06209_),
    .A2(_06213_),
    .B1(_06212_),
    .X(_06216_));
 sky130_fd_sc_hd__a22o_1 _16529_ (.A1(_05865_),
    .A2(_05868_),
    .B1(_05872_),
    .B2(_05870_),
    .X(_06217_));
 sky130_fd_sc_hd__xor2_1 _16530_ (.A(_06216_),
    .B(_06217_),
    .X(net89));
 sky130_fd_sc_hd__a21oi_1 _16531_ (.A1(_06207_),
    .A2(_05537_),
    .B1(_06205_),
    .Y(_06218_));
 sky130_fd_sc_hd__o21ai_2 _16532_ (.A1(_05876_),
    .A2(_06196_),
    .B1(_06199_),
    .Y(_06219_));
 sky130_fd_sc_hd__a21oi_1 _16533_ (.A1(_05877_),
    .A2(_06197_),
    .B1(_06198_),
    .Y(_06220_));
 sky130_fd_sc_hd__o2bb2ai_2 _16534_ (.A1_N(_06180_),
    .A2_N(_06186_),
    .B1(_06184_),
    .B2(_05971_),
    .Y(_06221_));
 sky130_fd_sc_hd__a31o_1 _16535_ (.A1(_05967_),
    .A2(_05969_),
    .A3(_06187_),
    .B1(_06184_),
    .X(_06222_));
 sky130_fd_sc_hd__o21ai_2 _16536_ (.A1(_06167_),
    .A2(_06163_),
    .B1(_06166_),
    .Y(_06223_));
 sky130_fd_sc_hd__a21o_1 _16537_ (.A1(_05937_),
    .A2(_05938_),
    .B1(_05934_),
    .X(_06224_));
 sky130_fd_sc_hd__a21oi_2 _16538_ (.A1(_05937_),
    .A2(_05938_),
    .B1(_05934_),
    .Y(_06226_));
 sky130_fd_sc_hd__a21oi_2 _16539_ (.A1(_05923_),
    .A2(_05927_),
    .B1(_05924_),
    .Y(_06227_));
 sky130_fd_sc_hd__a21o_1 _16540_ (.A1(_05923_),
    .A2(_05927_),
    .B1(_05924_),
    .X(_06228_));
 sky130_fd_sc_hd__a32o_2 _16541_ (.A1(_06129_),
    .A2(_06137_),
    .A3(_06139_),
    .B1(_06140_),
    .B2(_06152_),
    .X(_06229_));
 sky130_fd_sc_hd__o31a_1 _16542_ (.A1(_01879_),
    .A2(_02120_),
    .A3(_05755_),
    .B1(_05552_),
    .X(_06230_));
 sky130_fd_sc_hd__o21a_1 _16543_ (.A1(_05552_),
    .A2(_05914_),
    .B1(_05917_),
    .X(_06231_));
 sky130_fd_sc_hd__nor2_2 _16544_ (.A(_05756_),
    .B(_06145_),
    .Y(_06232_));
 sky130_fd_sc_hd__a31o_1 _16545_ (.A1(_06146_),
    .A2(net47),
    .A3(net32),
    .B1(_06143_),
    .X(_06233_));
 sky130_fd_sc_hd__o21a_1 _16546_ (.A1(_05756_),
    .A2(_06145_),
    .B1(_06144_),
    .X(_06234_));
 sky130_fd_sc_hd__nand2_2 _16547_ (.A(net29),
    .B(net51),
    .Y(_06235_));
 sky130_fd_sc_hd__a22oi_4 _16548_ (.A1(net31),
    .A2(net49),
    .B1(net50),
    .B2(net30),
    .Y(_06237_));
 sky130_fd_sc_hd__a22o_2 _16549_ (.A1(net31),
    .A2(net49),
    .B1(net50),
    .B2(net30),
    .X(_06238_));
 sky130_fd_sc_hd__and4_4 _16550_ (.A(net30),
    .B(net31),
    .C(net49),
    .D(net50),
    .X(_06239_));
 sky130_fd_sc_hd__nand4_4 _16551_ (.A(net30),
    .B(net31),
    .C(net49),
    .D(net50),
    .Y(_06240_));
 sky130_fd_sc_hd__o211ai_4 _16552_ (.A1(_01857_),
    .A2(_02152_),
    .B1(_06238_),
    .C1(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__o21bai_4 _16553_ (.A1(_06237_),
    .A2(_06239_),
    .B1_N(_06235_),
    .Y(_06242_));
 sky130_fd_sc_hd__nand4_2 _16554_ (.A(_06238_),
    .B(_06240_),
    .C(net29),
    .D(net51),
    .Y(_06243_));
 sky130_fd_sc_hd__o21ai_2 _16555_ (.A1(_06237_),
    .A2(_06239_),
    .B1(_06235_),
    .Y(_06244_));
 sky130_fd_sc_hd__a2bb2oi_4 _16556_ (.A1_N(_06143_),
    .A2_N(_06232_),
    .B1(_06241_),
    .B2(_06242_),
    .Y(_06245_));
 sky130_fd_sc_hd__o211ai_4 _16557_ (.A1(_06143_),
    .A2(_06232_),
    .B1(_06243_),
    .C1(_06244_),
    .Y(_06246_));
 sky130_fd_sc_hd__a21oi_1 _16558_ (.A1(_06243_),
    .A2(_06244_),
    .B1(_06233_),
    .Y(_06248_));
 sky130_fd_sc_hd__nand3_1 _16559_ (.A(_06234_),
    .B(_06241_),
    .C(_06242_),
    .Y(_06249_));
 sky130_fd_sc_hd__a31oi_4 _16560_ (.A1(_06234_),
    .A2(_06241_),
    .A3(_06242_),
    .B1(_06231_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand2_1 _16561_ (.A(_06250_),
    .B(_06246_),
    .Y(_06251_));
 sky130_fd_sc_hd__a2bb2oi_2 _16562_ (.A1_N(_05914_),
    .A2_N(_06230_),
    .B1(_06246_),
    .B2(_06249_),
    .Y(_06252_));
 sky130_fd_sc_hd__o22ai_2 _16563_ (.A1(_05914_),
    .A2(_06230_),
    .B1(_06245_),
    .B2(_06248_),
    .Y(_06253_));
 sky130_fd_sc_hd__a21oi_2 _16564_ (.A1(_06246_),
    .A2(_06250_),
    .B1(_06252_),
    .Y(_06254_));
 sky130_fd_sc_hd__a221oi_4 _16565_ (.A1(_06250_),
    .A2(_06246_),
    .B1(_06153_),
    .B2(_06141_),
    .C1(_06252_),
    .Y(_06255_));
 sky130_fd_sc_hd__a221o_2 _16566_ (.A1(_06250_),
    .A2(_06246_),
    .B1(_06153_),
    .B2(_06141_),
    .C1(_06252_),
    .X(_06256_));
 sky130_fd_sc_hd__a21oi_4 _16567_ (.A1(_06251_),
    .A2(_06253_),
    .B1(_06229_),
    .Y(_06257_));
 sky130_fd_sc_hd__o21ai_1 _16568_ (.A1(_06255_),
    .A2(_06257_),
    .B1(_06227_),
    .Y(_06259_));
 sky130_fd_sc_hd__o22a_1 _16569_ (.A1(_05924_),
    .A2(_05931_),
    .B1(_06229_),
    .B2(_06254_),
    .X(_06260_));
 sky130_fd_sc_hd__o22ai_4 _16570_ (.A1(_05924_),
    .A2(_05931_),
    .B1(_06229_),
    .B2(_06254_),
    .Y(_06261_));
 sky130_fd_sc_hd__nand3b_1 _16571_ (.A_N(_06257_),
    .B(_06227_),
    .C(_06256_),
    .Y(_06262_));
 sky130_fd_sc_hd__o21ai_1 _16572_ (.A1(_06255_),
    .A2(_06257_),
    .B1(_06228_),
    .Y(_06263_));
 sky130_fd_sc_hd__o211ai_4 _16573_ (.A1(_06261_),
    .A2(_06255_),
    .B1(_06226_),
    .C1(_06259_),
    .Y(_06264_));
 sky130_fd_sc_hd__nand3_4 _16574_ (.A(_06262_),
    .B(_06263_),
    .C(_06224_),
    .Y(_06265_));
 sky130_fd_sc_hd__o31a_2 _16575_ (.A1(_01802_),
    .A2(_02229_),
    .A3(_05519_),
    .B1(_05888_),
    .X(_06266_));
 sky130_fd_sc_hd__o21ai_2 _16576_ (.A1(_05520_),
    .A2(_05891_),
    .B1(_05893_),
    .Y(_06267_));
 sky130_fd_sc_hd__nor2_1 _16577_ (.A(_01791_),
    .B(_02207_),
    .Y(_06268_));
 sky130_fd_sc_hd__a22oi_4 _16578_ (.A1(net28),
    .A2(net52),
    .B1(net53),
    .B2(net27),
    .Y(_06270_));
 sky130_fd_sc_hd__a22o_1 _16579_ (.A1(net28),
    .A2(net52),
    .B1(net53),
    .B2(net27),
    .X(_06271_));
 sky130_fd_sc_hd__nand2_1 _16580_ (.A(net28),
    .B(net53),
    .Y(_06272_));
 sky130_fd_sc_hd__and4_1 _16581_ (.A(net28),
    .B(net27),
    .C(net52),
    .D(net53),
    .X(_06273_));
 sky130_fd_sc_hd__nand4_2 _16582_ (.A(net28),
    .B(net27),
    .C(net52),
    .D(net53),
    .Y(_06274_));
 sky130_fd_sc_hd__o211ai_1 _16583_ (.A1(_01791_),
    .A2(_02207_),
    .B1(_06271_),
    .C1(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__o21ai_1 _16584_ (.A1(_06270_),
    .A2(_06273_),
    .B1(_06268_),
    .Y(_06276_));
 sky130_fd_sc_hd__and4_2 _16585_ (.A(_06271_),
    .B(_06274_),
    .C(net26),
    .D(net54),
    .X(_06277_));
 sky130_fd_sc_hd__nand4_1 _16586_ (.A(_06271_),
    .B(_06274_),
    .C(net26),
    .D(net54),
    .Y(_06278_));
 sky130_fd_sc_hd__a22o_1 _16587_ (.A1(net26),
    .A2(net54),
    .B1(_06271_),
    .B2(_06274_),
    .X(_06279_));
 sky130_fd_sc_hd__nand2_2 _16588_ (.A(_06279_),
    .B(_06267_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand3_1 _16589_ (.A(_06279_),
    .B(_06267_),
    .C(_06278_),
    .Y(_06282_));
 sky130_fd_sc_hd__nand3b_2 _16590_ (.A_N(_06267_),
    .B(_06275_),
    .C(_06276_),
    .Y(_06283_));
 sky130_fd_sc_hd__and4_2 _16591_ (.A(_01824_),
    .B(net56),
    .C(net57),
    .D(net23),
    .X(_06284_));
 sky130_fd_sc_hd__o22a_1 _16592_ (.A1(net12),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01802_),
    .X(_06285_));
 sky130_fd_sc_hd__nor2_2 _16593_ (.A(_06284_),
    .B(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__a21o_2 _16594_ (.A1(_06282_),
    .A2(_06283_),
    .B1(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__o211ai_4 _16595_ (.A1(_06277_),
    .A2(_06281_),
    .B1(_06283_),
    .C1(_06286_),
    .Y(_06288_));
 sky130_fd_sc_hd__a21oi_2 _16596_ (.A1(_05889_),
    .A2(_05901_),
    .B1(_05898_),
    .Y(_06289_));
 sky130_fd_sc_hd__a21oi_4 _16597_ (.A1(_06287_),
    .A2(_06288_),
    .B1(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__and3_1 _16598_ (.A(_06287_),
    .B(_06288_),
    .C(_06289_),
    .X(_06292_));
 sky130_fd_sc_hd__nand3_2 _16599_ (.A(_06287_),
    .B(_06288_),
    .C(_06289_),
    .Y(_06293_));
 sky130_fd_sc_hd__o2bb2a_1 _16600_ (.A1_N(_05886_),
    .A2_N(_05888_),
    .B1(_06290_),
    .B2(_06292_),
    .X(_06294_));
 sky130_fd_sc_hd__o21bai_1 _16601_ (.A1(_06290_),
    .A2(_06292_),
    .B1_N(_06266_),
    .Y(_06295_));
 sky130_fd_sc_hd__and3b_1 _16602_ (.A_N(_06290_),
    .B(_06293_),
    .C(_06266_),
    .X(_06296_));
 sky130_fd_sc_hd__nand3b_1 _16603_ (.A_N(_06290_),
    .B(_06293_),
    .C(_06266_),
    .Y(_06297_));
 sky130_fd_sc_hd__o221a_1 _16604_ (.A1(_05519_),
    .A2(_05884_),
    .B1(_06290_),
    .B2(_06292_),
    .C1(_05888_),
    .X(_06298_));
 sky130_fd_sc_hd__a311oi_1 _16605_ (.A1(_06287_),
    .A2(_06288_),
    .A3(_06289_),
    .B1(_06290_),
    .C1(_06266_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2_1 _16606_ (.A(_06295_),
    .B(_06297_),
    .Y(_06300_));
 sky130_fd_sc_hd__nand4_2 _16607_ (.A(_06264_),
    .B(_06265_),
    .C(_06295_),
    .D(_06297_),
    .Y(_06301_));
 sky130_fd_sc_hd__o2bb2ai_1 _16608_ (.A1_N(_06264_),
    .A2_N(_06265_),
    .B1(_06294_),
    .B2(_06296_),
    .Y(_06303_));
 sky130_fd_sc_hd__o2bb2ai_2 _16609_ (.A1_N(_06264_),
    .A2_N(_06265_),
    .B1(_06298_),
    .B2(_06299_),
    .Y(_06304_));
 sky130_fd_sc_hd__nand3_2 _16610_ (.A(_06264_),
    .B(_06265_),
    .C(_06300_),
    .Y(_06305_));
 sky130_fd_sc_hd__o2111ai_4 _16611_ (.A1(_06167_),
    .A2(_06163_),
    .B1(_06166_),
    .C1(_06301_),
    .D1(_06303_),
    .Y(_06306_));
 sky130_fd_sc_hd__nand3_2 _16612_ (.A(_06304_),
    .B(_06305_),
    .C(_06223_),
    .Y(_06307_));
 sky130_fd_sc_hd__a31o_1 _16613_ (.A1(_05906_),
    .A2(_05910_),
    .A3(_05949_),
    .B1(_05947_),
    .X(_06308_));
 sky130_fd_sc_hd__a21o_2 _16614_ (.A1(_06306_),
    .A2(_06307_),
    .B1(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__o21a_1 _16615_ (.A1(_05947_),
    .A2(_05952_),
    .B1(_06306_),
    .X(_06310_));
 sky130_fd_sc_hd__o211ai_4 _16616_ (.A1(_05947_),
    .A2(_05952_),
    .B1(_06306_),
    .C1(_06307_),
    .Y(_06311_));
 sky130_fd_sc_hd__nand2_2 _16617_ (.A(_06309_),
    .B(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__a311oi_4 _16618_ (.A1(_06040_),
    .A2(_05682_),
    .A3(_06037_),
    .B1(_06090_),
    .C1(_06091_),
    .Y(_06314_));
 sky130_fd_sc_hd__o22ai_4 _16619_ (.A1(_06036_),
    .A2(_06041_),
    .B1(_06092_),
    .B2(_06044_),
    .Y(_06315_));
 sky130_fd_sc_hd__a21oi_4 _16620_ (.A1(_05993_),
    .A2(_06033_),
    .B1(_06031_),
    .Y(_06316_));
 sky130_fd_sc_hd__o21a_1 _16621_ (.A1(_06002_),
    .A2(_06005_),
    .B1(_06025_),
    .X(_06317_));
 sky130_fd_sc_hd__o21ai_2 _16622_ (.A1(_06007_),
    .A2(_06022_),
    .B1(_06025_),
    .Y(_06318_));
 sky130_fd_sc_hd__o31a_1 _16623_ (.A1(_06002_),
    .A2(_06005_),
    .A3(_06022_),
    .B1(_06025_),
    .X(_06319_));
 sky130_fd_sc_hd__nand2_1 _16624_ (.A(net60),
    .B(net20),
    .Y(_06320_));
 sky130_fd_sc_hd__a22oi_4 _16625_ (.A1(net59),
    .A2(net21),
    .B1(net22),
    .B2(net58),
    .Y(_06321_));
 sky130_fd_sc_hd__a22o_1 _16626_ (.A1(net59),
    .A2(net21),
    .B1(net22),
    .B2(net58),
    .X(_06322_));
 sky130_fd_sc_hd__and4_1 _16627_ (.A(net58),
    .B(net59),
    .C(net21),
    .D(net22),
    .X(_06323_));
 sky130_fd_sc_hd__nand4_1 _16628_ (.A(net58),
    .B(net59),
    .C(net21),
    .D(net22),
    .Y(_06325_));
 sky130_fd_sc_hd__o211a_1 _16629_ (.A1(_06321_),
    .A2(_06323_),
    .B1(net60),
    .C1(net20),
    .X(_06326_));
 sky130_fd_sc_hd__and3_1 _16630_ (.A(_06320_),
    .B(_06322_),
    .C(_06325_),
    .X(_06327_));
 sky130_fd_sc_hd__o22a_2 _16631_ (.A1(_01835_),
    .A2(_02163_),
    .B1(_06321_),
    .B2(_06323_),
    .X(_06328_));
 sky130_fd_sc_hd__o22ai_4 _16632_ (.A1(_01835_),
    .A2(_02163_),
    .B1(_06321_),
    .B2(_06323_),
    .Y(_06329_));
 sky130_fd_sc_hd__a41o_1 _16633_ (.A1(net58),
    .A2(net59),
    .A3(net21),
    .A4(net22),
    .B1(_06320_),
    .X(_06330_));
 sky130_fd_sc_hd__and4_2 _16634_ (.A(_06322_),
    .B(_06325_),
    .C(net60),
    .D(net20),
    .X(_06331_));
 sky130_fd_sc_hd__o21ai_1 _16635_ (.A1(_06321_),
    .A2(_06330_),
    .B1(_06329_),
    .Y(_06332_));
 sky130_fd_sc_hd__o21a_1 _16636_ (.A1(_06321_),
    .A2(_06330_),
    .B1(_06329_),
    .X(_06333_));
 sky130_fd_sc_hd__a31o_1 _16637_ (.A1(_06013_),
    .A2(net24),
    .A3(net44),
    .B1(_06014_),
    .X(_06334_));
 sky130_fd_sc_hd__o31a_2 _16638_ (.A1(_01759_),
    .A2(_02218_),
    .A3(_06012_),
    .B1(_06015_),
    .X(_06336_));
 sky130_fd_sc_hd__nand2_1 _16639_ (.A(net55),
    .B(net24),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _16640_ (.A(net44),
    .B(net25),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _16641_ (.A(net33),
    .B(net44),
    .Y(_06339_));
 sky130_fd_sc_hd__and3_1 _16642_ (.A(net33),
    .B(net44),
    .C(net25),
    .X(_06340_));
 sky130_fd_sc_hd__nand3_4 _16643_ (.A(net33),
    .B(net44),
    .C(net25),
    .Y(_06341_));
 sky130_fd_sc_hd__o21a_2 _16644_ (.A1(net33),
    .A2(net44),
    .B1(net25),
    .X(_06342_));
 sky130_fd_sc_hd__o2bb2ai_1 _16645_ (.A1_N(_06011_),
    .A2_N(_06338_),
    .B1(_06339_),
    .B2(_02251_),
    .Y(_06343_));
 sky130_fd_sc_hd__o221ai_4 _16646_ (.A1(_01780_),
    .A2(_02218_),
    .B1(_06011_),
    .B2(_01759_),
    .C1(_06342_),
    .Y(_06344_));
 sky130_fd_sc_hd__a21o_1 _16647_ (.A1(_06341_),
    .A2(_06342_),
    .B1(_06337_),
    .X(_06345_));
 sky130_fd_sc_hd__o2bb2ai_2 _16648_ (.A1_N(_06341_),
    .A2_N(_06342_),
    .B1(_01780_),
    .B2(_02218_),
    .Y(_06347_));
 sky130_fd_sc_hd__o2111ai_4 _16649_ (.A1(net33),
    .A2(net44),
    .B1(net55),
    .C1(net24),
    .D1(net25),
    .Y(_06348_));
 sky130_fd_sc_hd__o2111ai_1 _16650_ (.A1(_01759_),
    .A2(_06011_),
    .B1(_06342_),
    .C1(net55),
    .D1(net24),
    .Y(_06349_));
 sky130_fd_sc_hd__o221a_2 _16651_ (.A1(_06340_),
    .A2(_06348_),
    .B1(_06014_),
    .B2(_06018_),
    .C1(_06347_),
    .X(_06350_));
 sky130_fd_sc_hd__o221ai_4 _16652_ (.A1(_06340_),
    .A2(_06348_),
    .B1(_06014_),
    .B2(_06018_),
    .C1(_06347_),
    .Y(_06351_));
 sky130_fd_sc_hd__a21oi_2 _16653_ (.A1(_06347_),
    .A2(_06349_),
    .B1(_06334_),
    .Y(_06352_));
 sky130_fd_sc_hd__nand3_4 _16654_ (.A(_06336_),
    .B(_06344_),
    .C(_06345_),
    .Y(_06353_));
 sky130_fd_sc_hd__o211ai_4 _16655_ (.A1(_06328_),
    .A2(_06331_),
    .B1(_06351_),
    .C1(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__o22ai_4 _16656_ (.A1(_06326_),
    .A2(_06327_),
    .B1(_06350_),
    .B2(_06352_),
    .Y(_06355_));
 sky130_fd_sc_hd__and3_1 _16657_ (.A(_06333_),
    .B(_06351_),
    .C(_06353_),
    .X(_06356_));
 sky130_fd_sc_hd__o2111ai_4 _16658_ (.A1(_06330_),
    .A2(_06321_),
    .B1(_06329_),
    .C1(_06351_),
    .D1(_06353_),
    .Y(_06358_));
 sky130_fd_sc_hd__o22ai_4 _16659_ (.A1(_06328_),
    .A2(_06331_),
    .B1(_06350_),
    .B2(_06352_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand2_2 _16660_ (.A(_06359_),
    .B(_06318_),
    .Y(_06360_));
 sky130_fd_sc_hd__and3_1 _16661_ (.A(_06359_),
    .B(_06318_),
    .C(_06358_),
    .X(_06361_));
 sky130_fd_sc_hd__nand3_4 _16662_ (.A(_06359_),
    .B(_06318_),
    .C(_06358_),
    .Y(_06362_));
 sky130_fd_sc_hd__nand2_2 _16663_ (.A(net63),
    .B(net17),
    .Y(_06363_));
 sky130_fd_sc_hd__a22oi_4 _16664_ (.A1(net62),
    .A2(net18),
    .B1(net19),
    .B2(net61),
    .Y(_06364_));
 sky130_fd_sc_hd__a22o_1 _16665_ (.A1(net62),
    .A2(net18),
    .B1(net19),
    .B2(net61),
    .X(_06365_));
 sky130_fd_sc_hd__nand3_4 _16666_ (.A(net61),
    .B(net62),
    .C(net19),
    .Y(_06366_));
 sky130_fd_sc_hd__and4_1 _16667_ (.A(net61),
    .B(net62),
    .C(net18),
    .D(net19),
    .X(_06367_));
 sky130_fd_sc_hd__nand4_1 _16668_ (.A(net61),
    .B(net62),
    .C(net18),
    .D(net19),
    .Y(_06369_));
 sky130_fd_sc_hd__o21bai_1 _16669_ (.A1(_06364_),
    .A2(_06367_),
    .B1_N(_06363_),
    .Y(_06370_));
 sky130_fd_sc_hd__o211ai_2 _16670_ (.A1(_02131_),
    .A2(_06366_),
    .B1(_06365_),
    .C1(_06363_),
    .Y(_06371_));
 sky130_fd_sc_hd__o21ai_2 _16671_ (.A1(_06364_),
    .A2(_06367_),
    .B1(_06363_),
    .Y(_06372_));
 sky130_fd_sc_hd__and4_1 _16672_ (.A(_06365_),
    .B(_06369_),
    .C(net63),
    .D(net17),
    .X(_06373_));
 sky130_fd_sc_hd__o2111ai_4 _16673_ (.A1(_02131_),
    .A2(_06366_),
    .B1(net63),
    .C1(net17),
    .D1(_06365_),
    .Y(_06374_));
 sky130_fd_sc_hd__o21ai_2 _16674_ (.A1(_05657_),
    .A2(_05998_),
    .B1(_05997_),
    .Y(_06375_));
 sky130_fd_sc_hd__o22a_1 _16675_ (.A1(_05639_),
    .A2(_05996_),
    .B1(_05657_),
    .B2(_05998_),
    .X(_06376_));
 sky130_fd_sc_hd__nand3_4 _16676_ (.A(_06370_),
    .B(_06371_),
    .C(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand2_1 _16677_ (.A(_06372_),
    .B(_06375_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand3_4 _16678_ (.A(_06372_),
    .B(_06374_),
    .C(_06375_),
    .Y(_06380_));
 sky130_fd_sc_hd__a21oi_1 _16679_ (.A1(net62),
    .A2(net17),
    .B1(_05977_),
    .Y(_06381_));
 sky130_fd_sc_hd__and3_1 _16680_ (.A(_05976_),
    .B(net17),
    .C(net62),
    .X(_06382_));
 sky130_fd_sc_hd__a31o_1 _16681_ (.A1(_05976_),
    .A2(net17),
    .A3(net62),
    .B1(_05977_),
    .X(_06383_));
 sky130_fd_sc_hd__o2bb2ai_2 _16682_ (.A1_N(_06377_),
    .A2_N(_06380_),
    .B1(_06381_),
    .B2(_05975_),
    .Y(_06384_));
 sky130_fd_sc_hd__o211ai_4 _16683_ (.A1(_05977_),
    .A2(_06382_),
    .B1(_06380_),
    .C1(_06377_),
    .Y(_06385_));
 sky130_fd_sc_hd__o2bb2ai_1 _16684_ (.A1_N(_06377_),
    .A2_N(_06380_),
    .B1(_06382_),
    .B2(_05977_),
    .Y(_06386_));
 sky130_fd_sc_hd__o2111ai_1 _16685_ (.A1(_05621_),
    .A2(_05975_),
    .B1(_05978_),
    .C1(_06377_),
    .D1(_06380_),
    .Y(_06387_));
 sky130_fd_sc_hd__nand2_2 _16686_ (.A(_06386_),
    .B(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__nand2_4 _16687_ (.A(_06384_),
    .B(_06385_),
    .Y(_06389_));
 sky130_fd_sc_hd__a311o_1 _16688_ (.A1(_06333_),
    .A2(_06351_),
    .A3(_06353_),
    .B1(_06360_),
    .C1(_06389_),
    .X(_06391_));
 sky130_fd_sc_hd__a2bb2oi_2 _16689_ (.A1_N(_06022_),
    .A2_N(_06317_),
    .B1(_06358_),
    .B2(_06359_),
    .Y(_06392_));
 sky130_fd_sc_hd__o211ai_4 _16690_ (.A1(_06022_),
    .A2(_06317_),
    .B1(_06354_),
    .C1(_06355_),
    .Y(_06393_));
 sky130_fd_sc_hd__a21oi_2 _16691_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__o2111ai_1 _16692_ (.A1(_06022_),
    .A2(_06317_),
    .B1(_06354_),
    .C1(_06355_),
    .D1(_06389_),
    .Y(_06395_));
 sky130_fd_sc_hd__a31oi_1 _16693_ (.A1(_06319_),
    .A2(_06354_),
    .A3(_06355_),
    .B1(_06389_),
    .Y(_06396_));
 sky130_fd_sc_hd__nand2_2 _16694_ (.A(_06393_),
    .B(_06388_),
    .Y(_06397_));
 sky130_fd_sc_hd__o2bb2ai_4 _16695_ (.A1_N(_06388_),
    .A2_N(_06393_),
    .B1(_06356_),
    .B2(_06360_),
    .Y(_06398_));
 sky130_fd_sc_hd__o211ai_2 _16696_ (.A1(_06356_),
    .A2(_06360_),
    .B1(_06395_),
    .C1(_06397_),
    .Y(_06399_));
 sky130_fd_sc_hd__and3_1 _16697_ (.A(_06362_),
    .B(_06393_),
    .C(_06388_),
    .X(_06400_));
 sky130_fd_sc_hd__a22oi_1 _16698_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06393_),
    .B2(_06362_),
    .Y(_06402_));
 sky130_fd_sc_hd__a22o_1 _16699_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06393_),
    .B2(_06362_),
    .X(_06403_));
 sky130_fd_sc_hd__a221oi_1 _16700_ (.A1(_06032_),
    .A2(_06035_),
    .B1(_06396_),
    .B2(_06362_),
    .C1(_06402_),
    .Y(_06404_));
 sky130_fd_sc_hd__o221ai_4 _16701_ (.A1(_06031_),
    .A2(_06034_),
    .B1(_06361_),
    .B2(_06397_),
    .C1(_06403_),
    .Y(_06405_));
 sky130_fd_sc_hd__o221a_1 _16702_ (.A1(_06362_),
    .A2(_06389_),
    .B1(_06394_),
    .B2(_06398_),
    .C1(_06316_),
    .X(_06406_));
 sky130_fd_sc_hd__o221ai_4 _16703_ (.A1(_06362_),
    .A2(_06389_),
    .B1(_06394_),
    .B2(_06398_),
    .C1(_06316_),
    .Y(_06407_));
 sky130_fd_sc_hd__a31o_1 _16704_ (.A1(_06051_),
    .A2(net14),
    .A3(net34),
    .B1(_06052_),
    .X(_06408_));
 sky130_fd_sc_hd__o21a_1 _16705_ (.A1(_05696_),
    .A2(_06049_),
    .B1(_06053_),
    .X(_06409_));
 sky130_fd_sc_hd__nand2_1 _16706_ (.A(net35),
    .B(net14),
    .Y(_06410_));
 sky130_fd_sc_hd__a22oi_1 _16707_ (.A1(net34),
    .A2(net15),
    .B1(net16),
    .B2(net64),
    .Y(_06411_));
 sky130_fd_sc_hd__a22o_1 _16708_ (.A1(net34),
    .A2(net15),
    .B1(net16),
    .B2(net64),
    .X(_06413_));
 sky130_fd_sc_hd__nand4_4 _16709_ (.A(net64),
    .B(net34),
    .C(net15),
    .D(net16),
    .Y(_06414_));
 sky130_fd_sc_hd__o211ai_2 _16710_ (.A1(_01934_),
    .A2(_02065_),
    .B1(_06413_),
    .C1(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__a21o_1 _16711_ (.A1(_06413_),
    .A2(_06414_),
    .B1(_06410_),
    .X(_06416_));
 sky130_fd_sc_hd__nand4_2 _16712_ (.A(_06413_),
    .B(_06414_),
    .C(net35),
    .D(net14),
    .Y(_06417_));
 sky130_fd_sc_hd__a22o_1 _16713_ (.A1(net35),
    .A2(net14),
    .B1(_06413_),
    .B2(_06414_),
    .X(_06418_));
 sky130_fd_sc_hd__nand3_4 _16714_ (.A(_06408_),
    .B(_06417_),
    .C(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__nand3_4 _16715_ (.A(_06409_),
    .B(_06415_),
    .C(_06416_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand2_1 _16716_ (.A(net38),
    .B(net10),
    .Y(_06421_));
 sky130_fd_sc_hd__nand2_1 _16717_ (.A(net37),
    .B(net13),
    .Y(_06422_));
 sky130_fd_sc_hd__nand2_1 _16718_ (.A(net37),
    .B(net11),
    .Y(_06424_));
 sky130_fd_sc_hd__and4_2 _16719_ (.A(net36),
    .B(net37),
    .C(net11),
    .D(net13),
    .X(_06425_));
 sky130_fd_sc_hd__a22oi_4 _16720_ (.A1(net37),
    .A2(net11),
    .B1(net13),
    .B2(net36),
    .Y(_06426_));
 sky130_fd_sc_hd__a211oi_4 _16721_ (.A1(net38),
    .A2(net10),
    .B1(_06425_),
    .C1(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__o211a_2 _16722_ (.A1(_06425_),
    .A2(_06426_),
    .B1(net38),
    .C1(net10),
    .X(_06428_));
 sky130_fd_sc_hd__o2bb2a_1 _16723_ (.A1_N(net38),
    .A2_N(net10),
    .B1(_06425_),
    .B2(_06426_),
    .X(_06429_));
 sky130_fd_sc_hd__and4bb_1 _16724_ (.A_N(_06425_),
    .B_N(_06426_),
    .C(net38),
    .D(net10),
    .X(_06430_));
 sky130_fd_sc_hd__o2bb2ai_4 _16725_ (.A1_N(_06419_),
    .A2_N(_06420_),
    .B1(_06427_),
    .B2(_06428_),
    .Y(_06431_));
 sky130_fd_sc_hd__o211ai_4 _16726_ (.A1(_06429_),
    .A2(_06430_),
    .B1(_06419_),
    .C1(_06420_),
    .Y(_06432_));
 sky130_fd_sc_hd__o2bb2ai_1 _16727_ (.A1_N(_06419_),
    .A2_N(_06420_),
    .B1(_06429_),
    .B2(_06430_),
    .Y(_06433_));
 sky130_fd_sc_hd__o21ai_4 _16728_ (.A1(_06427_),
    .A2(_06428_),
    .B1(_06420_),
    .Y(_06435_));
 sky130_fd_sc_hd__o211ai_1 _16729_ (.A1(_06427_),
    .A2(_06428_),
    .B1(_06419_),
    .C1(_06420_),
    .Y(_06436_));
 sky130_fd_sc_hd__o21ai_1 _16730_ (.A1(_05988_),
    .A2(_05983_),
    .B1(_05986_),
    .Y(_06437_));
 sky130_fd_sc_hd__a21boi_4 _16731_ (.A1(_05985_),
    .A2(_05987_),
    .B1_N(_05986_),
    .Y(_06438_));
 sky130_fd_sc_hd__nand3_4 _16732_ (.A(_06431_),
    .B(_06432_),
    .C(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__a21oi_4 _16733_ (.A1(_06431_),
    .A2(_06432_),
    .B1(_06438_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand3_1 _16734_ (.A(_06433_),
    .B(_06437_),
    .C(_06436_),
    .Y(_06441_));
 sky130_fd_sc_hd__and3_1 _16735_ (.A(_06058_),
    .B(_06068_),
    .C(_06070_),
    .X(_06442_));
 sky130_fd_sc_hd__o21ai_2 _16736_ (.A1(_06067_),
    .A2(_06069_),
    .B1(_06060_),
    .Y(_06443_));
 sky130_fd_sc_hd__nand2_2 _16737_ (.A(_06058_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__o2bb2a_1 _16738_ (.A1_N(_06439_),
    .A2_N(_06441_),
    .B1(_06442_),
    .B2(_06059_),
    .X(_06446_));
 sky130_fd_sc_hd__o2bb2ai_2 _16739_ (.A1_N(_06439_),
    .A2_N(_06441_),
    .B1(_06442_),
    .B2(_06059_),
    .Y(_06447_));
 sky130_fd_sc_hd__a32oi_4 _16740_ (.A1(_06431_),
    .A2(_06432_),
    .A3(_06438_),
    .B1(_06443_),
    .B2(_06058_),
    .Y(_06448_));
 sky130_fd_sc_hd__nand2_1 _16741_ (.A(_06439_),
    .B(_06444_),
    .Y(_06449_));
 sky130_fd_sc_hd__and3_1 _16742_ (.A(_06439_),
    .B(_06441_),
    .C(_06444_),
    .X(_06450_));
 sky130_fd_sc_hd__o21ai_2 _16743_ (.A1(_06440_),
    .A2(_06449_),
    .B1(_06447_),
    .Y(_06451_));
 sky130_fd_sc_hd__o211ai_2 _16744_ (.A1(_06446_),
    .A2(_06450_),
    .B1(_06405_),
    .C1(_06407_),
    .Y(_06452_));
 sky130_fd_sc_hd__o21bai_1 _16745_ (.A1(_06404_),
    .A2(_06406_),
    .B1_N(_06451_),
    .Y(_06453_));
 sky130_fd_sc_hd__o2bb2ai_2 _16746_ (.A1_N(_06405_),
    .A2_N(_06407_),
    .B1(_06446_),
    .B2(_06450_),
    .Y(_06454_));
 sky130_fd_sc_hd__o2111ai_4 _16747_ (.A1(_06440_),
    .A2(_06449_),
    .B1(_06447_),
    .C1(_06405_),
    .D1(_06407_),
    .Y(_06455_));
 sky130_fd_sc_hd__a21oi_4 _16748_ (.A1(_06454_),
    .A2(_06455_),
    .B1(_06315_),
    .Y(_06457_));
 sky130_fd_sc_hd__o211ai_4 _16749_ (.A1(_06044_),
    .A2(_06314_),
    .B1(_06452_),
    .C1(_06453_),
    .Y(_06458_));
 sky130_fd_sc_hd__nand3_4 _16750_ (.A(_06315_),
    .B(_06454_),
    .C(_06455_),
    .Y(_06459_));
 sky130_fd_sc_hd__and2_1 _16751_ (.A(_06128_),
    .B(_06161_),
    .X(_06460_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(_06128_),
    .B(_06161_),
    .Y(_06461_));
 sky130_fd_sc_hd__a31oi_4 _16753_ (.A1(_06047_),
    .A2(_06076_),
    .A3(_06077_),
    .B1(_06082_),
    .Y(_06462_));
 sky130_fd_sc_hd__a31o_1 _16754_ (.A1(_06047_),
    .A2(_06076_),
    .A3(_06077_),
    .B1(_06085_),
    .X(_06463_));
 sky130_fd_sc_hd__a21oi_1 _16755_ (.A1(net4),
    .A2(net43),
    .B1(_06133_),
    .Y(_06464_));
 sky130_fd_sc_hd__nand2_2 _16756_ (.A(_05764_),
    .B(_06134_),
    .Y(_06465_));
 sky130_fd_sc_hd__nor2_1 _16757_ (.A(_05764_),
    .B(_06131_),
    .Y(_06466_));
 sky130_fd_sc_hd__nand2_1 _16758_ (.A(net4),
    .B(net45),
    .Y(_06468_));
 sky130_fd_sc_hd__nand4_4 _16759_ (.A(net5),
    .B(net6),
    .C(net42),
    .D(net43),
    .Y(_06469_));
 sky130_fd_sc_hd__a22oi_2 _16760_ (.A1(net6),
    .A2(net42),
    .B1(net43),
    .B2(net5),
    .Y(_06470_));
 sky130_fd_sc_hd__a22o_2 _16761_ (.A1(net6),
    .A2(net42),
    .B1(net43),
    .B2(net5),
    .X(_06471_));
 sky130_fd_sc_hd__a22oi_2 _16762_ (.A1(net4),
    .A2(net45),
    .B1(_06469_),
    .B2(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__o2bb2ai_4 _16763_ (.A1_N(_06469_),
    .A2_N(_06471_),
    .B1(_01945_),
    .B2(_02054_),
    .Y(_06473_));
 sky130_fd_sc_hd__nor3b_2 _16764_ (.A(_06470_),
    .B(_06468_),
    .C_N(_06469_),
    .Y(_06474_));
 sky130_fd_sc_hd__nand4_4 _16765_ (.A(_06471_),
    .B(net45),
    .C(net4),
    .D(_06469_),
    .Y(_06475_));
 sky130_fd_sc_hd__a22oi_4 _16766_ (.A1(_06132_),
    .A2(_06465_),
    .B1(_06473_),
    .B2(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__o22ai_4 _16767_ (.A1(_06131_),
    .A2(_06464_),
    .B1(_06472_),
    .B2(_06474_),
    .Y(_06477_));
 sky130_fd_sc_hd__o21ai_1 _16768_ (.A1(_06133_),
    .A2(_06466_),
    .B1(_06473_),
    .Y(_06479_));
 sky130_fd_sc_hd__nand4_4 _16769_ (.A(_06132_),
    .B(_06465_),
    .C(_06473_),
    .D(_06475_),
    .Y(_06480_));
 sky130_fd_sc_hd__nand2_1 _16770_ (.A(net2),
    .B(net47),
    .Y(_06481_));
 sky130_fd_sc_hd__a22oi_2 _16771_ (.A1(net3),
    .A2(net46),
    .B1(net47),
    .B2(net2),
    .Y(_06482_));
 sky130_fd_sc_hd__a22o_1 _16772_ (.A1(net3),
    .A2(net46),
    .B1(net47),
    .B2(net2),
    .X(_06483_));
 sky130_fd_sc_hd__nand2_1 _16773_ (.A(net3),
    .B(net47),
    .Y(_06484_));
 sky130_fd_sc_hd__and4_2 _16774_ (.A(net2),
    .B(net3),
    .C(net46),
    .D(net47),
    .X(_06485_));
 sky130_fd_sc_hd__nand4_2 _16775_ (.A(net2),
    .B(net3),
    .C(net46),
    .D(net47),
    .Y(_06486_));
 sky130_fd_sc_hd__nand2_1 _16776_ (.A(net32),
    .B(net48),
    .Y(_06487_));
 sky130_fd_sc_hd__a22oi_1 _16777_ (.A1(net32),
    .A2(net48),
    .B1(_06483_),
    .B2(_06486_),
    .Y(_06488_));
 sky130_fd_sc_hd__o21ai_1 _16778_ (.A1(_06482_),
    .A2(_06485_),
    .B1(_06487_),
    .Y(_06490_));
 sky130_fd_sc_hd__nor3_1 _16779_ (.A(_06482_),
    .B(_06487_),
    .C(_06485_),
    .Y(_06491_));
 sky130_fd_sc_hd__nand4_1 _16780_ (.A(_06483_),
    .B(_06486_),
    .C(net32),
    .D(net48),
    .Y(_06492_));
 sky130_fd_sc_hd__nor2_1 _16781_ (.A(_06488_),
    .B(_06491_),
    .Y(_06493_));
 sky130_fd_sc_hd__nand2_2 _16782_ (.A(_06490_),
    .B(_06492_),
    .Y(_06494_));
 sky130_fd_sc_hd__a21oi_4 _16783_ (.A1(_06477_),
    .A2(_06480_),
    .B1(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__o221a_2 _16784_ (.A1(_06488_),
    .A2(_06491_),
    .B1(_06474_),
    .B2(_06479_),
    .C1(_06477_),
    .X(_06496_));
 sky130_fd_sc_hd__a21oi_2 _16785_ (.A1(_06477_),
    .A2(_06480_),
    .B1(_06493_),
    .Y(_06497_));
 sky130_fd_sc_hd__and3_2 _16786_ (.A(_06477_),
    .B(_06480_),
    .C(_06493_),
    .X(_06498_));
 sky130_fd_sc_hd__nor2_1 _16787_ (.A(_06495_),
    .B(_06496_),
    .Y(_06499_));
 sky130_fd_sc_hd__nor2_1 _16788_ (.A(_06497_),
    .B(_06498_),
    .Y(_06501_));
 sky130_fd_sc_hd__o21ai_2 _16789_ (.A1(_06119_),
    .A2(_06113_),
    .B1(_06115_),
    .Y(_06502_));
 sky130_fd_sc_hd__a21boi_4 _16790_ (.A1(_06114_),
    .A2(_06118_),
    .B1_N(_06115_),
    .Y(_06503_));
 sky130_fd_sc_hd__a21oi_2 _16791_ (.A1(net7),
    .A2(net40),
    .B1(_06107_),
    .Y(_06504_));
 sky130_fd_sc_hd__and3_2 _16792_ (.A(_06106_),
    .B(net40),
    .C(net7),
    .X(_06505_));
 sky130_fd_sc_hd__a21oi_2 _16793_ (.A1(_06062_),
    .A2(_06063_),
    .B1(_05715_),
    .Y(_06506_));
 sky130_fd_sc_hd__o22ai_4 _16794_ (.A1(_05695_),
    .A2(_06065_),
    .B1(_05715_),
    .B2(_06064_),
    .Y(_06507_));
 sky130_fd_sc_hd__a22oi_4 _16795_ (.A1(net8),
    .A2(net40),
    .B1(net9),
    .B2(net39),
    .Y(_06508_));
 sky130_fd_sc_hd__a22o_1 _16796_ (.A1(net8),
    .A2(net40),
    .B1(net9),
    .B2(net39),
    .X(_06509_));
 sky130_fd_sc_hd__and4_1 _16797_ (.A(net39),
    .B(net8),
    .C(net40),
    .D(net9),
    .X(_06510_));
 sky130_fd_sc_hd__nand4_4 _16798_ (.A(net39),
    .B(net8),
    .C(net40),
    .D(net9),
    .Y(_06512_));
 sky130_fd_sc_hd__o211ai_2 _16799_ (.A1(_01977_),
    .A2(_02010_),
    .B1(_06509_),
    .C1(_06512_),
    .Y(_06513_));
 sky130_fd_sc_hd__o211ai_2 _16800_ (.A1(_06508_),
    .A2(_06510_),
    .B1(net7),
    .C1(net41),
    .Y(_06514_));
 sky130_fd_sc_hd__nand4_4 _16801_ (.A(_06509_),
    .B(_06512_),
    .C(net7),
    .D(net41),
    .Y(_06515_));
 sky130_fd_sc_hd__o22ai_4 _16802_ (.A1(_01977_),
    .A2(_02010_),
    .B1(_06508_),
    .B2(_06510_),
    .Y(_06516_));
 sky130_fd_sc_hd__o211a_2 _16803_ (.A1(_06066_),
    .A2(_06506_),
    .B1(_06515_),
    .C1(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__o211ai_4 _16804_ (.A1(_06066_),
    .A2(_06506_),
    .B1(_06515_),
    .C1(_06516_),
    .Y(_06518_));
 sky130_fd_sc_hd__a21oi_4 _16805_ (.A1(_06515_),
    .A2(_06516_),
    .B1(_06507_),
    .Y(_06519_));
 sky130_fd_sc_hd__nand3b_4 _16806_ (.A_N(_06507_),
    .B(_06513_),
    .C(_06514_),
    .Y(_06520_));
 sky130_fd_sc_hd__o22ai_4 _16807_ (.A1(_06107_),
    .A2(_06505_),
    .B1(_06517_),
    .B2(_06519_),
    .Y(_06521_));
 sky130_fd_sc_hd__o2111ai_4 _16808_ (.A1(_05793_),
    .A2(_06104_),
    .B1(_06108_),
    .C1(_06518_),
    .D1(_06520_),
    .Y(_06523_));
 sky130_fd_sc_hd__o211ai_4 _16809_ (.A1(_06107_),
    .A2(_06505_),
    .B1(_06518_),
    .C1(_06520_),
    .Y(_06524_));
 sky130_fd_sc_hd__o22ai_4 _16810_ (.A1(_06104_),
    .A2(_06504_),
    .B1(_06517_),
    .B2(_06519_),
    .Y(_06525_));
 sky130_fd_sc_hd__a21oi_4 _16811_ (.A1(_06521_),
    .A2(_06523_),
    .B1(_06503_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand3_4 _16812_ (.A(_06525_),
    .B(_06502_),
    .C(_06524_),
    .Y(_06527_));
 sky130_fd_sc_hd__a21oi_2 _16813_ (.A1(_06524_),
    .A2(_06525_),
    .B1(_06502_),
    .Y(_06528_));
 sky130_fd_sc_hd__nand3_4 _16814_ (.A(_06503_),
    .B(_06521_),
    .C(_06523_),
    .Y(_06529_));
 sky130_fd_sc_hd__nand2_1 _16815_ (.A(_06527_),
    .B(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__o211a_4 _16816_ (.A1(_06495_),
    .A2(_06496_),
    .B1(_06527_),
    .C1(_06529_),
    .X(_06531_));
 sky130_fd_sc_hd__o211ai_4 _16817_ (.A1(_06495_),
    .A2(_06496_),
    .B1(_06527_),
    .C1(_06529_),
    .Y(_06532_));
 sky130_fd_sc_hd__a21oi_1 _16818_ (.A1(_06527_),
    .A2(_06529_),
    .B1(_06501_),
    .Y(_06534_));
 sky130_fd_sc_hd__o22ai_4 _16819_ (.A1(_06497_),
    .A2(_06498_),
    .B1(_06526_),
    .B2(_06528_),
    .Y(_06535_));
 sky130_fd_sc_hd__o2bb2ai_2 _16820_ (.A1_N(_06499_),
    .A2_N(_06530_),
    .B1(_06080_),
    .B2(_06085_),
    .Y(_06536_));
 sky130_fd_sc_hd__and3_1 _16821_ (.A(_06463_),
    .B(_06532_),
    .C(_06535_),
    .X(_06537_));
 sky130_fd_sc_hd__o211ai_2 _16822_ (.A1(_06080_),
    .A2(_06085_),
    .B1(_06532_),
    .C1(_06535_),
    .Y(_06538_));
 sky130_fd_sc_hd__a2bb2oi_2 _16823_ (.A1_N(_06078_),
    .A2_N(_06462_),
    .B1(_06532_),
    .B2(_06535_),
    .Y(_06539_));
 sky130_fd_sc_hd__o22ai_4 _16824_ (.A1(_06078_),
    .A2(_06462_),
    .B1(_06531_),
    .B2(_06534_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand2_1 _16825_ (.A(_06461_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__and3_1 _16826_ (.A(_06461_),
    .B(_06538_),
    .C(_06540_),
    .X(_06542_));
 sky130_fd_sc_hd__a21oi_1 _16827_ (.A1(_06538_),
    .A2(_06540_),
    .B1(_06461_),
    .Y(_06543_));
 sky130_fd_sc_hd__a21o_1 _16828_ (.A1(_06538_),
    .A2(_06540_),
    .B1(_06461_),
    .X(_06545_));
 sky130_fd_sc_hd__a21oi_1 _16829_ (.A1(_06538_),
    .A2(_06540_),
    .B1(_06460_),
    .Y(_06546_));
 sky130_fd_sc_hd__a22o_1 _16830_ (.A1(_06128_),
    .A2(_06161_),
    .B1(_06538_),
    .B2(_06540_),
    .X(_06547_));
 sky130_fd_sc_hd__o211ai_4 _16831_ (.A1(_06531_),
    .A2(_06536_),
    .B1(_06460_),
    .C1(_06540_),
    .Y(_06548_));
 sky130_fd_sc_hd__inv_2 _16832_ (.A(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__o21ai_2 _16833_ (.A1(_06537_),
    .A2(_06541_),
    .B1(_06545_),
    .Y(_06550_));
 sky130_fd_sc_hd__o2bb2ai_4 _16834_ (.A1_N(_06458_),
    .A2_N(_06459_),
    .B1(_06542_),
    .B2(_06543_),
    .Y(_06551_));
 sky130_fd_sc_hd__o2111ai_4 _16835_ (.A1(_06537_),
    .A2(_06541_),
    .B1(_06545_),
    .C1(_06459_),
    .D1(_06458_),
    .Y(_06552_));
 sky130_fd_sc_hd__nand4_4 _16836_ (.A(_06458_),
    .B(_06459_),
    .C(_06547_),
    .D(_06548_),
    .Y(_06553_));
 sky130_fd_sc_hd__o2bb2ai_2 _16837_ (.A1_N(_06458_),
    .A2_N(_06459_),
    .B1(_06546_),
    .B2(_06549_),
    .Y(_06554_));
 sky130_fd_sc_hd__o2bb2ai_4 _16838_ (.A1_N(_06175_),
    .A2_N(_06099_),
    .B1(_06098_),
    .B2(_06100_),
    .Y(_06556_));
 sky130_fd_sc_hd__a21boi_2 _16839_ (.A1(_06099_),
    .A2(_06175_),
    .B1_N(_06101_),
    .Y(_06557_));
 sky130_fd_sc_hd__a21oi_1 _16840_ (.A1(_06551_),
    .A2(_06552_),
    .B1(_06556_),
    .Y(_06558_));
 sky130_fd_sc_hd__nand3_2 _16841_ (.A(_06553_),
    .B(_06554_),
    .C(_06557_),
    .Y(_06559_));
 sky130_fd_sc_hd__nand3_4 _16842_ (.A(_06551_),
    .B(_06552_),
    .C(_06556_),
    .Y(_06560_));
 sky130_fd_sc_hd__a21o_1 _16843_ (.A1(_06559_),
    .A2(_06560_),
    .B1(_06312_),
    .X(_06561_));
 sky130_fd_sc_hd__nand3_2 _16844_ (.A(_06312_),
    .B(_06559_),
    .C(_06560_),
    .Y(_06562_));
 sky130_fd_sc_hd__a22o_1 _16845_ (.A1(_06309_),
    .A2(_06311_),
    .B1(_06559_),
    .B2(_06560_),
    .X(_06563_));
 sky130_fd_sc_hd__nand4_2 _16846_ (.A(_06309_),
    .B(_06311_),
    .C(_06559_),
    .D(_06560_),
    .Y(_06564_));
 sky130_fd_sc_hd__a22oi_2 _16847_ (.A1(_06187_),
    .A2(_06189_),
    .B1(_06561_),
    .B2(_06562_),
    .Y(_06565_));
 sky130_fd_sc_hd__nand3_4 _16848_ (.A(_06563_),
    .B(_06564_),
    .C(_06221_),
    .Y(_06567_));
 sky130_fd_sc_hd__a21oi_1 _16849_ (.A1(_06563_),
    .A2(_06564_),
    .B1(_06221_),
    .Y(_06568_));
 sky130_fd_sc_hd__nand3_2 _16850_ (.A(_06222_),
    .B(_06561_),
    .C(_06562_),
    .Y(_06569_));
 sky130_fd_sc_hd__and3_1 _16851_ (.A(_05586_),
    .B(_05591_),
    .C(_05957_),
    .X(_06570_));
 sky130_fd_sc_hd__a31o_1 _16852_ (.A1(_05882_),
    .A2(_05953_),
    .A3(_05955_),
    .B1(_05961_),
    .X(_06571_));
 sky130_fd_sc_hd__a31o_1 _16853_ (.A1(_05586_),
    .A2(_05590_),
    .A3(_05957_),
    .B1(_05958_),
    .X(_06572_));
 sky130_fd_sc_hd__o22ai_2 _16854_ (.A1(_05956_),
    .A2(_05961_),
    .B1(_06565_),
    .B2(_06568_),
    .Y(_06573_));
 sky130_fd_sc_hd__o2111ai_4 _16855_ (.A1(_05880_),
    .A2(_05958_),
    .B1(_06567_),
    .C1(_06569_),
    .D1(_05957_),
    .Y(_06574_));
 sky130_fd_sc_hd__o2bb2ai_1 _16856_ (.A1_N(_06567_),
    .A2_N(_06569_),
    .B1(_06570_),
    .B2(_05958_),
    .Y(_06575_));
 sky130_fd_sc_hd__o211ai_2 _16857_ (.A1(_05956_),
    .A2(_05961_),
    .B1(_06567_),
    .C1(_06569_),
    .Y(_06576_));
 sky130_fd_sc_hd__nand3_4 _16858_ (.A(_06573_),
    .B(_06574_),
    .C(_06219_),
    .Y(_06578_));
 sky130_fd_sc_hd__and3_1 _16859_ (.A(_06220_),
    .B(_06575_),
    .C(_06576_),
    .X(_06579_));
 sky130_fd_sc_hd__nand3_1 _16860_ (.A(_06220_),
    .B(_06575_),
    .C(_06576_),
    .Y(_06580_));
 sky130_fd_sc_hd__a21o_1 _16861_ (.A1(_06578_),
    .A2(_06580_),
    .B1(_05910_),
    .X(_06581_));
 sky130_fd_sc_hd__o211ai_1 _16862_ (.A1(_05908_),
    .A2(_05903_),
    .B1(_06580_),
    .C1(_06578_),
    .Y(_06582_));
 sky130_fd_sc_hd__o2bb2ai_1 _16863_ (.A1_N(_06578_),
    .A2_N(_06580_),
    .B1(_05903_),
    .B2(_05908_),
    .Y(_06583_));
 sky130_fd_sc_hd__a31o_1 _16864_ (.A1(_06573_),
    .A2(_06574_),
    .A3(_06219_),
    .B1(_05910_),
    .X(_06584_));
 sky130_fd_sc_hd__nand3_1 _16865_ (.A(_06218_),
    .B(_06581_),
    .C(_06582_),
    .Y(_06585_));
 sky130_fd_sc_hd__o221ai_4 _16866_ (.A1(_06205_),
    .A2(_06208_),
    .B1(_06579_),
    .B2(_06584_),
    .C1(_06583_),
    .Y(_06586_));
 sky130_fd_sc_hd__and2_1 _16867_ (.A(_06585_),
    .B(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__o211a_2 _16868_ (.A1(_06209_),
    .A2(_06213_),
    .B1(_05870_),
    .C1(_06212_),
    .X(_06589_));
 sky130_fd_sc_hd__nand4_1 _16869_ (.A(_05514_),
    .B(_05870_),
    .C(_06212_),
    .D(_06214_),
    .Y(_06590_));
 sky130_fd_sc_hd__nand4_4 _16870_ (.A(_04500_),
    .B(_04502_),
    .C(_04818_),
    .D(_04819_),
    .Y(_06591_));
 sky130_fd_sc_hd__o21bai_4 _16871_ (.A1(_04506_),
    .A2(_06591_),
    .B1_N(_05164_),
    .Y(_06592_));
 sky130_fd_sc_hd__nand4_1 _16872_ (.A(_06212_),
    .B(_06214_),
    .C(_05870_),
    .D(_05871_),
    .Y(_06593_));
 sky130_fd_sc_hd__o211ai_1 _16873_ (.A1(_05866_),
    .A2(_05869_),
    .B1(_06210_),
    .C1(_06211_),
    .Y(_06594_));
 sky130_fd_sc_hd__nand2_1 _16874_ (.A(_06593_),
    .B(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__a31oi_4 _16875_ (.A1(_05514_),
    .A2(_06589_),
    .A3(_06592_),
    .B1(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__nor3_4 _16876_ (.A(_03862_),
    .B(_04174_),
    .C(_06591_),
    .Y(_06597_));
 sky130_fd_sc_hd__nand4_4 _16877_ (.A(_03869_),
    .B(_05514_),
    .C(_06589_),
    .D(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__nand4b_4 _16878_ (.A_N(_06590_),
    .B(_01763_),
    .C(_03864_),
    .D(_06597_),
    .Y(_06600_));
 sky130_fd_sc_hd__nand3_4 _16879_ (.A(_06596_),
    .B(_06598_),
    .C(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__xor2_1 _16880_ (.A(_06587_),
    .B(_06601_),
    .X(net90));
 sky130_fd_sc_hd__a31oi_2 _16881_ (.A1(_06223_),
    .A2(_06304_),
    .A3(_06305_),
    .B1(_06310_),
    .Y(_06602_));
 sky130_fd_sc_hd__a31o_1 _16882_ (.A1(_06223_),
    .A2(_06304_),
    .A3(_06305_),
    .B1(_06310_),
    .X(_06603_));
 sky130_fd_sc_hd__a32oi_4 _16883_ (.A1(_06551_),
    .A2(_06556_),
    .A3(_06552_),
    .B1(_06309_),
    .B2(_06311_),
    .Y(_06604_));
 sky130_fd_sc_hd__a32oi_4 _16884_ (.A1(_06553_),
    .A2(_06554_),
    .A3(_06557_),
    .B1(_06560_),
    .B2(_06312_),
    .Y(_06605_));
 sky130_fd_sc_hd__a32o_1 _16885_ (.A1(_06553_),
    .A2(_06554_),
    .A3(_06557_),
    .B1(_06560_),
    .B2(_06312_),
    .X(_06606_));
 sky130_fd_sc_hd__o2bb2ai_2 _16886_ (.A1_N(_06286_),
    .A2_N(_06283_),
    .B1(_06281_),
    .B2(_06277_),
    .Y(_06607_));
 sky130_fd_sc_hd__o21a_1 _16887_ (.A1(_01791_),
    .A2(_02207_),
    .B1(_06274_),
    .X(_06608_));
 sky130_fd_sc_hd__a31o_1 _16888_ (.A1(_06271_),
    .A2(net54),
    .A3(net26),
    .B1(_06273_),
    .X(_06610_));
 sky130_fd_sc_hd__nand2_1 _16889_ (.A(net27),
    .B(net54),
    .Y(_06611_));
 sky130_fd_sc_hd__nand2_2 _16890_ (.A(net29),
    .B(net52),
    .Y(_06612_));
 sky130_fd_sc_hd__and4_1 _16891_ (.A(net28),
    .B(net29),
    .C(net52),
    .D(net53),
    .X(_06613_));
 sky130_fd_sc_hd__nand4_2 _16892_ (.A(net28),
    .B(net29),
    .C(net52),
    .D(net53),
    .Y(_06614_));
 sky130_fd_sc_hd__a22oi_1 _16893_ (.A1(net29),
    .A2(net52),
    .B1(net53),
    .B2(net28),
    .Y(_06615_));
 sky130_fd_sc_hd__a22o_2 _16894_ (.A1(net29),
    .A2(net52),
    .B1(net53),
    .B2(net28),
    .X(_06616_));
 sky130_fd_sc_hd__a22oi_2 _16895_ (.A1(net27),
    .A2(net54),
    .B1(_06614_),
    .B2(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__o21ai_1 _16896_ (.A1(_06613_),
    .A2(_06615_),
    .B1(_06611_),
    .Y(_06618_));
 sky130_fd_sc_hd__and4_2 _16897_ (.A(_06616_),
    .B(net54),
    .C(net27),
    .D(_06614_),
    .X(_06619_));
 sky130_fd_sc_hd__nand4_1 _16898_ (.A(_06616_),
    .B(net54),
    .C(net27),
    .D(_06614_),
    .Y(_06621_));
 sky130_fd_sc_hd__a21oi_1 _16899_ (.A1(_06618_),
    .A2(_06621_),
    .B1(_06610_),
    .Y(_06622_));
 sky130_fd_sc_hd__o22ai_4 _16900_ (.A1(_06270_),
    .A2(_06608_),
    .B1(_06617_),
    .B2(_06619_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand2_1 _16901_ (.A(_06610_),
    .B(_06618_),
    .Y(_06624_));
 sky130_fd_sc_hd__nand3_1 _16902_ (.A(_06610_),
    .B(_06618_),
    .C(_06621_),
    .Y(_06625_));
 sky130_fd_sc_hd__nand2_1 _16903_ (.A(net26),
    .B(net56),
    .Y(_06626_));
 sky130_fd_sc_hd__and4b_1 _16904_ (.A_N(net23),
    .B(net56),
    .C(net57),
    .D(net26),
    .X(_06627_));
 sky130_fd_sc_hd__or4_2 _16905_ (.A(net23),
    .B(_02229_),
    .C(_02240_),
    .D(_01791_),
    .X(_06628_));
 sky130_fd_sc_hd__a22oi_1 _16906_ (.A1(net26),
    .A2(net56),
    .B1(_01802_),
    .B2(net57),
    .Y(_06629_));
 sky130_fd_sc_hd__nor2_1 _16907_ (.A(_06627_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__or2_1 _16908_ (.A(_06627_),
    .B(_06629_),
    .X(_06632_));
 sky130_fd_sc_hd__a21oi_2 _16909_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_06630_),
    .Y(_06633_));
 sky130_fd_sc_hd__a21o_1 _16910_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_06630_),
    .X(_06634_));
 sky130_fd_sc_hd__and3_1 _16911_ (.A(_06623_),
    .B(_06625_),
    .C(_06630_),
    .X(_06635_));
 sky130_fd_sc_hd__o211ai_2 _16912_ (.A1(_06619_),
    .A2(_06624_),
    .B1(_06630_),
    .C1(_06623_),
    .Y(_06636_));
 sky130_fd_sc_hd__o221a_1 _16913_ (.A1(_06277_),
    .A2(_06281_),
    .B1(_06633_),
    .B2(_06635_),
    .C1(_06288_),
    .X(_06637_));
 sky130_fd_sc_hd__o21bai_4 _16914_ (.A1(_06633_),
    .A2(_06635_),
    .B1_N(_06607_),
    .Y(_06638_));
 sky130_fd_sc_hd__nand3_4 _16915_ (.A(_06607_),
    .B(_06634_),
    .C(_06636_),
    .Y(_06639_));
 sky130_fd_sc_hd__a21oi_2 _16916_ (.A1(_06638_),
    .A2(_06639_),
    .B1(_06284_),
    .Y(_06640_));
 sky130_fd_sc_hd__a21o_1 _16917_ (.A1(_06638_),
    .A2(_06639_),
    .B1(_06284_),
    .X(_06641_));
 sky130_fd_sc_hd__and3_1 _16918_ (.A(_06638_),
    .B(_06639_),
    .C(_06284_),
    .X(_06643_));
 sky130_fd_sc_hd__nand3_1 _16919_ (.A(_06638_),
    .B(_06639_),
    .C(_06284_),
    .Y(_06644_));
 sky130_fd_sc_hd__o311a_1 _16920_ (.A1(net12),
    .A2(_02240_),
    .A3(_05884_),
    .B1(_06638_),
    .C1(_06639_),
    .X(_06645_));
 sky130_fd_sc_hd__a21boi_1 _16921_ (.A1(_06638_),
    .A2(_06639_),
    .B1_N(_06284_),
    .Y(_06646_));
 sky130_fd_sc_hd__a21oi_1 _16922_ (.A1(_06254_),
    .A2(_06229_),
    .B1(_06228_),
    .Y(_06647_));
 sky130_fd_sc_hd__a31o_2 _16923_ (.A1(_06233_),
    .A2(_06243_),
    .A3(_06244_),
    .B1(_06250_),
    .X(_06648_));
 sky130_fd_sc_hd__nand2_1 _16924_ (.A(_06477_),
    .B(_06493_),
    .Y(_06649_));
 sky130_fd_sc_hd__o22ai_2 _16925_ (.A1(_06474_),
    .A2(_06479_),
    .B1(_06494_),
    .B2(_06476_),
    .Y(_06650_));
 sky130_fd_sc_hd__and3_1 _16926_ (.A(_06238_),
    .B(net51),
    .C(net29),
    .X(_06651_));
 sky130_fd_sc_hd__a31o_1 _16927_ (.A1(_06238_),
    .A2(net51),
    .A3(net29),
    .B1(_06239_),
    .X(_06652_));
 sky130_fd_sc_hd__a21oi_2 _16928_ (.A1(_06142_),
    .A2(_06481_),
    .B1(_06487_),
    .Y(_06654_));
 sky130_fd_sc_hd__o21ai_2 _16929_ (.A1(_06487_),
    .A2(_06482_),
    .B1(_06486_),
    .Y(_06655_));
 sky130_fd_sc_hd__nand2_1 _16930_ (.A(net30),
    .B(net51),
    .Y(_06656_));
 sky130_fd_sc_hd__a22oi_4 _16931_ (.A1(net32),
    .A2(net49),
    .B1(net50),
    .B2(net31),
    .Y(_06657_));
 sky130_fd_sc_hd__a22o_1 _16932_ (.A1(net32),
    .A2(net49),
    .B1(net50),
    .B2(net31),
    .X(_06658_));
 sky130_fd_sc_hd__and4_4 _16933_ (.A(net31),
    .B(net32),
    .C(net49),
    .D(net50),
    .X(_06659_));
 sky130_fd_sc_hd__nand4_4 _16934_ (.A(net31),
    .B(net32),
    .C(net49),
    .D(net50),
    .Y(_06660_));
 sky130_fd_sc_hd__o211ai_2 _16935_ (.A1(_01868_),
    .A2(_02152_),
    .B1(_06658_),
    .C1(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__o21bai_2 _16936_ (.A1(_06657_),
    .A2(_06659_),
    .B1_N(_06656_),
    .Y(_06662_));
 sky130_fd_sc_hd__nand4_4 _16937_ (.A(_06658_),
    .B(_06660_),
    .C(net30),
    .D(net51),
    .Y(_06663_));
 sky130_fd_sc_hd__o22ai_4 _16938_ (.A1(_01868_),
    .A2(_02152_),
    .B1(_06657_),
    .B2(_06659_),
    .Y(_06665_));
 sky130_fd_sc_hd__o211a_2 _16939_ (.A1(_06485_),
    .A2(_06654_),
    .B1(_06663_),
    .C1(_06665_),
    .X(_06666_));
 sky130_fd_sc_hd__o211ai_4 _16940_ (.A1(_06485_),
    .A2(_06654_),
    .B1(_06663_),
    .C1(_06665_),
    .Y(_06667_));
 sky130_fd_sc_hd__a21oi_4 _16941_ (.A1(_06663_),
    .A2(_06665_),
    .B1(_06655_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand3b_4 _16942_ (.A_N(_06655_),
    .B(_06661_),
    .C(_06662_),
    .Y(_06669_));
 sky130_fd_sc_hd__nor2_1 _16943_ (.A(_06666_),
    .B(_06668_),
    .Y(_06670_));
 sky130_fd_sc_hd__o21a_1 _16944_ (.A1(_06239_),
    .A2(_06651_),
    .B1(_06669_),
    .X(_06671_));
 sky130_fd_sc_hd__and3_1 _16945_ (.A(_06669_),
    .B(_06652_),
    .C(_06667_),
    .X(_06672_));
 sky130_fd_sc_hd__a2bb2oi_1 _16946_ (.A1_N(_06239_),
    .A2_N(_06651_),
    .B1(_06667_),
    .B2(_06669_),
    .Y(_06673_));
 sky130_fd_sc_hd__o22ai_4 _16947_ (.A1(_06239_),
    .A2(_06651_),
    .B1(_06666_),
    .B2(_06668_),
    .Y(_06674_));
 sky130_fd_sc_hd__o2111a_1 _16948_ (.A1(_06235_),
    .A2(_06237_),
    .B1(_06240_),
    .C1(_06667_),
    .D1(_06669_),
    .X(_06676_));
 sky130_fd_sc_hd__o2111ai_4 _16949_ (.A1(_06235_),
    .A2(_06237_),
    .B1(_06240_),
    .C1(_06667_),
    .D1(_06669_),
    .Y(_06677_));
 sky130_fd_sc_hd__o2bb2ai_2 _16950_ (.A1_N(_06480_),
    .A2_N(_06649_),
    .B1(_06652_),
    .B2(_06670_),
    .Y(_06678_));
 sky130_fd_sc_hd__a22oi_4 _16951_ (.A1(_06480_),
    .A2(_06649_),
    .B1(_06674_),
    .B2(_06677_),
    .Y(_06679_));
 sky130_fd_sc_hd__o21ai_1 _16952_ (.A1(_06673_),
    .A2(_06676_),
    .B1(_06650_),
    .Y(_06680_));
 sky130_fd_sc_hd__nor3_2 _16953_ (.A(_06650_),
    .B(_06673_),
    .C(_06676_),
    .Y(_06681_));
 sky130_fd_sc_hd__o2111ai_4 _16954_ (.A1(_06494_),
    .A2(_06476_),
    .B1(_06480_),
    .C1(_06674_),
    .D1(_06677_),
    .Y(_06682_));
 sky130_fd_sc_hd__o221ai_4 _16955_ (.A1(_06245_),
    .A2(_06250_),
    .B1(_06672_),
    .B2(_06678_),
    .C1(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__o21bai_4 _16956_ (.A1(_06679_),
    .A2(_06681_),
    .B1_N(_06648_),
    .Y(_06684_));
 sky130_fd_sc_hd__o22ai_4 _16957_ (.A1(_06245_),
    .A2(_06250_),
    .B1(_06679_),
    .B2(_06681_),
    .Y(_06685_));
 sky130_fd_sc_hd__nand3b_2 _16958_ (.A_N(_06648_),
    .B(_06680_),
    .C(_06682_),
    .Y(_06687_));
 sky130_fd_sc_hd__a22oi_4 _16959_ (.A1(_06256_),
    .A2(_06261_),
    .B1(_06685_),
    .B2(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__o211ai_4 _16960_ (.A1(_06255_),
    .A2(_06260_),
    .B1(_06683_),
    .C1(_06684_),
    .Y(_06689_));
 sky130_fd_sc_hd__a2bb2oi_4 _16961_ (.A1_N(_06257_),
    .A2_N(_06647_),
    .B1(_06683_),
    .B2(_06684_),
    .Y(_06690_));
 sky130_fd_sc_hd__o2111ai_4 _16962_ (.A1(_06227_),
    .A2(_06257_),
    .B1(_06685_),
    .C1(_06687_),
    .D1(_06256_),
    .Y(_06691_));
 sky130_fd_sc_hd__o22ai_2 _16963_ (.A1(_06645_),
    .A2(_06646_),
    .B1(_06688_),
    .B2(_06690_),
    .Y(_06692_));
 sky130_fd_sc_hd__o211ai_2 _16964_ (.A1(_06640_),
    .A2(_06643_),
    .B1(_06689_),
    .C1(_06691_),
    .Y(_06693_));
 sky130_fd_sc_hd__o22ai_2 _16965_ (.A1(_06640_),
    .A2(_06643_),
    .B1(_06688_),
    .B2(_06690_),
    .Y(_06694_));
 sky130_fd_sc_hd__and3_1 _16966_ (.A(_06641_),
    .B(_06644_),
    .C(_06691_),
    .X(_06695_));
 sky130_fd_sc_hd__o211ai_2 _16967_ (.A1(_06645_),
    .A2(_06646_),
    .B1(_06689_),
    .C1(_06691_),
    .Y(_06696_));
 sky130_fd_sc_hd__a31oi_2 _16968_ (.A1(_06463_),
    .A2(_06532_),
    .A3(_06535_),
    .B1(_06461_),
    .Y(_06698_));
 sky130_fd_sc_hd__o22ai_2 _16969_ (.A1(_06536_),
    .A2(_06531_),
    .B1(_06460_),
    .B2(_06539_),
    .Y(_06699_));
 sky130_fd_sc_hd__o211ai_4 _16970_ (.A1(_06539_),
    .A2(_06698_),
    .B1(_06693_),
    .C1(_06692_),
    .Y(_06700_));
 sky130_fd_sc_hd__and3_2 _16971_ (.A(_06694_),
    .B(_06699_),
    .C(_06696_),
    .X(_06701_));
 sky130_fd_sc_hd__nand3_2 _16972_ (.A(_06694_),
    .B(_06699_),
    .C(_06696_),
    .Y(_06702_));
 sky130_fd_sc_hd__a21bo_1 _16973_ (.A1(_06265_),
    .A2(_06300_),
    .B1_N(_06264_),
    .X(_06703_));
 sky130_fd_sc_hd__a21o_2 _16974_ (.A1(_06700_),
    .A2(_06702_),
    .B1(_06703_),
    .X(_06704_));
 sky130_fd_sc_hd__nand2_2 _16975_ (.A(_06700_),
    .B(_06703_),
    .Y(_06705_));
 sky130_fd_sc_hd__and3_1 _16976_ (.A(_06700_),
    .B(_06702_),
    .C(_06703_),
    .X(_06706_));
 sky130_fd_sc_hd__nand3_2 _16977_ (.A(_06700_),
    .B(_06702_),
    .C(_06703_),
    .Y(_06707_));
 sky130_fd_sc_hd__o21ai_4 _16978_ (.A1(_06701_),
    .A2(_06705_),
    .B1(_06704_),
    .Y(_06709_));
 sky130_fd_sc_hd__a31oi_4 _16979_ (.A1(_06459_),
    .A2(_06547_),
    .A3(_06548_),
    .B1(_06457_),
    .Y(_06710_));
 sky130_fd_sc_hd__o21a_1 _16980_ (.A1(_01977_),
    .A2(_02010_),
    .B1(_06512_),
    .X(_06711_));
 sky130_fd_sc_hd__a31o_1 _16981_ (.A1(_06509_),
    .A2(net41),
    .A3(net7),
    .B1(_06510_),
    .X(_06712_));
 sky130_fd_sc_hd__a21oi_2 _16982_ (.A1(_06065_),
    .A2(_06424_),
    .B1(_06421_),
    .Y(_06713_));
 sky130_fd_sc_hd__o22ai_1 _16983_ (.A1(_06063_),
    .A2(_06422_),
    .B1(_06421_),
    .B2(_06426_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(net8),
    .B(net41),
    .Y(_06715_));
 sky130_fd_sc_hd__a22oi_4 _16985_ (.A1(net40),
    .A2(net9),
    .B1(net10),
    .B2(net39),
    .Y(_06716_));
 sky130_fd_sc_hd__a22o_1 _16986_ (.A1(net40),
    .A2(net9),
    .B1(net10),
    .B2(net39),
    .X(_06717_));
 sky130_fd_sc_hd__and4_2 _16987_ (.A(net39),
    .B(net40),
    .C(net9),
    .D(net10),
    .X(_06718_));
 sky130_fd_sc_hd__nand4_4 _16988_ (.A(net39),
    .B(net40),
    .C(net9),
    .D(net10),
    .Y(_06720_));
 sky130_fd_sc_hd__o211ai_1 _16989_ (.A1(_01988_),
    .A2(_02010_),
    .B1(_06717_),
    .C1(_06720_),
    .Y(_06721_));
 sky130_fd_sc_hd__o21bai_1 _16990_ (.A1(_06716_),
    .A2(_06718_),
    .B1_N(_06715_),
    .Y(_06722_));
 sky130_fd_sc_hd__nand4_2 _16991_ (.A(_06717_),
    .B(_06720_),
    .C(net8),
    .D(net41),
    .Y(_06723_));
 sky130_fd_sc_hd__o22ai_4 _16992_ (.A1(_01988_),
    .A2(_02010_),
    .B1(_06716_),
    .B2(_06718_),
    .Y(_06724_));
 sky130_fd_sc_hd__o211a_1 _16993_ (.A1(_06425_),
    .A2(_06713_),
    .B1(_06723_),
    .C1(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__o211ai_4 _16994_ (.A1(_06425_),
    .A2(_06713_),
    .B1(_06723_),
    .C1(_06724_),
    .Y(_06726_));
 sky130_fd_sc_hd__a21oi_1 _16995_ (.A1(_06723_),
    .A2(_06724_),
    .B1(_06714_),
    .Y(_06727_));
 sky130_fd_sc_hd__nand3b_2 _16996_ (.A_N(_06714_),
    .B(_06721_),
    .C(_06722_),
    .Y(_06728_));
 sky130_fd_sc_hd__nand3_4 _16997_ (.A(_06728_),
    .B(_06712_),
    .C(_06726_),
    .Y(_06729_));
 sky130_fd_sc_hd__o22ai_4 _16998_ (.A1(_06508_),
    .A2(_06711_),
    .B1(_06725_),
    .B2(_06727_),
    .Y(_06731_));
 sky130_fd_sc_hd__o211a_1 _16999_ (.A1(_05793_),
    .A2(_06104_),
    .B1(_06108_),
    .C1(_06518_),
    .X(_06732_));
 sky130_fd_sc_hd__o21ai_2 _17000_ (.A1(_06104_),
    .A2(_06504_),
    .B1(_06518_),
    .Y(_06733_));
 sky130_fd_sc_hd__o2bb2ai_4 _17001_ (.A1_N(_06729_),
    .A2_N(_06731_),
    .B1(_06732_),
    .B2(_06519_),
    .Y(_06734_));
 sky130_fd_sc_hd__nand4_4 _17002_ (.A(_06520_),
    .B(_06729_),
    .C(_06731_),
    .D(_06733_),
    .Y(_06735_));
 sky130_fd_sc_hd__o21ai_2 _17003_ (.A1(_06468_),
    .A2(_06470_),
    .B1(_06469_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_1 _17004_ (.A(net5),
    .B(net45),
    .Y(_06737_));
 sky130_fd_sc_hd__a22oi_4 _17005_ (.A1(net7),
    .A2(net42),
    .B1(net43),
    .B2(net6),
    .Y(_06738_));
 sky130_fd_sc_hd__a22o_1 _17006_ (.A1(net7),
    .A2(net42),
    .B1(net43),
    .B2(net6),
    .X(_06739_));
 sky130_fd_sc_hd__and4_1 _17007_ (.A(net6),
    .B(net7),
    .C(net42),
    .D(net43),
    .X(_06740_));
 sky130_fd_sc_hd__nand4_2 _17008_ (.A(net6),
    .B(net7),
    .C(net42),
    .D(net43),
    .Y(_06742_));
 sky130_fd_sc_hd__a22oi_2 _17009_ (.A1(net5),
    .A2(net45),
    .B1(_06739_),
    .B2(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__o21ai_1 _17010_ (.A1(_06738_),
    .A2(_06740_),
    .B1(_06737_),
    .Y(_06744_));
 sky130_fd_sc_hd__a41o_1 _17011_ (.A1(net6),
    .A2(net7),
    .A3(net42),
    .A4(net43),
    .B1(_06737_),
    .X(_06745_));
 sky130_fd_sc_hd__nor3_1 _17012_ (.A(_06737_),
    .B(_06738_),
    .C(_06740_),
    .Y(_06746_));
 sky130_fd_sc_hd__o21bai_4 _17013_ (.A1(_06743_),
    .A2(_06746_),
    .B1_N(_06736_),
    .Y(_06747_));
 sky130_fd_sc_hd__o211ai_4 _17014_ (.A1(_06738_),
    .A2(_06745_),
    .B1(_06736_),
    .C1(_06744_),
    .Y(_06748_));
 sky130_fd_sc_hd__nand2_1 _17015_ (.A(net2),
    .B(net48),
    .Y(_06749_));
 sky130_fd_sc_hd__nand2_1 _17016_ (.A(net4),
    .B(net46),
    .Y(_06750_));
 sky130_fd_sc_hd__and4_2 _17017_ (.A(net3),
    .B(net4),
    .C(net46),
    .D(net47),
    .X(_06751_));
 sky130_fd_sc_hd__nand4_2 _17018_ (.A(net3),
    .B(net4),
    .C(net46),
    .D(net47),
    .Y(_06753_));
 sky130_fd_sc_hd__a22oi_2 _17019_ (.A1(net4),
    .A2(net46),
    .B1(net47),
    .B2(net3),
    .Y(_06754_));
 sky130_fd_sc_hd__a22o_1 _17020_ (.A1(net4),
    .A2(net46),
    .B1(net47),
    .B2(net3),
    .X(_06755_));
 sky130_fd_sc_hd__o311a_1 _17021_ (.A1(_01945_),
    .A2(_02087_),
    .A3(_06142_),
    .B1(_06749_),
    .C1(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__o211ai_2 _17022_ (.A1(_01901_),
    .A2(_02109_),
    .B1(_06753_),
    .C1(_06755_),
    .Y(_06757_));
 sky130_fd_sc_hd__o211a_1 _17023_ (.A1(_06751_),
    .A2(_06754_),
    .B1(net2),
    .C1(net48),
    .X(_06758_));
 sky130_fd_sc_hd__o21bai_2 _17024_ (.A1(_06751_),
    .A2(_06754_),
    .B1_N(_06749_),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_2 _17025_ (.A(_06757_),
    .B(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__and3_2 _17026_ (.A(_06747_),
    .B(_06748_),
    .C(_06760_),
    .X(_06761_));
 sky130_fd_sc_hd__a21oi_4 _17027_ (.A1(_06747_),
    .A2(_06748_),
    .B1(_06760_),
    .Y(_06762_));
 sky130_fd_sc_hd__nand4_2 _17028_ (.A(_06747_),
    .B(_06748_),
    .C(_06757_),
    .D(_06759_),
    .Y(_06764_));
 sky130_fd_sc_hd__inv_2 _17029_ (.A(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__o2bb2ai_2 _17030_ (.A1_N(_06747_),
    .A2_N(_06748_),
    .B1(_06756_),
    .B2(_06758_),
    .Y(_06766_));
 sky130_fd_sc_hd__inv_2 _17031_ (.A(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__nand2_2 _17032_ (.A(_06764_),
    .B(_06766_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand3_2 _17033_ (.A(_06734_),
    .B(_06768_),
    .C(_06735_),
    .Y(_06769_));
 sky130_fd_sc_hd__o2bb2ai_4 _17034_ (.A1_N(_06734_),
    .A2_N(_06735_),
    .B1(_06761_),
    .B2(_06762_),
    .Y(_06770_));
 sky130_fd_sc_hd__o211ai_4 _17035_ (.A1(_06761_),
    .A2(_06762_),
    .B1(_06734_),
    .C1(_06735_),
    .Y(_06771_));
 sky130_fd_sc_hd__o2bb2ai_4 _17036_ (.A1_N(_06734_),
    .A2_N(_06735_),
    .B1(_06765_),
    .B2(_06767_),
    .Y(_06772_));
 sky130_fd_sc_hd__a21oi_4 _17037_ (.A1(_06439_),
    .A2(_06444_),
    .B1(_06440_),
    .Y(_06773_));
 sky130_fd_sc_hd__a32o_1 _17038_ (.A1(_06433_),
    .A2(_06436_),
    .A3(_06437_),
    .B1(_06439_),
    .B2(_06444_),
    .X(_06775_));
 sky130_fd_sc_hd__and3_1 _17039_ (.A(_06771_),
    .B(_06772_),
    .C(_06773_),
    .X(_06776_));
 sky130_fd_sc_hd__nand3_2 _17040_ (.A(_06771_),
    .B(_06772_),
    .C(_06773_),
    .Y(_06777_));
 sky130_fd_sc_hd__and3_1 _17041_ (.A(_06769_),
    .B(_06770_),
    .C(_06775_),
    .X(_06778_));
 sky130_fd_sc_hd__o211ai_4 _17042_ (.A1(_06440_),
    .A2(_06448_),
    .B1(_06769_),
    .C1(_06770_),
    .Y(_06779_));
 sky130_fd_sc_hd__a21oi_4 _17043_ (.A1(_06501_),
    .A2(_06529_),
    .B1(_06526_),
    .Y(_06780_));
 sky130_fd_sc_hd__o21ai_2 _17044_ (.A1(_06499_),
    .A2(_06528_),
    .B1(_06527_),
    .Y(_06781_));
 sky130_fd_sc_hd__a31o_1 _17045_ (.A1(_06771_),
    .A2(_06772_),
    .A3(_06773_),
    .B1(_06780_),
    .X(_06782_));
 sky130_fd_sc_hd__o211ai_4 _17046_ (.A1(_06526_),
    .A2(_06531_),
    .B1(_06777_),
    .C1(_06779_),
    .Y(_06783_));
 sky130_fd_sc_hd__a21o_1 _17047_ (.A1(_06777_),
    .A2(_06779_),
    .B1(_06781_),
    .X(_06784_));
 sky130_fd_sc_hd__a21oi_2 _17048_ (.A1(_06777_),
    .A2(_06779_),
    .B1(_06780_),
    .Y(_06786_));
 sky130_fd_sc_hd__and3_1 _17049_ (.A(_06777_),
    .B(_06779_),
    .C(_06780_),
    .X(_06787_));
 sky130_fd_sc_hd__o21ai_2 _17050_ (.A1(_06778_),
    .A2(_06782_),
    .B1(_06784_),
    .Y(_06788_));
 sky130_fd_sc_hd__o21ai_1 _17051_ (.A1(_06410_),
    .A2(_06411_),
    .B1(_06414_),
    .Y(_06789_));
 sky130_fd_sc_hd__o31a_2 _17052_ (.A1(_01934_),
    .A2(_02065_),
    .A3(_06411_),
    .B1(_06414_),
    .X(_06790_));
 sky130_fd_sc_hd__nand2_1 _17053_ (.A(net35),
    .B(net15),
    .Y(_06791_));
 sky130_fd_sc_hd__a22oi_2 _17054_ (.A1(net34),
    .A2(net16),
    .B1(net17),
    .B2(net64),
    .Y(_06792_));
 sky130_fd_sc_hd__a22o_1 _17055_ (.A1(net34),
    .A2(net16),
    .B1(net17),
    .B2(net64),
    .X(_06793_));
 sky130_fd_sc_hd__and4_1 _17056_ (.A(net64),
    .B(net34),
    .C(net16),
    .D(net17),
    .X(_06794_));
 sky130_fd_sc_hd__nand4_4 _17057_ (.A(net64),
    .B(net34),
    .C(net16),
    .D(net17),
    .Y(_06795_));
 sky130_fd_sc_hd__o211ai_2 _17058_ (.A1(_01934_),
    .A2(_02076_),
    .B1(_06793_),
    .C1(_06795_),
    .Y(_06797_));
 sky130_fd_sc_hd__o21bai_2 _17059_ (.A1(_06792_),
    .A2(_06794_),
    .B1_N(_06791_),
    .Y(_06798_));
 sky130_fd_sc_hd__a22o_1 _17060_ (.A1(net35),
    .A2(net15),
    .B1(_06793_),
    .B2(_06795_),
    .X(_06799_));
 sky130_fd_sc_hd__nand4_2 _17061_ (.A(_06793_),
    .B(_06795_),
    .C(net35),
    .D(net15),
    .Y(_06800_));
 sky130_fd_sc_hd__nand2_1 _17062_ (.A(_06799_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__nand3_4 _17063_ (.A(_06790_),
    .B(_06797_),
    .C(_06798_),
    .Y(_06802_));
 sky130_fd_sc_hd__nand3_4 _17064_ (.A(_06799_),
    .B(_06800_),
    .C(_06789_),
    .Y(_06803_));
 sky130_fd_sc_hd__nand2_1 _17065_ (.A(net38),
    .B(net11),
    .Y(_06804_));
 sky130_fd_sc_hd__nand2_1 _17066_ (.A(net36),
    .B(net14),
    .Y(_06805_));
 sky130_fd_sc_hd__a22oi_4 _17067_ (.A1(net37),
    .A2(net13),
    .B1(net14),
    .B2(net36),
    .Y(_06806_));
 sky130_fd_sc_hd__a22o_1 _17068_ (.A1(net37),
    .A2(net13),
    .B1(net14),
    .B2(net36),
    .X(_06808_));
 sky130_fd_sc_hd__and4_2 _17069_ (.A(net36),
    .B(net37),
    .C(net13),
    .D(net14),
    .X(_06809_));
 sky130_fd_sc_hd__nand4_2 _17070_ (.A(net36),
    .B(net37),
    .C(net13),
    .D(net14),
    .Y(_06810_));
 sky130_fd_sc_hd__and3_1 _17071_ (.A(_06804_),
    .B(_06808_),
    .C(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__a211o_1 _17072_ (.A1(net38),
    .A2(net11),
    .B1(_06806_),
    .C1(_06809_),
    .X(_06812_));
 sky130_fd_sc_hd__o211a_1 _17073_ (.A1(_06806_),
    .A2(_06809_),
    .B1(net38),
    .C1(net11),
    .X(_06813_));
 sky130_fd_sc_hd__a21o_1 _17074_ (.A1(_06808_),
    .A2(_06810_),
    .B1(_06804_),
    .X(_06814_));
 sky130_fd_sc_hd__o2bb2a_1 _17075_ (.A1_N(net38),
    .A2_N(net11),
    .B1(_06806_),
    .B2(_06809_),
    .X(_06815_));
 sky130_fd_sc_hd__and4_1 _17076_ (.A(_06808_),
    .B(_06810_),
    .C(net38),
    .D(net11),
    .X(_06816_));
 sky130_fd_sc_hd__o2bb2ai_1 _17077_ (.A1_N(_06802_),
    .A2_N(_06803_),
    .B1(_06811_),
    .B2(_06813_),
    .Y(_06817_));
 sky130_fd_sc_hd__o211ai_1 _17078_ (.A1(_06815_),
    .A2(_06816_),
    .B1(_06802_),
    .C1(_06803_),
    .Y(_06819_));
 sky130_fd_sc_hd__o2bb2ai_4 _17079_ (.A1_N(_06802_),
    .A2_N(_06803_),
    .B1(_06815_),
    .B2(_06816_),
    .Y(_06820_));
 sky130_fd_sc_hd__o211ai_4 _17080_ (.A1(_06811_),
    .A2(_06813_),
    .B1(_06802_),
    .C1(_06803_),
    .Y(_06821_));
 sky130_fd_sc_hd__o2bb2ai_4 _17081_ (.A1_N(_06383_),
    .A2_N(_06377_),
    .B1(_06373_),
    .B2(_06378_),
    .Y(_06822_));
 sky130_fd_sc_hd__a21boi_1 _17082_ (.A1(_06377_),
    .A2(_06383_),
    .B1_N(_06380_),
    .Y(_06823_));
 sky130_fd_sc_hd__a21oi_4 _17083_ (.A1(_06820_),
    .A2(_06821_),
    .B1(_06822_),
    .Y(_06824_));
 sky130_fd_sc_hd__nand3_2 _17084_ (.A(_06817_),
    .B(_06819_),
    .C(_06823_),
    .Y(_06825_));
 sky130_fd_sc_hd__nand3_4 _17085_ (.A(_06820_),
    .B(_06821_),
    .C(_06822_),
    .Y(_06826_));
 sky130_fd_sc_hd__nand2_2 _17086_ (.A(_06419_),
    .B(_06435_),
    .Y(_06827_));
 sky130_fd_sc_hd__a22oi_4 _17087_ (.A1(_06419_),
    .A2(_06435_),
    .B1(_06825_),
    .B2(_06826_),
    .Y(_06828_));
 sky130_fd_sc_hd__and3b_1 _17088_ (.A_N(_06827_),
    .B(_06826_),
    .C(_06825_),
    .X(_06830_));
 sky130_fd_sc_hd__a21oi_2 _17089_ (.A1(_06825_),
    .A2(_06826_),
    .B1(_06827_),
    .Y(_06831_));
 sky130_fd_sc_hd__and3_1 _17090_ (.A(_06825_),
    .B(_06826_),
    .C(_06827_),
    .X(_06832_));
 sky130_fd_sc_hd__nor2_1 _17091_ (.A(_06831_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__a21o_1 _17092_ (.A1(_06320_),
    .A2(_06325_),
    .B1(_06321_),
    .X(_06834_));
 sky130_fd_sc_hd__a21oi_1 _17093_ (.A1(_06320_),
    .A2(_06325_),
    .B1(_06321_),
    .Y(_06835_));
 sky130_fd_sc_hd__nand2_1 _17094_ (.A(net63),
    .B(net18),
    .Y(_06836_));
 sky130_fd_sc_hd__a22oi_4 _17095_ (.A1(net62),
    .A2(net19),
    .B1(net20),
    .B2(net61),
    .Y(_06837_));
 sky130_fd_sc_hd__a22o_1 _17096_ (.A1(net62),
    .A2(net19),
    .B1(net20),
    .B2(net61),
    .X(_06838_));
 sky130_fd_sc_hd__and4_2 _17097_ (.A(net61),
    .B(net62),
    .C(net19),
    .D(net20),
    .X(_06839_));
 sky130_fd_sc_hd__o221ai_4 _17098_ (.A1(_01890_),
    .A2(_02131_),
    .B1(_02163_),
    .B2(_06366_),
    .C1(_06838_),
    .Y(_06841_));
 sky130_fd_sc_hd__o21bai_1 _17099_ (.A1(_06837_),
    .A2(_06839_),
    .B1_N(_06836_),
    .Y(_06842_));
 sky130_fd_sc_hd__o22a_1 _17100_ (.A1(_01890_),
    .A2(_02131_),
    .B1(_06837_),
    .B2(_06839_),
    .X(_06843_));
 sky130_fd_sc_hd__o22ai_2 _17101_ (.A1(_01890_),
    .A2(_02131_),
    .B1(_06837_),
    .B2(_06839_),
    .Y(_06844_));
 sky130_fd_sc_hd__a41o_1 _17102_ (.A1(net61),
    .A2(net62),
    .A3(net19),
    .A4(net20),
    .B1(_06836_),
    .X(_06845_));
 sky130_fd_sc_hd__nand3_2 _17103_ (.A(_06842_),
    .B(_06834_),
    .C(_06841_),
    .Y(_06846_));
 sky130_fd_sc_hd__o21ai_1 _17104_ (.A1(_06837_),
    .A2(_06845_),
    .B1(_06835_),
    .Y(_06847_));
 sky130_fd_sc_hd__o211a_1 _17105_ (.A1(_06845_),
    .A2(_06837_),
    .B1(_06835_),
    .C1(_06844_),
    .X(_06848_));
 sky130_fd_sc_hd__o211ai_2 _17106_ (.A1(_06845_),
    .A2(_06837_),
    .B1(_06835_),
    .C1(_06844_),
    .Y(_06849_));
 sky130_fd_sc_hd__o2bb2a_1 _17107_ (.A1_N(net63),
    .A2_N(net17),
    .B1(_02131_),
    .B2(_06366_),
    .X(_06850_));
 sky130_fd_sc_hd__a21o_1 _17108_ (.A1(_06363_),
    .A2(_06369_),
    .B1(_06364_),
    .X(_06852_));
 sky130_fd_sc_hd__a21oi_1 _17109_ (.A1(_06363_),
    .A2(_06369_),
    .B1(_06364_),
    .Y(_06853_));
 sky130_fd_sc_hd__a21oi_2 _17110_ (.A1(_06846_),
    .A2(_06849_),
    .B1(_06852_),
    .Y(_06854_));
 sky130_fd_sc_hd__and3_1 _17111_ (.A(_06846_),
    .B(_06849_),
    .C(_06852_),
    .X(_06855_));
 sky130_fd_sc_hd__o2bb2ai_1 _17112_ (.A1_N(_06846_),
    .A2_N(_06849_),
    .B1(_06850_),
    .B2(_06364_),
    .Y(_06856_));
 sky130_fd_sc_hd__a31o_1 _17113_ (.A1(_06842_),
    .A2(_06834_),
    .A3(_06841_),
    .B1(_06852_),
    .X(_06857_));
 sky130_fd_sc_hd__o21ai_4 _17114_ (.A1(_06848_),
    .A2(_06857_),
    .B1(_06856_),
    .Y(_06858_));
 sky130_fd_sc_hd__nand2_1 _17115_ (.A(net60),
    .B(net21),
    .Y(_06859_));
 sky130_fd_sc_hd__nand4_4 _17116_ (.A(net58),
    .B(net59),
    .C(net22),
    .D(net24),
    .Y(_06860_));
 sky130_fd_sc_hd__a22oi_2 _17117_ (.A1(net59),
    .A2(net22),
    .B1(net24),
    .B2(net58),
    .Y(_06861_));
 sky130_fd_sc_hd__a22o_1 _17118_ (.A1(net59),
    .A2(net22),
    .B1(net24),
    .B2(net58),
    .X(_06863_));
 sky130_fd_sc_hd__a22oi_4 _17119_ (.A1(net60),
    .A2(net21),
    .B1(_06860_),
    .B2(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__o2bb2ai_1 _17120_ (.A1_N(_06860_),
    .A2_N(_06863_),
    .B1(_01835_),
    .B2(_02185_),
    .Y(_06865_));
 sky130_fd_sc_hd__and3_1 _17121_ (.A(_06860_),
    .B(net21),
    .C(net60),
    .X(_06866_));
 sky130_fd_sc_hd__a41o_1 _17122_ (.A1(net58),
    .A2(net59),
    .A3(net22),
    .A4(net24),
    .B1(_06859_),
    .X(_06867_));
 sky130_fd_sc_hd__and4_1 _17123_ (.A(_06863_),
    .B(net21),
    .C(net60),
    .D(_06860_),
    .X(_06868_));
 sky130_fd_sc_hd__o21ai_1 _17124_ (.A1(_06861_),
    .A2(_06867_),
    .B1(_06865_),
    .Y(_06869_));
 sky130_fd_sc_hd__a21oi_1 _17125_ (.A1(_06863_),
    .A2(_06866_),
    .B1(_06864_),
    .Y(_06870_));
 sky130_fd_sc_hd__a22o_1 _17126_ (.A1(_06011_),
    .A2(_06338_),
    .B1(_06341_),
    .B2(_06337_),
    .X(_06871_));
 sky130_fd_sc_hd__and2_1 _17127_ (.A(net55),
    .B(net25),
    .X(_06872_));
 sky130_fd_sc_hd__o211ai_1 _17128_ (.A1(_01780_),
    .A2(_02251_),
    .B1(_06341_),
    .C1(_06342_),
    .Y(_06874_));
 sky130_fd_sc_hd__nand2_1 _17129_ (.A(_06343_),
    .B(_06872_),
    .Y(_06875_));
 sky130_fd_sc_hd__o2bb2ai_1 _17130_ (.A1_N(_06341_),
    .A2_N(_06342_),
    .B1(_01780_),
    .B2(_02251_),
    .Y(_06876_));
 sky130_fd_sc_hd__nand4_1 _17131_ (.A(_06342_),
    .B(net25),
    .C(net55),
    .D(_06341_),
    .Y(_06877_));
 sky130_fd_sc_hd__a21boi_1 _17132_ (.A1(_06876_),
    .A2(_06877_),
    .B1_N(_06871_),
    .Y(_06878_));
 sky130_fd_sc_hd__nand3_1 _17133_ (.A(_06871_),
    .B(_06874_),
    .C(_06875_),
    .Y(_06879_));
 sky130_fd_sc_hd__and4_4 _17134_ (.A(net33),
    .B(net44),
    .C(net55),
    .D(net25),
    .X(_06880_));
 sky130_fd_sc_hd__nand4_4 _17135_ (.A(net33),
    .B(net44),
    .C(net55),
    .D(net25),
    .Y(_06881_));
 sky130_fd_sc_hd__nand3_2 _17136_ (.A(_06871_),
    .B(_06876_),
    .C(_06877_),
    .Y(_06882_));
 sky130_fd_sc_hd__a21oi_2 _17137_ (.A1(_06343_),
    .A2(_06872_),
    .B1(_06871_),
    .Y(_06883_));
 sky130_fd_sc_hd__a22o_1 _17138_ (.A1(_06341_),
    .A2(_06348_),
    .B1(_06343_),
    .B2(_06872_),
    .X(_06885_));
 sky130_fd_sc_hd__nand3_4 _17139_ (.A(_06870_),
    .B(_06879_),
    .C(_06881_),
    .Y(_06886_));
 sky130_fd_sc_hd__o21ai_2 _17140_ (.A1(_06864_),
    .A2(_06868_),
    .B1(_06882_),
    .Y(_06887_));
 sky130_fd_sc_hd__o211ai_4 _17141_ (.A1(_06864_),
    .A2(_06868_),
    .B1(_06882_),
    .C1(_06885_),
    .Y(_06888_));
 sky130_fd_sc_hd__a32oi_4 _17142_ (.A1(_06336_),
    .A2(_06344_),
    .A3(_06345_),
    .B1(_06351_),
    .B2(_06332_),
    .Y(_06889_));
 sky130_fd_sc_hd__a21oi_4 _17143_ (.A1(_06886_),
    .A2(_06888_),
    .B1(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__a21o_1 _17144_ (.A1(_06886_),
    .A2(_06888_),
    .B1(_06889_),
    .X(_06891_));
 sky130_fd_sc_hd__o211a_2 _17145_ (.A1(_06883_),
    .A2(_06887_),
    .B1(_06886_),
    .C1(_06889_),
    .X(_06892_));
 sky130_fd_sc_hd__o211ai_4 _17146_ (.A1(_06883_),
    .A2(_06887_),
    .B1(_06886_),
    .C1(_06889_),
    .Y(_06893_));
 sky130_fd_sc_hd__o22ai_4 _17147_ (.A1(_06854_),
    .A2(_06855_),
    .B1(_06890_),
    .B2(_06892_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand3_2 _17148_ (.A(_06891_),
    .B(_06893_),
    .C(_06858_),
    .Y(_06896_));
 sky130_fd_sc_hd__nor2_1 _17149_ (.A(_06858_),
    .B(_06890_),
    .Y(_06897_));
 sky130_fd_sc_hd__o21ai_1 _17150_ (.A1(_06854_),
    .A2(_06855_),
    .B1(_06893_),
    .Y(_06898_));
 sky130_fd_sc_hd__o21ai_1 _17151_ (.A1(_06890_),
    .A2(_06892_),
    .B1(_06858_),
    .Y(_06899_));
 sky130_fd_sc_hd__a22oi_4 _17152_ (.A1(_06362_),
    .A2(_06397_),
    .B1(_06894_),
    .B2(_06896_),
    .Y(_06900_));
 sky130_fd_sc_hd__o211ai_4 _17153_ (.A1(_06890_),
    .A2(_06898_),
    .B1(_06899_),
    .C1(_06398_),
    .Y(_06901_));
 sky130_fd_sc_hd__o2111a_1 _17154_ (.A1(_06392_),
    .A2(_06389_),
    .B1(_06362_),
    .C1(_06896_),
    .D1(_06894_),
    .X(_06902_));
 sky130_fd_sc_hd__o2111ai_4 _17155_ (.A1(_06392_),
    .A2(_06389_),
    .B1(_06362_),
    .C1(_06896_),
    .D1(_06894_),
    .Y(_06903_));
 sky130_fd_sc_hd__o22ai_4 _17156_ (.A1(_06831_),
    .A2(_06832_),
    .B1(_06900_),
    .B2(_06902_),
    .Y(_06904_));
 sky130_fd_sc_hd__o21a_1 _17157_ (.A1(_06828_),
    .A2(_06830_),
    .B1(_06903_),
    .X(_06905_));
 sky130_fd_sc_hd__o21ai_2 _17158_ (.A1(_06828_),
    .A2(_06830_),
    .B1(_06903_),
    .Y(_06907_));
 sky130_fd_sc_hd__and3_1 _17159_ (.A(_06833_),
    .B(_06901_),
    .C(_06903_),
    .X(_06908_));
 sky130_fd_sc_hd__o211ai_4 _17160_ (.A1(_06828_),
    .A2(_06830_),
    .B1(_06901_),
    .C1(_06903_),
    .Y(_06909_));
 sky130_fd_sc_hd__a21oi_2 _17161_ (.A1(_06833_),
    .A2(_06903_),
    .B1(_06900_),
    .Y(_06910_));
 sky130_fd_sc_hd__o31a_1 _17162_ (.A1(_06402_),
    .A2(_06316_),
    .A3(_06400_),
    .B1(_06451_),
    .X(_06911_));
 sky130_fd_sc_hd__a32oi_4 _17163_ (.A1(_06316_),
    .A2(_06391_),
    .A3(_06399_),
    .B1(_06405_),
    .B2(_06451_),
    .Y(_06912_));
 sky130_fd_sc_hd__a21oi_4 _17164_ (.A1(_06904_),
    .A2(_06909_),
    .B1(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__o2bb2ai_2 _17165_ (.A1_N(_06904_),
    .A2_N(_06909_),
    .B1(_06911_),
    .B2(_06406_),
    .Y(_06914_));
 sky130_fd_sc_hd__nand2_1 _17166_ (.A(_06912_),
    .B(_06904_),
    .Y(_06915_));
 sky130_fd_sc_hd__o211a_2 _17167_ (.A1(_06900_),
    .A2(_06907_),
    .B1(_06904_),
    .C1(_06912_),
    .X(_06916_));
 sky130_fd_sc_hd__o211ai_2 _17168_ (.A1(_06900_),
    .A2(_06907_),
    .B1(_06904_),
    .C1(_06912_),
    .Y(_06918_));
 sky130_fd_sc_hd__o21ai_2 _17169_ (.A1(_06786_),
    .A2(_06787_),
    .B1(_06914_),
    .Y(_06919_));
 sky130_fd_sc_hd__o211a_2 _17170_ (.A1(_06786_),
    .A2(_06787_),
    .B1(_06914_),
    .C1(_06918_),
    .X(_06920_));
 sky130_fd_sc_hd__o2bb2ai_2 _17171_ (.A1_N(_06783_),
    .A2_N(_06784_),
    .B1(_06913_),
    .B2(_06916_),
    .Y(_06921_));
 sky130_fd_sc_hd__o211ai_2 _17172_ (.A1(_06908_),
    .A2(_06915_),
    .B1(_06914_),
    .C1(_06788_),
    .Y(_06922_));
 sky130_fd_sc_hd__o22ai_2 _17173_ (.A1(_06786_),
    .A2(_06787_),
    .B1(_06913_),
    .B2(_06916_),
    .Y(_06923_));
 sky130_fd_sc_hd__nand2_2 _17174_ (.A(_06710_),
    .B(_06921_),
    .Y(_06924_));
 sky130_fd_sc_hd__o211a_1 _17175_ (.A1(_06916_),
    .A2(_06919_),
    .B1(_06921_),
    .C1(_06710_),
    .X(_06925_));
 sky130_fd_sc_hd__o211ai_4 _17176_ (.A1(_06916_),
    .A2(_06919_),
    .B1(_06921_),
    .C1(_06710_),
    .Y(_06926_));
 sky130_fd_sc_hd__o2111a_1 _17177_ (.A1(_06550_),
    .A2(_06457_),
    .B1(_06459_),
    .C1(_06922_),
    .D1(_06923_),
    .X(_06927_));
 sky130_fd_sc_hd__o2111ai_4 _17178_ (.A1(_06550_),
    .A2(_06457_),
    .B1(_06459_),
    .C1(_06922_),
    .D1(_06923_),
    .Y(_06929_));
 sky130_fd_sc_hd__o211ai_4 _17179_ (.A1(_06920_),
    .A2(_06924_),
    .B1(_06929_),
    .C1(_06709_),
    .Y(_06930_));
 sky130_fd_sc_hd__a21o_1 _17180_ (.A1(_06926_),
    .A2(_06929_),
    .B1(_06709_),
    .X(_06931_));
 sky130_fd_sc_hd__o211ai_4 _17181_ (.A1(_06705_),
    .A2(_06701_),
    .B1(_06704_),
    .C1(_06929_),
    .Y(_06932_));
 sky130_fd_sc_hd__a22o_1 _17182_ (.A1(_06704_),
    .A2(_06707_),
    .B1(_06926_),
    .B2(_06929_),
    .X(_06933_));
 sky130_fd_sc_hd__o211a_1 _17183_ (.A1(_06925_),
    .A2(_06932_),
    .B1(_06933_),
    .C1(_06605_),
    .X(_06934_));
 sky130_fd_sc_hd__o211ai_2 _17184_ (.A1(_06925_),
    .A2(_06932_),
    .B1(_06933_),
    .C1(_06605_),
    .Y(_06935_));
 sky130_fd_sc_hd__o211ai_4 _17185_ (.A1(_06558_),
    .A2(_06604_),
    .B1(_06930_),
    .C1(_06931_),
    .Y(_06936_));
 sky130_fd_sc_hd__a22o_1 _17186_ (.A1(_06307_),
    .A2(_06311_),
    .B1(_06935_),
    .B2(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__nand4_2 _17187_ (.A(_06307_),
    .B(_06311_),
    .C(_06935_),
    .D(_06936_),
    .Y(_06938_));
 sky130_fd_sc_hd__a21o_1 _17188_ (.A1(_06935_),
    .A2(_06936_),
    .B1(_06603_),
    .X(_06940_));
 sky130_fd_sc_hd__a31oi_4 _17189_ (.A1(_06606_),
    .A2(_06930_),
    .A3(_06931_),
    .B1(_06602_),
    .Y(_06941_));
 sky130_fd_sc_hd__nand3_1 _17190_ (.A(_06603_),
    .B(_06935_),
    .C(_06936_),
    .Y(_06942_));
 sky130_fd_sc_hd__a32oi_4 _17191_ (.A1(_06222_),
    .A2(_06561_),
    .A3(_06562_),
    .B1(_06567_),
    .B2(_06572_),
    .Y(_06943_));
 sky130_fd_sc_hd__a21oi_2 _17192_ (.A1(_06569_),
    .A2(_06571_),
    .B1(_06565_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand3_4 _17193_ (.A(_06937_),
    .B(_06938_),
    .C(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__and3_1 _17194_ (.A(_06940_),
    .B(_06943_),
    .C(_06942_),
    .X(_06946_));
 sky130_fd_sc_hd__nand3_2 _17195_ (.A(_06940_),
    .B(_06942_),
    .C(_06943_),
    .Y(_06947_));
 sky130_fd_sc_hd__o311a_1 _17196_ (.A1(_01802_),
    .A2(_02229_),
    .A3(_05519_),
    .B1(_05888_),
    .C1(_06293_),
    .X(_06948_));
 sky130_fd_sc_hd__o21a_1 _17197_ (.A1(_06266_),
    .A2(_06290_),
    .B1(_06293_),
    .X(_06949_));
 sky130_fd_sc_hd__o2bb2ai_1 _17198_ (.A1_N(_06945_),
    .A2_N(_06947_),
    .B1(_06948_),
    .B2(_06290_),
    .Y(_06951_));
 sky130_fd_sc_hd__a31oi_1 _17199_ (.A1(_06937_),
    .A2(_06938_),
    .A3(_06944_),
    .B1(_06949_),
    .Y(_06952_));
 sky130_fd_sc_hd__nand3b_1 _17200_ (.A_N(_06949_),
    .B(_06947_),
    .C(_06945_),
    .Y(_06953_));
 sky130_fd_sc_hd__a21o_1 _17201_ (.A1(_06945_),
    .A2(_06947_),
    .B1(_06949_),
    .X(_06954_));
 sky130_fd_sc_hd__o2111ai_4 _17202_ (.A1(_06266_),
    .A2(_06290_),
    .B1(_06293_),
    .C1(_06945_),
    .D1(_06947_),
    .Y(_06955_));
 sky130_fd_sc_hd__a31o_1 _17203_ (.A1(_06220_),
    .A2(_06575_),
    .A3(_06576_),
    .B1(_05909_),
    .X(_06956_));
 sky130_fd_sc_hd__a21boi_2 _17204_ (.A1(_05909_),
    .A2(_06578_),
    .B1_N(_06580_),
    .Y(_06957_));
 sky130_fd_sc_hd__nand3_1 _17205_ (.A(_06954_),
    .B(_06955_),
    .C(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__nand4_4 _17206_ (.A(_06578_),
    .B(_06951_),
    .C(_06953_),
    .D(_06956_),
    .Y(_06959_));
 sky130_fd_sc_hd__nand2_1 _17207_ (.A(_06958_),
    .B(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__a21bo_1 _17208_ (.A1(_06585_),
    .A2(_06601_),
    .B1_N(_06586_),
    .X(_06962_));
 sky130_fd_sc_hd__xnor2_1 _17209_ (.A(_06960_),
    .B(_06962_),
    .Y(net91));
 sky130_fd_sc_hd__o21ai_1 _17210_ (.A1(_06290_),
    .A2(_06948_),
    .B1(_06947_),
    .Y(_06963_));
 sky130_fd_sc_hd__a21oi_1 _17211_ (.A1(_06603_),
    .A2(_06936_),
    .B1(_06934_),
    .Y(_06964_));
 sky130_fd_sc_hd__a21oi_2 _17212_ (.A1(_06700_),
    .A2(_06703_),
    .B1(_06701_),
    .Y(_06965_));
 sky130_fd_sc_hd__a31o_1 _17213_ (.A1(_06694_),
    .A2(_06696_),
    .A3(_06699_),
    .B1(_06706_),
    .X(_06966_));
 sky130_fd_sc_hd__a31oi_2 _17214_ (.A1(_06704_),
    .A2(_06707_),
    .A3(_06929_),
    .B1(_06925_),
    .Y(_06967_));
 sky130_fd_sc_hd__o22ai_4 _17215_ (.A1(_06920_),
    .A2(_06924_),
    .B1(_06709_),
    .B2(_06927_),
    .Y(_06968_));
 sky130_fd_sc_hd__a21oi_2 _17216_ (.A1(_06641_),
    .A2(_06644_),
    .B1(_06688_),
    .Y(_06969_));
 sky130_fd_sc_hd__o31a_2 _17217_ (.A1(_06640_),
    .A2(_06643_),
    .A3(_06690_),
    .B1(_06689_),
    .X(_06970_));
 sky130_fd_sc_hd__a31oi_4 _17218_ (.A1(_06769_),
    .A2(_06770_),
    .A3(_06775_),
    .B1(_06781_),
    .Y(_06972_));
 sky130_fd_sc_hd__a32oi_4 _17219_ (.A1(_06771_),
    .A2(_06772_),
    .A3(_06773_),
    .B1(_06779_),
    .B2(_06780_),
    .Y(_06973_));
 sky130_fd_sc_hd__a31o_1 _17220_ (.A1(_06771_),
    .A2(_06772_),
    .A3(_06773_),
    .B1(_06972_),
    .X(_06974_));
 sky130_fd_sc_hd__o22ai_4 _17221_ (.A1(_06619_),
    .A2(_06624_),
    .B1(_06632_),
    .B2(_06622_),
    .Y(_06975_));
 sky130_fd_sc_hd__a22o_1 _17222_ (.A1(net27),
    .A2(net56),
    .B1(_01791_),
    .B2(net57),
    .X(_06976_));
 sky130_fd_sc_hd__nand3_2 _17223_ (.A(_01791_),
    .B(net56),
    .C(net27),
    .Y(_06977_));
 sky130_fd_sc_hd__and4_1 _17224_ (.A(_01791_),
    .B(net56),
    .C(net57),
    .D(net27),
    .X(_06978_));
 sky130_fd_sc_hd__or2_1 _17225_ (.A(_02240_),
    .B(_06977_),
    .X(_06979_));
 sky130_fd_sc_hd__o21ai_2 _17226_ (.A1(_02240_),
    .A2(_06977_),
    .B1(_06976_),
    .Y(_06980_));
 sky130_fd_sc_hd__o21ai_1 _17227_ (.A1(_06272_),
    .A2(_06612_),
    .B1(_06611_),
    .Y(_06981_));
 sky130_fd_sc_hd__a21oi_2 _17228_ (.A1(_06272_),
    .A2(_06612_),
    .B1(_06611_),
    .Y(_06983_));
 sky130_fd_sc_hd__o31a_1 _17229_ (.A1(_01769_),
    .A2(_02207_),
    .A3(_06615_),
    .B1(_06614_),
    .X(_06984_));
 sky130_fd_sc_hd__nand2_1 _17230_ (.A(net28),
    .B(net54),
    .Y(_06985_));
 sky130_fd_sc_hd__nand2_2 _17231_ (.A(net30),
    .B(net53),
    .Y(_06986_));
 sky130_fd_sc_hd__nand2_1 _17232_ (.A(net30),
    .B(net52),
    .Y(_06987_));
 sky130_fd_sc_hd__and4_1 _17233_ (.A(net29),
    .B(net30),
    .C(net52),
    .D(net53),
    .X(_06988_));
 sky130_fd_sc_hd__a22oi_4 _17234_ (.A1(net30),
    .A2(net52),
    .B1(net53),
    .B2(net29),
    .Y(_06989_));
 sky130_fd_sc_hd__a22o_1 _17235_ (.A1(net30),
    .A2(net52),
    .B1(net53),
    .B2(net29),
    .X(_06990_));
 sky130_fd_sc_hd__o21ai_1 _17236_ (.A1(_06612_),
    .A2(_06986_),
    .B1(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__o221ai_1 _17237_ (.A1(_01748_),
    .A2(_02207_),
    .B1(_06612_),
    .B2(_06986_),
    .C1(_06990_),
    .Y(_06992_));
 sky130_fd_sc_hd__nand3_1 _17238_ (.A(_06991_),
    .B(net54),
    .C(net28),
    .Y(_06994_));
 sky130_fd_sc_hd__o22ai_4 _17239_ (.A1(_01748_),
    .A2(_02207_),
    .B1(_06988_),
    .B2(_06989_),
    .Y(_06995_));
 sky130_fd_sc_hd__o2111ai_4 _17240_ (.A1(_06612_),
    .A2(_06986_),
    .B1(net28),
    .C1(net54),
    .D1(_06990_),
    .Y(_06996_));
 sky130_fd_sc_hd__a22oi_4 _17241_ (.A1(_06616_),
    .A2(_06981_),
    .B1(_06995_),
    .B2(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__nand3_1 _17242_ (.A(_06984_),
    .B(_06992_),
    .C(_06994_),
    .Y(_06998_));
 sky130_fd_sc_hd__a2bb2oi_1 _17243_ (.A1_N(_06613_),
    .A2_N(_06983_),
    .B1(_06985_),
    .B2(_06991_),
    .Y(_06999_));
 sky130_fd_sc_hd__o211ai_4 _17244_ (.A1(_06613_),
    .A2(_06983_),
    .B1(_06995_),
    .C1(_06996_),
    .Y(_07000_));
 sky130_fd_sc_hd__a22oi_2 _17245_ (.A1(_06976_),
    .A2(_06979_),
    .B1(_06998_),
    .B2(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__a22o_1 _17246_ (.A1(_06976_),
    .A2(_06979_),
    .B1(_06998_),
    .B2(_07000_),
    .X(_07002_));
 sky130_fd_sc_hd__a211oi_2 _17247_ (.A1(_06999_),
    .A2(_06996_),
    .B1(_06980_),
    .C1(_06997_),
    .Y(_07003_));
 sky130_fd_sc_hd__a211o_1 _17248_ (.A1(_06999_),
    .A2(_06996_),
    .B1(_06980_),
    .C1(_06997_),
    .X(_07005_));
 sky130_fd_sc_hd__o21bai_4 _17249_ (.A1(_07001_),
    .A2(_07003_),
    .B1_N(_06975_),
    .Y(_07006_));
 sky130_fd_sc_hd__inv_2 _17250_ (.A(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__nand3_4 _17251_ (.A(_06975_),
    .B(_07002_),
    .C(_07005_),
    .Y(_07008_));
 sky130_fd_sc_hd__o31a_1 _17252_ (.A1(net23),
    .A2(_02240_),
    .A3(_06626_),
    .B1(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__o311a_1 _17253_ (.A1(net23),
    .A2(_02240_),
    .A3(_06626_),
    .B1(_07006_),
    .C1(_07008_),
    .X(_07010_));
 sky130_fd_sc_hd__nand3_1 _17254_ (.A(_06628_),
    .B(_07006_),
    .C(_07008_),
    .Y(_07011_));
 sky130_fd_sc_hd__a21oi_2 _17255_ (.A1(_07006_),
    .A2(_07008_),
    .B1(_06628_),
    .Y(_07012_));
 sky130_fd_sc_hd__a21o_1 _17256_ (.A1(_07006_),
    .A2(_07008_),
    .B1(_06628_),
    .X(_07013_));
 sky130_fd_sc_hd__a21oi_2 _17257_ (.A1(_07006_),
    .A2(_07008_),
    .B1(_06627_),
    .Y(_07014_));
 sky130_fd_sc_hd__and3_1 _17258_ (.A(_07006_),
    .B(_07008_),
    .C(_06627_),
    .X(_07016_));
 sky130_fd_sc_hd__o2bb2ai_2 _17259_ (.A1_N(_06648_),
    .A2_N(_06682_),
    .B1(_06678_),
    .B2(_06672_),
    .Y(_07017_));
 sky130_fd_sc_hd__a21oi_4 _17260_ (.A1(_06648_),
    .A2(_06682_),
    .B1(_06679_),
    .Y(_07018_));
 sky130_fd_sc_hd__o311a_2 _17261_ (.A1(_01857_),
    .A2(_02152_),
    .A3(_06237_),
    .B1(_06240_),
    .C1(_06667_),
    .X(_07019_));
 sky130_fd_sc_hd__a21oi_4 _17262_ (.A1(_06669_),
    .A2(_06652_),
    .B1(_06666_),
    .Y(_07020_));
 sky130_fd_sc_hd__a21boi_4 _17263_ (.A1(_06747_),
    .A2(_06760_),
    .B1_N(_06748_),
    .Y(_07021_));
 sky130_fd_sc_hd__a21bo_1 _17264_ (.A1(_06747_),
    .A2(_06760_),
    .B1_N(_06748_),
    .X(_07022_));
 sky130_fd_sc_hd__o21a_1 _17265_ (.A1(_01868_),
    .A2(_02152_),
    .B1(_06660_),
    .X(_07023_));
 sky130_fd_sc_hd__and3_1 _17266_ (.A(_06658_),
    .B(net51),
    .C(net30),
    .X(_07024_));
 sky130_fd_sc_hd__a21oi_2 _17267_ (.A1(_06484_),
    .A2(_06750_),
    .B1(_06749_),
    .Y(_07025_));
 sky130_fd_sc_hd__o21ai_2 _17268_ (.A1(_06749_),
    .A2(_06754_),
    .B1(_06753_),
    .Y(_07027_));
 sky130_fd_sc_hd__nand2_1 _17269_ (.A(net31),
    .B(net51),
    .Y(_07028_));
 sky130_fd_sc_hd__a22oi_4 _17270_ (.A1(net2),
    .A2(net49),
    .B1(net50),
    .B2(net32),
    .Y(_07029_));
 sky130_fd_sc_hd__a22o_2 _17271_ (.A1(net2),
    .A2(net49),
    .B1(net50),
    .B2(net32),
    .X(_07030_));
 sky130_fd_sc_hd__and4_2 _17272_ (.A(net2),
    .B(net32),
    .C(net49),
    .D(net50),
    .X(_07031_));
 sky130_fd_sc_hd__nand4_4 _17273_ (.A(net2),
    .B(net32),
    .C(net49),
    .D(net50),
    .Y(_07032_));
 sky130_fd_sc_hd__o211ai_1 _17274_ (.A1(_01879_),
    .A2(_02152_),
    .B1(_07030_),
    .C1(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__a21o_1 _17275_ (.A1(_07030_),
    .A2(_07032_),
    .B1(_07028_),
    .X(_07034_));
 sky130_fd_sc_hd__nand4_4 _17276_ (.A(_07030_),
    .B(_07032_),
    .C(net31),
    .D(net51),
    .Y(_07035_));
 sky130_fd_sc_hd__o22ai_4 _17277_ (.A1(_01879_),
    .A2(_02152_),
    .B1(_07029_),
    .B2(_07031_),
    .Y(_07036_));
 sky130_fd_sc_hd__o211a_1 _17278_ (.A1(_06751_),
    .A2(_07025_),
    .B1(_07035_),
    .C1(_07036_),
    .X(_07038_));
 sky130_fd_sc_hd__o211ai_4 _17279_ (.A1(_06751_),
    .A2(_07025_),
    .B1(_07035_),
    .C1(_07036_),
    .Y(_07039_));
 sky130_fd_sc_hd__a21oi_4 _17280_ (.A1(_07035_),
    .A2(_07036_),
    .B1(_07027_),
    .Y(_07040_));
 sky130_fd_sc_hd__nand3b_2 _17281_ (.A_N(_07027_),
    .B(_07033_),
    .C(_07034_),
    .Y(_07041_));
 sky130_fd_sc_hd__o211ai_2 _17282_ (.A1(_06659_),
    .A2(_07024_),
    .B1(_07039_),
    .C1(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__o22ai_2 _17283_ (.A1(_06657_),
    .A2(_07023_),
    .B1(_07038_),
    .B2(_07040_),
    .Y(_07043_));
 sky130_fd_sc_hd__o22ai_4 _17284_ (.A1(_06659_),
    .A2(_07024_),
    .B1(_07038_),
    .B2(_07040_),
    .Y(_07044_));
 sky130_fd_sc_hd__o2111ai_4 _17285_ (.A1(_06656_),
    .A2(_06657_),
    .B1(_06660_),
    .C1(_07039_),
    .D1(_07041_),
    .Y(_07045_));
 sky130_fd_sc_hd__a21oi_4 _17286_ (.A1(_07044_),
    .A2(_07045_),
    .B1(_07021_),
    .Y(_07046_));
 sky130_fd_sc_hd__nand3_2 _17287_ (.A(_07022_),
    .B(_07042_),
    .C(_07043_),
    .Y(_07047_));
 sky130_fd_sc_hd__a21oi_2 _17288_ (.A1(_07042_),
    .A2(_07043_),
    .B1(_07022_),
    .Y(_07049_));
 sky130_fd_sc_hd__nand3_1 _17289_ (.A(_07021_),
    .B(_07044_),
    .C(_07045_),
    .Y(_07050_));
 sky130_fd_sc_hd__a31oi_4 _17290_ (.A1(_07021_),
    .A2(_07044_),
    .A3(_07045_),
    .B1(_07020_),
    .Y(_07051_));
 sky130_fd_sc_hd__nand2_1 _17291_ (.A(_07051_),
    .B(_07047_),
    .Y(_07052_));
 sky130_fd_sc_hd__o22ai_4 _17292_ (.A1(_06668_),
    .A2(_07019_),
    .B1(_07046_),
    .B2(_07049_),
    .Y(_07053_));
 sky130_fd_sc_hd__o22ai_4 _17293_ (.A1(_06666_),
    .A2(_06671_),
    .B1(_07046_),
    .B2(_07049_),
    .Y(_07054_));
 sky130_fd_sc_hd__o211ai_4 _17294_ (.A1(_06668_),
    .A2(_07019_),
    .B1(_07047_),
    .C1(_07050_),
    .Y(_07055_));
 sky130_fd_sc_hd__a21oi_4 _17295_ (.A1(_07054_),
    .A2(_07055_),
    .B1(_07018_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand3_4 _17296_ (.A(_07053_),
    .B(_07017_),
    .C(_07052_),
    .Y(_07057_));
 sky130_fd_sc_hd__a21oi_1 _17297_ (.A1(_07052_),
    .A2(_07053_),
    .B1(_07017_),
    .Y(_07058_));
 sky130_fd_sc_hd__nand3_2 _17298_ (.A(_07018_),
    .B(_07054_),
    .C(_07055_),
    .Y(_07060_));
 sky130_fd_sc_hd__a32oi_2 _17299_ (.A1(_07018_),
    .A2(_07054_),
    .A3(_07055_),
    .B1(_07013_),
    .B2(_07011_),
    .Y(_07061_));
 sky130_fd_sc_hd__o21ai_4 _17300_ (.A1(_07010_),
    .A2(_07012_),
    .B1(_07060_),
    .Y(_07062_));
 sky130_fd_sc_hd__o211a_1 _17301_ (.A1(_07010_),
    .A2(_07012_),
    .B1(_07057_),
    .C1(_07060_),
    .X(_07063_));
 sky130_fd_sc_hd__a2bb2oi_2 _17302_ (.A1_N(_07014_),
    .A2_N(_07016_),
    .B1(_07057_),
    .B2(_07060_),
    .Y(_07064_));
 sky130_fd_sc_hd__o22ai_4 _17303_ (.A1(_07014_),
    .A2(_07016_),
    .B1(_07056_),
    .B2(_07058_),
    .Y(_07065_));
 sky130_fd_sc_hd__o21ai_1 _17304_ (.A1(_07056_),
    .A2(_07062_),
    .B1(_07065_),
    .Y(_07066_));
 sky130_fd_sc_hd__o211a_2 _17305_ (.A1(_07056_),
    .A2(_07062_),
    .B1(_06973_),
    .C1(_07065_),
    .X(_07067_));
 sky130_fd_sc_hd__o211ai_4 _17306_ (.A1(_07056_),
    .A2(_07062_),
    .B1(_06973_),
    .C1(_07065_),
    .Y(_07068_));
 sky130_fd_sc_hd__o22a_2 _17307_ (.A1(_06776_),
    .A2(_06972_),
    .B1(_07063_),
    .B2(_07064_),
    .X(_07069_));
 sky130_fd_sc_hd__o22ai_4 _17308_ (.A1(_06776_),
    .A2(_06972_),
    .B1(_07063_),
    .B2(_07064_),
    .Y(_07071_));
 sky130_fd_sc_hd__a2bb2oi_2 _17309_ (.A1_N(_06690_),
    .A2_N(_06969_),
    .B1(_07068_),
    .B2(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__o22ai_1 _17310_ (.A1(_06690_),
    .A2(_06969_),
    .B1(_07067_),
    .B2(_07069_),
    .Y(_07073_));
 sky130_fd_sc_hd__a2bb2oi_2 _17311_ (.A1_N(_06688_),
    .A2_N(_06695_),
    .B1(_06974_),
    .B2(_07066_),
    .Y(_07074_));
 sky130_fd_sc_hd__o21ai_1 _17312_ (.A1(_06688_),
    .A2(_06695_),
    .B1(_07071_),
    .Y(_07075_));
 sky130_fd_sc_hd__o211a_1 _17313_ (.A1(_06688_),
    .A2(_06695_),
    .B1(_07068_),
    .C1(_07071_),
    .X(_07076_));
 sky130_fd_sc_hd__o211a_1 _17314_ (.A1(_06690_),
    .A2(_06969_),
    .B1(_07068_),
    .C1(_07071_),
    .X(_07077_));
 sky130_fd_sc_hd__a21oi_2 _17315_ (.A1(_07068_),
    .A2(_07071_),
    .B1(_06970_),
    .Y(_07078_));
 sky130_fd_sc_hd__a21oi_1 _17316_ (.A1(_07074_),
    .A2(_07068_),
    .B1(_07072_),
    .Y(_07079_));
 sky130_fd_sc_hd__o21ai_2 _17317_ (.A1(_07067_),
    .A2(_07075_),
    .B1(_07073_),
    .Y(_07080_));
 sky130_fd_sc_hd__o21ai_2 _17318_ (.A1(_06791_),
    .A2(_06792_),
    .B1(_06795_),
    .Y(_07082_));
 sky130_fd_sc_hd__o21a_1 _17319_ (.A1(_06791_),
    .A2(_06792_),
    .B1(_06795_),
    .X(_07083_));
 sky130_fd_sc_hd__nand2_1 _17320_ (.A(net35),
    .B(net16),
    .Y(_07084_));
 sky130_fd_sc_hd__a22oi_4 _17321_ (.A1(net34),
    .A2(net17),
    .B1(net18),
    .B2(net64),
    .Y(_07085_));
 sky130_fd_sc_hd__a22o_1 _17322_ (.A1(net34),
    .A2(net17),
    .B1(net18),
    .B2(net64),
    .X(_07086_));
 sky130_fd_sc_hd__and4_1 _17323_ (.A(net64),
    .B(net34),
    .C(net17),
    .D(net18),
    .X(_07087_));
 sky130_fd_sc_hd__nand4_2 _17324_ (.A(net64),
    .B(net34),
    .C(net17),
    .D(net18),
    .Y(_07088_));
 sky130_fd_sc_hd__o211ai_1 _17325_ (.A1(_01934_),
    .A2(_02098_),
    .B1(_07086_),
    .C1(_07088_),
    .Y(_07089_));
 sky130_fd_sc_hd__o21bai_1 _17326_ (.A1(_07085_),
    .A2(_07087_),
    .B1_N(_07084_),
    .Y(_07090_));
 sky130_fd_sc_hd__a22o_1 _17327_ (.A1(net35),
    .A2(net16),
    .B1(_07086_),
    .B2(_07088_),
    .X(_07091_));
 sky130_fd_sc_hd__a41o_1 _17328_ (.A1(net64),
    .A2(net34),
    .A3(net17),
    .A4(net18),
    .B1(_07084_),
    .X(_07093_));
 sky130_fd_sc_hd__nand3_2 _17329_ (.A(_07083_),
    .B(_07089_),
    .C(_07090_),
    .Y(_07094_));
 sky130_fd_sc_hd__o211ai_4 _17330_ (.A1(_07085_),
    .A2(_07093_),
    .B1(_07082_),
    .C1(_07091_),
    .Y(_07095_));
 sky130_fd_sc_hd__nand2_1 _17331_ (.A(net38),
    .B(net13),
    .Y(_07096_));
 sky130_fd_sc_hd__a22oi_2 _17332_ (.A1(net37),
    .A2(net14),
    .B1(net15),
    .B2(net36),
    .Y(_07097_));
 sky130_fd_sc_hd__a22o_1 _17333_ (.A1(net37),
    .A2(net14),
    .B1(net15),
    .B2(net36),
    .X(_07098_));
 sky130_fd_sc_hd__nand2_1 _17334_ (.A(net37),
    .B(net15),
    .Y(_07099_));
 sky130_fd_sc_hd__and4_1 _17335_ (.A(net36),
    .B(net37),
    .C(net14),
    .D(net15),
    .X(_07100_));
 sky130_fd_sc_hd__nand4_1 _17336_ (.A(net36),
    .B(net37),
    .C(net14),
    .D(net15),
    .Y(_07101_));
 sky130_fd_sc_hd__and3_1 _17337_ (.A(_07096_),
    .B(_07098_),
    .C(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__o211a_1 _17338_ (.A1(_07097_),
    .A2(_07100_),
    .B1(net38),
    .C1(net13),
    .X(_07104_));
 sky130_fd_sc_hd__o2bb2a_1 _17339_ (.A1_N(net38),
    .A2_N(net13),
    .B1(_07097_),
    .B2(_07100_),
    .X(_07105_));
 sky130_fd_sc_hd__and4_1 _17340_ (.A(_07098_),
    .B(_07101_),
    .C(net38),
    .D(net13),
    .X(_07106_));
 sky130_fd_sc_hd__nor2_1 _17341_ (.A(_07105_),
    .B(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__o2bb2ai_1 _17342_ (.A1_N(_07094_),
    .A2_N(_07095_),
    .B1(_07102_),
    .B2(_07104_),
    .Y(_07108_));
 sky130_fd_sc_hd__o211ai_1 _17343_ (.A1(_07105_),
    .A2(_07106_),
    .B1(_07094_),
    .C1(_07095_),
    .Y(_07109_));
 sky130_fd_sc_hd__o2bb2ai_2 _17344_ (.A1_N(_07094_),
    .A2_N(_07095_),
    .B1(_07105_),
    .B2(_07106_),
    .Y(_07110_));
 sky130_fd_sc_hd__o211ai_2 _17345_ (.A1(_07102_),
    .A2(_07104_),
    .B1(_07094_),
    .C1(_07095_),
    .Y(_07111_));
 sky130_fd_sc_hd__o2bb2ai_2 _17346_ (.A1_N(_06846_),
    .A2_N(_06853_),
    .B1(_06847_),
    .B2(_06843_),
    .Y(_07112_));
 sky130_fd_sc_hd__a21oi_1 _17347_ (.A1(_06846_),
    .A2(_06853_),
    .B1(_06848_),
    .Y(_07113_));
 sky130_fd_sc_hd__a21oi_1 _17348_ (.A1(_07110_),
    .A2(_07111_),
    .B1(_07112_),
    .Y(_07115_));
 sky130_fd_sc_hd__nand3_1 _17349_ (.A(_07108_),
    .B(_07109_),
    .C(_07113_),
    .Y(_07116_));
 sky130_fd_sc_hd__nand3_4 _17350_ (.A(_07110_),
    .B(_07111_),
    .C(_07112_),
    .Y(_07117_));
 sky130_fd_sc_hd__a32o_1 _17351_ (.A1(_06790_),
    .A2(_06797_),
    .A3(_06798_),
    .B1(_06812_),
    .B2(_06814_),
    .X(_07118_));
 sky130_fd_sc_hd__o21ai_1 _17352_ (.A1(_06790_),
    .A2(_06801_),
    .B1(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__a21boi_2 _17353_ (.A1(_07116_),
    .A2(_07117_),
    .B1_N(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__o2111a_1 _17354_ (.A1(_06801_),
    .A2(_06790_),
    .B1(_07117_),
    .C1(_07116_),
    .D1(_07118_),
    .X(_07121_));
 sky130_fd_sc_hd__a21oi_1 _17355_ (.A1(_07116_),
    .A2(_07117_),
    .B1(_07119_),
    .Y(_07122_));
 sky130_fd_sc_hd__a32o_1 _17356_ (.A1(_07108_),
    .A2(_07109_),
    .A3(_07113_),
    .B1(_07118_),
    .B2(_06803_),
    .X(_07123_));
 sky130_fd_sc_hd__and3_1 _17357_ (.A(_07116_),
    .B(_07117_),
    .C(_07119_),
    .X(_07124_));
 sky130_fd_sc_hd__o21ai_2 _17358_ (.A1(_06858_),
    .A2(_06890_),
    .B1(_06893_),
    .Y(_07126_));
 sky130_fd_sc_hd__o31ai_4 _17359_ (.A1(net33),
    .A2(net44),
    .A3(net55),
    .B1(net25),
    .Y(_07127_));
 sky130_fd_sc_hd__o31a_1 _17360_ (.A1(net33),
    .A2(net44),
    .A3(net55),
    .B1(net25),
    .X(_07128_));
 sky130_fd_sc_hd__o311a_4 _17361_ (.A1(net33),
    .A2(net44),
    .A3(net55),
    .B1(net25),
    .C1(_06881_),
    .X(_07129_));
 sky130_fd_sc_hd__nand2_1 _17362_ (.A(net60),
    .B(net22),
    .Y(_07130_));
 sky130_fd_sc_hd__a22oi_4 _17363_ (.A1(net59),
    .A2(net24),
    .B1(net25),
    .B2(net58),
    .Y(_07131_));
 sky130_fd_sc_hd__a22o_1 _17364_ (.A1(net59),
    .A2(net24),
    .B1(net25),
    .B2(net58),
    .X(_07132_));
 sky130_fd_sc_hd__and3_4 _17365_ (.A(net58),
    .B(net59),
    .C(net25),
    .X(_07133_));
 sky130_fd_sc_hd__nand3_4 _17366_ (.A(net58),
    .B(net59),
    .C(net25),
    .Y(_07134_));
 sky130_fd_sc_hd__and4_1 _17367_ (.A(net58),
    .B(net59),
    .C(net24),
    .D(net25),
    .X(_07135_));
 sky130_fd_sc_hd__nand4_4 _17368_ (.A(net58),
    .B(net59),
    .C(net24),
    .D(net25),
    .Y(_07137_));
 sky130_fd_sc_hd__o221ai_2 _17369_ (.A1(_01835_),
    .A2(_02196_),
    .B1(_02218_),
    .B2(_07134_),
    .C1(_07132_),
    .Y(_07138_));
 sky130_fd_sc_hd__o21bai_1 _17370_ (.A1(_07131_),
    .A2(_07135_),
    .B1_N(_07130_),
    .Y(_07139_));
 sky130_fd_sc_hd__a22oi_4 _17371_ (.A1(net60),
    .A2(net22),
    .B1(_07132_),
    .B2(_07137_),
    .Y(_07140_));
 sky130_fd_sc_hd__nand3_1 _17372_ (.A(_07137_),
    .B(net22),
    .C(net60),
    .Y(_07141_));
 sky130_fd_sc_hd__o211ai_2 _17373_ (.A1(_06880_),
    .A2(_07127_),
    .B1(_07138_),
    .C1(_07139_),
    .Y(_07142_));
 sky130_fd_sc_hd__o21ai_4 _17374_ (.A1(_07131_),
    .A2(_07141_),
    .B1(_07129_),
    .Y(_07143_));
 sky130_fd_sc_hd__o21a_1 _17375_ (.A1(_07140_),
    .A2(_07143_),
    .B1(_07142_),
    .X(_07144_));
 sky130_fd_sc_hd__o21ai_4 _17376_ (.A1(_07140_),
    .A2(_07143_),
    .B1(_07142_),
    .Y(_07145_));
 sky130_fd_sc_hd__o32a_2 _17377_ (.A1(_01737_),
    .A2(_01780_),
    .A3(_06338_),
    .B1(_06869_),
    .B2(_06878_),
    .X(_07146_));
 sky130_fd_sc_hd__o22ai_2 _17378_ (.A1(_01780_),
    .A2(_06341_),
    .B1(_06869_),
    .B2(_06878_),
    .Y(_07148_));
 sky130_fd_sc_hd__nand2_2 _17379_ (.A(_07148_),
    .B(_07144_),
    .Y(_07149_));
 sky130_fd_sc_hd__o311a_2 _17380_ (.A1(_01759_),
    .A2(_01780_),
    .A3(_06011_),
    .B1(_06886_),
    .C1(_07145_),
    .X(_07150_));
 sky130_fd_sc_hd__o211ai_4 _17381_ (.A1(_01780_),
    .A2(_06341_),
    .B1(_06886_),
    .C1(_07145_),
    .Y(_07151_));
 sky130_fd_sc_hd__o21ai_2 _17382_ (.A1(_06859_),
    .A2(_06861_),
    .B1(_06860_),
    .Y(_07152_));
 sky130_fd_sc_hd__o21a_1 _17383_ (.A1(_06859_),
    .A2(_06861_),
    .B1(_06860_),
    .X(_07153_));
 sky130_fd_sc_hd__nand2_1 _17384_ (.A(net63),
    .B(net19),
    .Y(_07154_));
 sky130_fd_sc_hd__a22oi_2 _17385_ (.A1(net62),
    .A2(net20),
    .B1(net21),
    .B2(net61),
    .Y(_07155_));
 sky130_fd_sc_hd__a22o_1 _17386_ (.A1(net62),
    .A2(net20),
    .B1(net21),
    .B2(net61),
    .X(_07156_));
 sky130_fd_sc_hd__and4_2 _17387_ (.A(net61),
    .B(net62),
    .C(net20),
    .D(net21),
    .X(_07157_));
 sky130_fd_sc_hd__nand4_2 _17388_ (.A(net61),
    .B(net62),
    .C(net20),
    .D(net21),
    .Y(_07159_));
 sky130_fd_sc_hd__o211ai_2 _17389_ (.A1(_01890_),
    .A2(_02142_),
    .B1(_07156_),
    .C1(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__o21bai_1 _17390_ (.A1(_07155_),
    .A2(_07157_),
    .B1_N(_07154_),
    .Y(_07161_));
 sky130_fd_sc_hd__o21ai_2 _17391_ (.A1(_07155_),
    .A2(_07157_),
    .B1(_07154_),
    .Y(_07162_));
 sky130_fd_sc_hd__nand4_2 _17392_ (.A(_07156_),
    .B(_07159_),
    .C(net63),
    .D(net19),
    .Y(_07163_));
 sky130_fd_sc_hd__a21oi_1 _17393_ (.A1(_07162_),
    .A2(_07163_),
    .B1(_07152_),
    .Y(_07164_));
 sky130_fd_sc_hd__nand3_4 _17394_ (.A(_07153_),
    .B(_07160_),
    .C(_07161_),
    .Y(_07165_));
 sky130_fd_sc_hd__nand3_4 _17395_ (.A(_07162_),
    .B(_07163_),
    .C(_07152_),
    .Y(_07166_));
 sky130_fd_sc_hd__o22a_1 _17396_ (.A1(_01890_),
    .A2(_02131_),
    .B1(_02163_),
    .B2(_06366_),
    .X(_07167_));
 sky130_fd_sc_hd__and3_1 _17397_ (.A(_06838_),
    .B(net18),
    .C(net63),
    .X(_07168_));
 sky130_fd_sc_hd__a31o_1 _17398_ (.A1(_06838_),
    .A2(net18),
    .A3(net63),
    .B1(_06839_),
    .X(_07170_));
 sky130_fd_sc_hd__o22a_1 _17399_ (.A1(_02163_),
    .A2(_06366_),
    .B1(_06836_),
    .B2(_06837_),
    .X(_07171_));
 sky130_fd_sc_hd__a21oi_1 _17400_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07170_),
    .Y(_07172_));
 sky130_fd_sc_hd__o2bb2ai_1 _17401_ (.A1_N(_07165_),
    .A2_N(_07166_),
    .B1(_07167_),
    .B2(_06837_),
    .Y(_07173_));
 sky130_fd_sc_hd__and3_1 _17402_ (.A(_07165_),
    .B(_07166_),
    .C(_07170_),
    .X(_07174_));
 sky130_fd_sc_hd__o211ai_1 _17403_ (.A1(_06839_),
    .A2(_07168_),
    .B1(_07166_),
    .C1(_07165_),
    .Y(_07175_));
 sky130_fd_sc_hd__and3_1 _17404_ (.A(_07165_),
    .B(_07166_),
    .C(_07171_),
    .X(_07176_));
 sky130_fd_sc_hd__o211ai_1 _17405_ (.A1(_06837_),
    .A2(_07167_),
    .B1(_07166_),
    .C1(_07165_),
    .Y(_07177_));
 sky130_fd_sc_hd__o2bb2a_1 _17406_ (.A1_N(_07165_),
    .A2_N(_07166_),
    .B1(_07168_),
    .B2(_06839_),
    .X(_07178_));
 sky130_fd_sc_hd__o2bb2ai_1 _17407_ (.A1_N(_07165_),
    .A2_N(_07166_),
    .B1(_07168_),
    .B2(_06839_),
    .Y(_07179_));
 sky130_fd_sc_hd__nand2_1 _17408_ (.A(_07173_),
    .B(_07175_),
    .Y(_07181_));
 sky130_fd_sc_hd__o211ai_2 _17409_ (.A1(_07172_),
    .A2(_07174_),
    .B1(_07149_),
    .C1(_07151_),
    .Y(_07182_));
 sky130_fd_sc_hd__o2bb2ai_1 _17410_ (.A1_N(_07149_),
    .A2_N(_07151_),
    .B1(_07176_),
    .B2(_07178_),
    .Y(_07183_));
 sky130_fd_sc_hd__o2bb2ai_2 _17411_ (.A1_N(_07149_),
    .A2_N(_07151_),
    .B1(_07172_),
    .B2(_07174_),
    .Y(_07184_));
 sky130_fd_sc_hd__a22o_1 _17412_ (.A1(_07148_),
    .A2(_07144_),
    .B1(_07179_),
    .B2(_07177_),
    .X(_07185_));
 sky130_fd_sc_hd__o221a_1 _17413_ (.A1(_07145_),
    .A2(_07146_),
    .B1(_07176_),
    .B2(_07178_),
    .C1(_07151_),
    .X(_07186_));
 sky130_fd_sc_hd__o221ai_4 _17414_ (.A1(_07145_),
    .A2(_07146_),
    .B1(_07176_),
    .B2(_07178_),
    .C1(_07151_),
    .Y(_07187_));
 sky130_fd_sc_hd__o2111ai_4 _17415_ (.A1(_06858_),
    .A2(_06890_),
    .B1(_06893_),
    .C1(_07182_),
    .D1(_07183_),
    .Y(_07188_));
 sky130_fd_sc_hd__o21ai_1 _17416_ (.A1(_06892_),
    .A2(_06897_),
    .B1(_07184_),
    .Y(_07189_));
 sky130_fd_sc_hd__o221a_2 _17417_ (.A1(_07150_),
    .A2(_07185_),
    .B1(_06892_),
    .B2(_06897_),
    .C1(_07184_),
    .X(_07190_));
 sky130_fd_sc_hd__o211ai_2 _17418_ (.A1(_07150_),
    .A2(_07185_),
    .B1(_07184_),
    .C1(_07126_),
    .Y(_07192_));
 sky130_fd_sc_hd__o21ai_4 _17419_ (.A1(_07120_),
    .A2(_07121_),
    .B1(_07188_),
    .Y(_07193_));
 sky130_fd_sc_hd__o211a_1 _17420_ (.A1(_07120_),
    .A2(_07121_),
    .B1(_07188_),
    .C1(_07192_),
    .X(_07194_));
 sky130_fd_sc_hd__a31o_1 _17421_ (.A1(_07126_),
    .A2(_07184_),
    .A3(_07187_),
    .B1(_07193_),
    .X(_07195_));
 sky130_fd_sc_hd__a2bb2oi_2 _17422_ (.A1_N(_07122_),
    .A2_N(_07124_),
    .B1(_07188_),
    .B2(_07192_),
    .Y(_07196_));
 sky130_fd_sc_hd__a2bb2o_2 _17423_ (.A1_N(_07122_),
    .A2_N(_07124_),
    .B1(_07188_),
    .B2(_07192_),
    .X(_07197_));
 sky130_fd_sc_hd__o21ai_2 _17424_ (.A1(_07190_),
    .A2(_07193_),
    .B1(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__a21oi_1 _17425_ (.A1(_06901_),
    .A2(_06907_),
    .B1(_07196_),
    .Y(_07199_));
 sky130_fd_sc_hd__o221a_2 _17426_ (.A1(_07190_),
    .A2(_07193_),
    .B1(_06900_),
    .B2(_06905_),
    .C1(_07197_),
    .X(_07200_));
 sky130_fd_sc_hd__o221ai_4 _17427_ (.A1(_07190_),
    .A2(_07193_),
    .B1(_06900_),
    .B2(_06905_),
    .C1(_07197_),
    .Y(_07201_));
 sky130_fd_sc_hd__o21ai_4 _17428_ (.A1(_07194_),
    .A2(_07196_),
    .B1(_06910_),
    .Y(_07203_));
 sky130_fd_sc_hd__a21bo_1 _17429_ (.A1(_06734_),
    .A2(_06768_),
    .B1_N(_06735_),
    .X(_07204_));
 sky130_fd_sc_hd__a21boi_4 _17430_ (.A1(_06734_),
    .A2(_06768_),
    .B1_N(_06735_),
    .Y(_07205_));
 sky130_fd_sc_hd__a31oi_4 _17431_ (.A1(_06820_),
    .A2(_06821_),
    .A3(_06822_),
    .B1(_06827_),
    .Y(_07206_));
 sky130_fd_sc_hd__a31oi_4 _17432_ (.A1(_06419_),
    .A2(_06435_),
    .A3(_06826_),
    .B1(_06824_),
    .Y(_07207_));
 sky130_fd_sc_hd__o21ai_2 _17433_ (.A1(_06737_),
    .A2(_06738_),
    .B1(_06742_),
    .Y(_07208_));
 sky130_fd_sc_hd__nand2_1 _17434_ (.A(net6),
    .B(net45),
    .Y(_07209_));
 sky130_fd_sc_hd__a22oi_4 _17435_ (.A1(net8),
    .A2(net42),
    .B1(net43),
    .B2(net7),
    .Y(_07210_));
 sky130_fd_sc_hd__a22o_1 _17436_ (.A1(net8),
    .A2(net42),
    .B1(net43),
    .B2(net7),
    .X(_07211_));
 sky130_fd_sc_hd__and4_2 _17437_ (.A(net7),
    .B(net8),
    .C(net42),
    .D(net43),
    .X(_07212_));
 sky130_fd_sc_hd__nand4_1 _17438_ (.A(net7),
    .B(net8),
    .C(net42),
    .D(net43),
    .Y(_07214_));
 sky130_fd_sc_hd__o211ai_2 _17439_ (.A1(_01966_),
    .A2(_02054_),
    .B1(_07211_),
    .C1(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__o21bai_2 _17440_ (.A1(_07210_),
    .A2(_07212_),
    .B1_N(_07209_),
    .Y(_07216_));
 sky130_fd_sc_hd__o22a_2 _17441_ (.A1(_01966_),
    .A2(_02054_),
    .B1(_07210_),
    .B2(_07212_),
    .X(_07217_));
 sky130_fd_sc_hd__nand3b_4 _17442_ (.A_N(_07208_),
    .B(_07215_),
    .C(_07216_),
    .Y(_07218_));
 sky130_fd_sc_hd__o31ai_4 _17443_ (.A1(_07209_),
    .A2(_07210_),
    .A3(_07212_),
    .B1(_07208_),
    .Y(_07219_));
 sky130_fd_sc_hd__nor2_1 _17444_ (.A(_07217_),
    .B(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__a21bo_1 _17445_ (.A1(_07215_),
    .A2(_07216_),
    .B1_N(_07208_),
    .X(_07221_));
 sky130_fd_sc_hd__nand2_1 _17446_ (.A(net3),
    .B(net48),
    .Y(_07222_));
 sky130_fd_sc_hd__nand4_4 _17447_ (.A(net4),
    .B(net5),
    .C(net46),
    .D(net47),
    .Y(_07223_));
 sky130_fd_sc_hd__a22oi_1 _17448_ (.A1(net5),
    .A2(net46),
    .B1(net47),
    .B2(net4),
    .Y(_07225_));
 sky130_fd_sc_hd__a22o_1 _17449_ (.A1(net5),
    .A2(net46),
    .B1(net47),
    .B2(net4),
    .X(_07226_));
 sky130_fd_sc_hd__o211ai_2 _17450_ (.A1(_01923_),
    .A2(_02109_),
    .B1(_07223_),
    .C1(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__a21o_1 _17451_ (.A1(_07223_),
    .A2(_07226_),
    .B1(_07222_),
    .X(_07228_));
 sky130_fd_sc_hd__a22o_1 _17452_ (.A1(net3),
    .A2(net48),
    .B1(_07223_),
    .B2(_07226_),
    .X(_07229_));
 sky130_fd_sc_hd__nand4_1 _17453_ (.A(_07226_),
    .B(net48),
    .C(net3),
    .D(_07223_),
    .Y(_07230_));
 sky130_fd_sc_hd__nand2_1 _17454_ (.A(_07229_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__nand2_1 _17455_ (.A(_07227_),
    .B(_07228_),
    .Y(_07232_));
 sky130_fd_sc_hd__a21oi_1 _17456_ (.A1(_07218_),
    .A2(_07221_),
    .B1(_07231_),
    .Y(_07233_));
 sky130_fd_sc_hd__and3_1 _17457_ (.A(_07218_),
    .B(_07221_),
    .C(_07231_),
    .X(_07234_));
 sky130_fd_sc_hd__o2111ai_2 _17458_ (.A1(_07217_),
    .A2(_07219_),
    .B1(_07227_),
    .C1(_07228_),
    .D1(_07218_),
    .Y(_07236_));
 sky130_fd_sc_hd__a22o_1 _17459_ (.A1(_07218_),
    .A2(_07221_),
    .B1(_07229_),
    .B2(_07230_),
    .X(_07237_));
 sky130_fd_sc_hd__nand2_1 _17460_ (.A(_07218_),
    .B(_07232_),
    .Y(_07238_));
 sky130_fd_sc_hd__o21ai_2 _17461_ (.A1(_07220_),
    .A2(_07238_),
    .B1(_07237_),
    .Y(_07239_));
 sky130_fd_sc_hd__a21oi_1 _17462_ (.A1(_06728_),
    .A2(_06712_),
    .B1(_06725_),
    .Y(_07240_));
 sky130_fd_sc_hd__o21a_1 _17463_ (.A1(_01988_),
    .A2(_02010_),
    .B1(_06720_),
    .X(_07241_));
 sky130_fd_sc_hd__and3_1 _17464_ (.A(_06717_),
    .B(net41),
    .C(net8),
    .X(_07242_));
 sky130_fd_sc_hd__o31a_1 _17465_ (.A1(_01988_),
    .A2(_02010_),
    .A3(_06716_),
    .B1(_06720_),
    .X(_07243_));
 sky130_fd_sc_hd__a21oi_2 _17466_ (.A1(_06422_),
    .A2(_06805_),
    .B1(_06804_),
    .Y(_07244_));
 sky130_fd_sc_hd__o21ai_1 _17467_ (.A1(_06804_),
    .A2(_06806_),
    .B1(_06810_),
    .Y(_07245_));
 sky130_fd_sc_hd__o21a_1 _17468_ (.A1(_06804_),
    .A2(_06806_),
    .B1(_06810_),
    .X(_07247_));
 sky130_fd_sc_hd__nor2_1 _17469_ (.A(_01999_),
    .B(_02010_),
    .Y(_07248_));
 sky130_fd_sc_hd__a22oi_4 _17470_ (.A1(net40),
    .A2(net10),
    .B1(net11),
    .B2(net39),
    .Y(_07249_));
 sky130_fd_sc_hd__a22o_1 _17471_ (.A1(net40),
    .A2(net10),
    .B1(net11),
    .B2(net39),
    .X(_07250_));
 sky130_fd_sc_hd__and4_1 _17472_ (.A(net39),
    .B(net40),
    .C(net10),
    .D(net11),
    .X(_07251_));
 sky130_fd_sc_hd__nand4_2 _17473_ (.A(net39),
    .B(net40),
    .C(net10),
    .D(net11),
    .Y(_07252_));
 sky130_fd_sc_hd__o211ai_2 _17474_ (.A1(_01999_),
    .A2(_02010_),
    .B1(_07250_),
    .C1(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__o21ai_1 _17475_ (.A1(_07249_),
    .A2(_07251_),
    .B1(_07248_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand4_2 _17476_ (.A(_07250_),
    .B(_07252_),
    .C(net9),
    .D(net41),
    .Y(_07255_));
 sky130_fd_sc_hd__o22ai_4 _17477_ (.A1(_01999_),
    .A2(_02010_),
    .B1(_07249_),
    .B2(_07251_),
    .Y(_07256_));
 sky130_fd_sc_hd__o211a_1 _17478_ (.A1(_06809_),
    .A2(_07244_),
    .B1(_07255_),
    .C1(_07256_),
    .X(_07258_));
 sky130_fd_sc_hd__o211ai_4 _17479_ (.A1(_06809_),
    .A2(_07244_),
    .B1(_07255_),
    .C1(_07256_),
    .Y(_07259_));
 sky130_fd_sc_hd__a21oi_1 _17480_ (.A1(_07255_),
    .A2(_07256_),
    .B1(_07245_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand3_2 _17481_ (.A(_07247_),
    .B(_07253_),
    .C(_07254_),
    .Y(_07261_));
 sky130_fd_sc_hd__a31oi_2 _17482_ (.A1(_07247_),
    .A2(_07253_),
    .A3(_07254_),
    .B1(_07243_),
    .Y(_07262_));
 sky130_fd_sc_hd__a2bb2oi_2 _17483_ (.A1_N(_06718_),
    .A2_N(_07242_),
    .B1(_07259_),
    .B2(_07261_),
    .Y(_07263_));
 sky130_fd_sc_hd__o22ai_2 _17484_ (.A1(_06718_),
    .A2(_07242_),
    .B1(_07258_),
    .B2(_07260_),
    .Y(_07264_));
 sky130_fd_sc_hd__o211a_1 _17485_ (.A1(_06716_),
    .A2(_07241_),
    .B1(_07259_),
    .C1(_07261_),
    .X(_07265_));
 sky130_fd_sc_hd__o2111ai_2 _17486_ (.A1(_06715_),
    .A2(_06716_),
    .B1(_06720_),
    .C1(_07259_),
    .D1(_07261_),
    .Y(_07266_));
 sky130_fd_sc_hd__a21oi_1 _17487_ (.A1(_07264_),
    .A2(_07266_),
    .B1(_07240_),
    .Y(_07267_));
 sky130_fd_sc_hd__o21bai_4 _17488_ (.A1(_07263_),
    .A2(_07265_),
    .B1_N(_07240_),
    .Y(_07269_));
 sky130_fd_sc_hd__nor3b_2 _17489_ (.A(_07263_),
    .B(_07265_),
    .C_N(_07240_),
    .Y(_07270_));
 sky130_fd_sc_hd__nand4_2 _17490_ (.A(_06726_),
    .B(_06729_),
    .C(_07264_),
    .D(_07266_),
    .Y(_07271_));
 sky130_fd_sc_hd__o2111ai_4 _17491_ (.A1(_07238_),
    .A2(_07220_),
    .B1(_07237_),
    .C1(_07269_),
    .D1(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__o21ai_2 _17492_ (.A1(_07267_),
    .A2(_07270_),
    .B1(_07239_),
    .Y(_07273_));
 sky130_fd_sc_hd__nand4b_2 _17493_ (.A_N(_07233_),
    .B(_07236_),
    .C(_07269_),
    .D(_07271_),
    .Y(_07274_));
 sky130_fd_sc_hd__o22ai_2 _17494_ (.A1(_07233_),
    .A2(_07234_),
    .B1(_07267_),
    .B2(_07270_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand3_4 _17495_ (.A(_07273_),
    .B(_07207_),
    .C(_07272_),
    .Y(_07276_));
 sky130_fd_sc_hd__o211a_1 _17496_ (.A1(_06824_),
    .A2(_07206_),
    .B1(_07274_),
    .C1(_07275_),
    .X(_07277_));
 sky130_fd_sc_hd__o211ai_4 _17497_ (.A1(_06824_),
    .A2(_07206_),
    .B1(_07274_),
    .C1(_07275_),
    .Y(_07278_));
 sky130_fd_sc_hd__a21oi_2 _17498_ (.A1(_07276_),
    .A2(_07278_),
    .B1(_07204_),
    .Y(_07280_));
 sky130_fd_sc_hd__and3_1 _17499_ (.A(_07276_),
    .B(_07278_),
    .C(_07204_),
    .X(_07281_));
 sky130_fd_sc_hd__a21oi_2 _17500_ (.A1(_07276_),
    .A2(_07278_),
    .B1(_07205_),
    .Y(_07282_));
 sky130_fd_sc_hd__a21o_1 _17501_ (.A1(_07276_),
    .A2(_07278_),
    .B1(_07205_),
    .X(_07283_));
 sky130_fd_sc_hd__and3_1 _17502_ (.A(_07205_),
    .B(_07276_),
    .C(_07278_),
    .X(_07284_));
 sky130_fd_sc_hd__nand3_2 _17503_ (.A(_07205_),
    .B(_07276_),
    .C(_07278_),
    .Y(_07285_));
 sky130_fd_sc_hd__nand2_1 _17504_ (.A(_07283_),
    .B(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__o2bb2ai_2 _17505_ (.A1_N(_07201_),
    .A2_N(_07203_),
    .B1(_07282_),
    .B2(_07284_),
    .Y(_07287_));
 sky130_fd_sc_hd__o211ai_4 _17506_ (.A1(_07280_),
    .A2(_07281_),
    .B1(_07201_),
    .C1(_07203_),
    .Y(_07288_));
 sky130_fd_sc_hd__o2bb2ai_2 _17507_ (.A1_N(_07201_),
    .A2_N(_07203_),
    .B1(_07280_),
    .B2(_07281_),
    .Y(_07289_));
 sky130_fd_sc_hd__a22oi_4 _17508_ (.A1(_07283_),
    .A2(_07285_),
    .B1(_07198_),
    .B2(_06910_),
    .Y(_07291_));
 sky130_fd_sc_hd__o21ai_1 _17509_ (.A1(_07282_),
    .A2(_07284_),
    .B1(_07203_),
    .Y(_07292_));
 sky130_fd_sc_hd__and3_2 _17510_ (.A(_07286_),
    .B(_07203_),
    .C(_07201_),
    .X(_07293_));
 sky130_fd_sc_hd__o211ai_2 _17511_ (.A1(_07282_),
    .A2(_07284_),
    .B1(_07201_),
    .C1(_07203_),
    .Y(_07294_));
 sky130_fd_sc_hd__a32oi_4 _17512_ (.A1(_06904_),
    .A2(_06909_),
    .A3(_06912_),
    .B1(_06784_),
    .B2(_06783_),
    .Y(_07295_));
 sky130_fd_sc_hd__o22ai_4 _17513_ (.A1(_06908_),
    .A2(_06915_),
    .B1(_06913_),
    .B2(_06788_),
    .Y(_07296_));
 sky130_fd_sc_hd__a21oi_4 _17514_ (.A1(_07289_),
    .A2(_07294_),
    .B1(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__o211ai_4 _17515_ (.A1(_06913_),
    .A2(_07295_),
    .B1(_07288_),
    .C1(_07287_),
    .Y(_07298_));
 sky130_fd_sc_hd__nand2_2 _17516_ (.A(_07296_),
    .B(_07289_),
    .Y(_07299_));
 sky130_fd_sc_hd__o211a_2 _17517_ (.A1(_07200_),
    .A2(_07292_),
    .B1(_07289_),
    .C1(_07296_),
    .X(_07300_));
 sky130_fd_sc_hd__a22o_1 _17518_ (.A1(_06918_),
    .A2(_06919_),
    .B1(_07287_),
    .B2(_07288_),
    .X(_07302_));
 sky130_fd_sc_hd__o22ai_4 _17519_ (.A1(_07077_),
    .A2(_07078_),
    .B1(_07297_),
    .B2(_07300_),
    .Y(_07303_));
 sky130_fd_sc_hd__o221ai_4 _17520_ (.A1(_07072_),
    .A2(_07076_),
    .B1(_07293_),
    .B2(_07299_),
    .C1(_07298_),
    .Y(_07304_));
 sky130_fd_sc_hd__o21ai_2 _17521_ (.A1(_07077_),
    .A2(_07078_),
    .B1(_07298_),
    .Y(_07305_));
 sky130_fd_sc_hd__o211ai_1 _17522_ (.A1(_07077_),
    .A2(_07078_),
    .B1(_07298_),
    .C1(_07302_),
    .Y(_07306_));
 sky130_fd_sc_hd__o22ai_2 _17523_ (.A1(_07072_),
    .A2(_07076_),
    .B1(_07297_),
    .B2(_07300_),
    .Y(_07307_));
 sky130_fd_sc_hd__a22oi_4 _17524_ (.A1(_06926_),
    .A2(_06932_),
    .B1(_07303_),
    .B2(_07304_),
    .Y(_07308_));
 sky130_fd_sc_hd__o211ai_4 _17525_ (.A1(_07305_),
    .A2(_07300_),
    .B1(_06968_),
    .C1(_07307_),
    .Y(_07309_));
 sky130_fd_sc_hd__a21oi_1 _17526_ (.A1(_07306_),
    .A2(_07307_),
    .B1(_06968_),
    .Y(_07310_));
 sky130_fd_sc_hd__nand3_4 _17527_ (.A(_06967_),
    .B(_07303_),
    .C(_07304_),
    .Y(_07311_));
 sky130_fd_sc_hd__nand2_1 _17528_ (.A(_07309_),
    .B(_06965_),
    .Y(_07313_));
 sky130_fd_sc_hd__a31o_2 _17529_ (.A1(_06967_),
    .A2(_07303_),
    .A3(_07304_),
    .B1(_06965_),
    .X(_07314_));
 sky130_fd_sc_hd__and3_1 _17530_ (.A(_06966_),
    .B(_07309_),
    .C(_07311_),
    .X(_07315_));
 sky130_fd_sc_hd__a21oi_1 _17531_ (.A1(_06966_),
    .A2(_07311_),
    .B1(_07308_),
    .Y(_07316_));
 sky130_fd_sc_hd__o22ai_2 _17532_ (.A1(_06701_),
    .A2(_06706_),
    .B1(_07308_),
    .B2(_07310_),
    .Y(_07317_));
 sky130_fd_sc_hd__nand4_2 _17533_ (.A(_06702_),
    .B(_06707_),
    .C(_07309_),
    .D(_07311_),
    .Y(_07318_));
 sky130_fd_sc_hd__o21ai_2 _17534_ (.A1(_07308_),
    .A2(_07310_),
    .B1(_06965_),
    .Y(_07319_));
 sky130_fd_sc_hd__nand3_2 _17535_ (.A(_06964_),
    .B(_07317_),
    .C(_07318_),
    .Y(_07320_));
 sky130_fd_sc_hd__o21ai_1 _17536_ (.A1(_06934_),
    .A2(_06941_),
    .B1(_07319_),
    .Y(_07321_));
 sky130_fd_sc_hd__o221a_1 _17537_ (.A1(_06934_),
    .A2(_06941_),
    .B1(_07308_),
    .B2(_07314_),
    .C1(_07319_),
    .X(_07322_));
 sky130_fd_sc_hd__o221ai_4 _17538_ (.A1(_06934_),
    .A2(_06941_),
    .B1(_07308_),
    .B2(_07314_),
    .C1(_07319_),
    .Y(_07324_));
 sky130_fd_sc_hd__o31a_1 _17539_ (.A1(net12),
    .A2(_02240_),
    .A3(_05884_),
    .B1(_06639_),
    .X(_07325_));
 sky130_fd_sc_hd__nand2_1 _17540_ (.A(_06639_),
    .B(_06644_),
    .Y(_07326_));
 sky130_fd_sc_hd__inv_2 _17541_ (.A(_07326_),
    .Y(_07327_));
 sky130_fd_sc_hd__a21oi_1 _17542_ (.A1(_07320_),
    .A2(_07324_),
    .B1(_07326_),
    .Y(_07328_));
 sky130_fd_sc_hd__o2bb2ai_1 _17543_ (.A1_N(_07320_),
    .A2_N(_07324_),
    .B1(_07325_),
    .B2(_06637_),
    .Y(_07329_));
 sky130_fd_sc_hd__a31oi_2 _17544_ (.A1(_06964_),
    .A2(_07317_),
    .A3(_07318_),
    .B1(_07327_),
    .Y(_07330_));
 sky130_fd_sc_hd__and3_1 _17545_ (.A(_07320_),
    .B(_07324_),
    .C(_07326_),
    .X(_07331_));
 sky130_fd_sc_hd__o21ai_2 _17546_ (.A1(_07315_),
    .A2(_07321_),
    .B1(_07330_),
    .Y(_07332_));
 sky130_fd_sc_hd__a22oi_1 _17547_ (.A1(_06945_),
    .A2(_06963_),
    .B1(_07329_),
    .B2(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__o2bb2ai_1 _17548_ (.A1_N(_06945_),
    .A2_N(_06963_),
    .B1(_07328_),
    .B2(_07331_),
    .Y(_07335_));
 sky130_fd_sc_hd__o21a_1 _17549_ (.A1(_06946_),
    .A2(_06952_),
    .B1(_07329_),
    .X(_07336_));
 sky130_fd_sc_hd__o211ai_1 _17550_ (.A1(_06946_),
    .A2(_06952_),
    .B1(_07329_),
    .C1(_07332_),
    .Y(_07337_));
 sky130_fd_sc_hd__a21oi_1 _17551_ (.A1(_07336_),
    .A2(_07332_),
    .B1(_07333_),
    .Y(_07338_));
 sky130_fd_sc_hd__a21o_1 _17552_ (.A1(_07336_),
    .A2(_07332_),
    .B1(_07333_),
    .X(_07339_));
 sky130_fd_sc_hd__a32oi_4 _17553_ (.A1(_06954_),
    .A2(_06955_),
    .A3(_06957_),
    .B1(_06959_),
    .B2(_06586_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand4_1 _17554_ (.A(_06585_),
    .B(_06586_),
    .C(_06958_),
    .D(_06959_),
    .Y(_07341_));
 sky130_fd_sc_hd__a41oi_2 _17555_ (.A1(_06601_),
    .A2(_06958_),
    .A3(_06959_),
    .A4(_06587_),
    .B1(_07340_),
    .Y(_07342_));
 sky130_fd_sc_hd__xor2_1 _17556_ (.A(_07339_),
    .B(_07342_),
    .X(net92));
 sky130_fd_sc_hd__a21oi_2 _17557_ (.A1(_07079_),
    .A2(_07298_),
    .B1(_07300_),
    .Y(_07343_));
 sky130_fd_sc_hd__o22ai_4 _17558_ (.A1(_07293_),
    .A2(_07299_),
    .B1(_07297_),
    .B2(_07080_),
    .Y(_07345_));
 sky130_fd_sc_hd__a311o_1 _17559_ (.A1(_07126_),
    .A2(_07184_),
    .A3(_07187_),
    .B1(_07121_),
    .C1(_07120_),
    .X(_07346_));
 sky130_fd_sc_hd__o21ai_4 _17560_ (.A1(_07186_),
    .A2(_07189_),
    .B1(_07193_),
    .Y(_07347_));
 sky130_fd_sc_hd__o21ai_4 _17561_ (.A1(_07084_),
    .A2(_07085_),
    .B1(_07088_),
    .Y(_07348_));
 sky130_fd_sc_hd__nand2_1 _17562_ (.A(net35),
    .B(net17),
    .Y(_07349_));
 sky130_fd_sc_hd__a22oi_2 _17563_ (.A1(net34),
    .A2(net18),
    .B1(net19),
    .B2(net64),
    .Y(_07350_));
 sky130_fd_sc_hd__a22o_1 _17564_ (.A1(net34),
    .A2(net18),
    .B1(net19),
    .B2(net64),
    .X(_07351_));
 sky130_fd_sc_hd__and4_1 _17565_ (.A(net64),
    .B(net34),
    .C(net18),
    .D(net19),
    .X(_07352_));
 sky130_fd_sc_hd__nand4_4 _17566_ (.A(net64),
    .B(net34),
    .C(net18),
    .D(net19),
    .Y(_07353_));
 sky130_fd_sc_hd__nand3_1 _17567_ (.A(_07349_),
    .B(_07351_),
    .C(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__o21bai_1 _17568_ (.A1(_07350_),
    .A2(_07352_),
    .B1_N(_07349_),
    .Y(_07356_));
 sky130_fd_sc_hd__a22o_1 _17569_ (.A1(net35),
    .A2(net17),
    .B1(_07351_),
    .B2(_07353_),
    .X(_07357_));
 sky130_fd_sc_hd__nand4_4 _17570_ (.A(_07351_),
    .B(_07353_),
    .C(net35),
    .D(net17),
    .Y(_07358_));
 sky130_fd_sc_hd__nand3b_4 _17571_ (.A_N(_07348_),
    .B(_07354_),
    .C(_07356_),
    .Y(_07359_));
 sky130_fd_sc_hd__nand3_2 _17572_ (.A(_07357_),
    .B(_07358_),
    .C(_07348_),
    .Y(_07360_));
 sky130_fd_sc_hd__nand2_1 _17573_ (.A(_07359_),
    .B(_07360_),
    .Y(_07361_));
 sky130_fd_sc_hd__nand2_2 _17574_ (.A(net38),
    .B(net14),
    .Y(_07362_));
 sky130_fd_sc_hd__nand2_1 _17575_ (.A(net36),
    .B(net16),
    .Y(_07363_));
 sky130_fd_sc_hd__a22oi_4 _17576_ (.A1(net37),
    .A2(net15),
    .B1(net16),
    .B2(net36),
    .Y(_07364_));
 sky130_fd_sc_hd__and4_1 _17577_ (.A(net36),
    .B(net37),
    .C(net15),
    .D(net16),
    .X(_07365_));
 sky130_fd_sc_hd__nand4_2 _17578_ (.A(net36),
    .B(net37),
    .C(net15),
    .D(net16),
    .Y(_07367_));
 sky130_fd_sc_hd__o21ai_1 _17579_ (.A1(_07364_),
    .A2(_07365_),
    .B1(_07362_),
    .Y(_07368_));
 sky130_fd_sc_hd__a41o_1 _17580_ (.A1(net36),
    .A2(net37),
    .A3(net15),
    .A4(net16),
    .B1(_07362_),
    .X(_07369_));
 sky130_fd_sc_hd__o21a_2 _17581_ (.A1(_07364_),
    .A2(_07369_),
    .B1(_07368_),
    .X(_07370_));
 sky130_fd_sc_hd__nand2_1 _17582_ (.A(_07361_),
    .B(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__nand3b_1 _17583_ (.A_N(_07370_),
    .B(_07360_),
    .C(_07359_),
    .Y(_07372_));
 sky130_fd_sc_hd__a21o_1 _17584_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07370_),
    .X(_07373_));
 sky130_fd_sc_hd__nand2_1 _17585_ (.A(_07359_),
    .B(_07370_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand3_1 _17586_ (.A(_07359_),
    .B(_07360_),
    .C(_07370_),
    .Y(_07375_));
 sky130_fd_sc_hd__nand2_1 _17587_ (.A(_07373_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__o21ai_1 _17588_ (.A1(_07171_),
    .A2(_07164_),
    .B1(_07166_),
    .Y(_07378_));
 sky130_fd_sc_hd__a21boi_2 _17589_ (.A1(_07165_),
    .A2(_07170_),
    .B1_N(_07166_),
    .Y(_07379_));
 sky130_fd_sc_hd__nand3_2 _17590_ (.A(_07371_),
    .B(_07372_),
    .C(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__nand3_2 _17591_ (.A(_07373_),
    .B(_07375_),
    .C(_07378_),
    .Y(_07381_));
 sky130_fd_sc_hd__a21bo_2 _17592_ (.A1(_07094_),
    .A2(_07107_),
    .B1_N(_07095_),
    .X(_07382_));
 sky130_fd_sc_hd__and3_1 _17593_ (.A(_07380_),
    .B(_07381_),
    .C(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__nand3_4 _17594_ (.A(_07380_),
    .B(_07381_),
    .C(_07382_),
    .Y(_07384_));
 sky130_fd_sc_hd__a21oi_1 _17595_ (.A1(_07380_),
    .A2(_07381_),
    .B1(_07382_),
    .Y(_07385_));
 sky130_fd_sc_hd__a21o_1 _17596_ (.A1(_07380_),
    .A2(_07381_),
    .B1(_07382_),
    .X(_07386_));
 sky130_fd_sc_hd__o21ai_4 _17597_ (.A1(net58),
    .A2(net59),
    .B1(net25),
    .Y(_07387_));
 sky130_fd_sc_hd__o21a_4 _17598_ (.A1(net58),
    .A2(net59),
    .B1(net25),
    .X(_07389_));
 sky130_fd_sc_hd__nand2_1 _17599_ (.A(_07134_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__a22oi_2 _17600_ (.A1(net60),
    .A2(net24),
    .B1(_07134_),
    .B2(_07389_),
    .Y(_07391_));
 sky130_fd_sc_hd__o22ai_4 _17601_ (.A1(_01835_),
    .A2(_02218_),
    .B1(_07133_),
    .B2(_07387_),
    .Y(_07392_));
 sky130_fd_sc_hd__and4_2 _17602_ (.A(_07389_),
    .B(net24),
    .C(net60),
    .D(_07134_),
    .X(_07393_));
 sky130_fd_sc_hd__nand4_2 _17603_ (.A(_07389_),
    .B(net24),
    .C(net60),
    .D(_07134_),
    .Y(_07394_));
 sky130_fd_sc_hd__o22ai_4 _17604_ (.A1(_06880_),
    .A2(_07127_),
    .B1(_07391_),
    .B2(_07393_),
    .Y(_07395_));
 sky130_fd_sc_hd__nand2_1 _17605_ (.A(_07392_),
    .B(_07129_),
    .Y(_07396_));
 sky130_fd_sc_hd__nand3_2 _17606_ (.A(_07392_),
    .B(_07394_),
    .C(_07129_),
    .Y(_07397_));
 sky130_fd_sc_hd__o22ai_4 _17607_ (.A1(_01780_),
    .A2(_06341_),
    .B1(_07140_),
    .B2(_07143_),
    .Y(_07398_));
 sky130_fd_sc_hd__a21oi_4 _17608_ (.A1(_07395_),
    .A2(_07397_),
    .B1(_07398_),
    .Y(_07400_));
 sky130_fd_sc_hd__a21o_1 _17609_ (.A1(_07395_),
    .A2(_07397_),
    .B1(_07398_),
    .X(_07401_));
 sky130_fd_sc_hd__o211a_2 _17610_ (.A1(_07393_),
    .A2(_07396_),
    .B1(_07398_),
    .C1(_07395_),
    .X(_07402_));
 sky130_fd_sc_hd__o211ai_4 _17611_ (.A1(_07393_),
    .A2(_07396_),
    .B1(_07398_),
    .C1(_07395_),
    .Y(_07403_));
 sky130_fd_sc_hd__o21ai_2 _17612_ (.A1(_07130_),
    .A2(_07131_),
    .B1(_07137_),
    .Y(_07404_));
 sky130_fd_sc_hd__o22a_2 _17613_ (.A1(_02218_),
    .A2(_07134_),
    .B1(_07130_),
    .B2(_07131_),
    .X(_07405_));
 sky130_fd_sc_hd__nand2_1 _17614_ (.A(net63),
    .B(net20),
    .Y(_07406_));
 sky130_fd_sc_hd__a22oi_4 _17615_ (.A1(net62),
    .A2(net21),
    .B1(net22),
    .B2(net61),
    .Y(_07407_));
 sky130_fd_sc_hd__a22o_1 _17616_ (.A1(net62),
    .A2(net21),
    .B1(net22),
    .B2(net61),
    .X(_07408_));
 sky130_fd_sc_hd__and4_2 _17617_ (.A(net61),
    .B(net62),
    .C(net21),
    .D(net22),
    .X(_07409_));
 sky130_fd_sc_hd__nand4_4 _17618_ (.A(net61),
    .B(net62),
    .C(net21),
    .D(net22),
    .Y(_07411_));
 sky130_fd_sc_hd__o211ai_4 _17619_ (.A1(_01890_),
    .A2(_02163_),
    .B1(_07408_),
    .C1(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__o21bai_2 _17620_ (.A1(_07407_),
    .A2(_07409_),
    .B1_N(_07406_),
    .Y(_07413_));
 sky130_fd_sc_hd__o21ai_2 _17621_ (.A1(_07407_),
    .A2(_07409_),
    .B1(_07406_),
    .Y(_07414_));
 sky130_fd_sc_hd__nand4_2 _17622_ (.A(_07408_),
    .B(_07411_),
    .C(net63),
    .D(net20),
    .Y(_07415_));
 sky130_fd_sc_hd__nand3_2 _17623_ (.A(_07405_),
    .B(_07412_),
    .C(_07413_),
    .Y(_07416_));
 sky130_fd_sc_hd__and3_4 _17624_ (.A(_07414_),
    .B(_07415_),
    .C(_07404_),
    .X(_07417_));
 sky130_fd_sc_hd__nand3_2 _17625_ (.A(_07414_),
    .B(_07415_),
    .C(_07404_),
    .Y(_07418_));
 sky130_fd_sc_hd__and3_1 _17626_ (.A(_07156_),
    .B(net19),
    .C(net63),
    .X(_07419_));
 sky130_fd_sc_hd__a31o_1 _17627_ (.A1(_07156_),
    .A2(net19),
    .A3(net63),
    .B1(_07157_),
    .X(_07420_));
 sky130_fd_sc_hd__o31a_1 _17628_ (.A1(_01890_),
    .A2(_02142_),
    .A3(_07155_),
    .B1(_07159_),
    .X(_07422_));
 sky130_fd_sc_hd__a21oi_2 _17629_ (.A1(_07416_),
    .A2(_07418_),
    .B1(_07420_),
    .Y(_07423_));
 sky130_fd_sc_hd__a21o_2 _17630_ (.A1(_07416_),
    .A2(_07418_),
    .B1(_07420_),
    .X(_07424_));
 sky130_fd_sc_hd__a31oi_4 _17631_ (.A1(_07405_),
    .A2(_07412_),
    .A3(_07413_),
    .B1(_07422_),
    .Y(_07425_));
 sky130_fd_sc_hd__a31o_1 _17632_ (.A1(_07405_),
    .A2(_07412_),
    .A3(_07413_),
    .B1(_07422_),
    .X(_07426_));
 sky130_fd_sc_hd__o211a_1 _17633_ (.A1(_07157_),
    .A2(_07419_),
    .B1(_07418_),
    .C1(_07416_),
    .X(_07427_));
 sky130_fd_sc_hd__o211ai_2 _17634_ (.A1(_07157_),
    .A2(_07419_),
    .B1(_07418_),
    .C1(_07416_),
    .Y(_07428_));
 sky130_fd_sc_hd__o221ai_4 _17635_ (.A1(_07417_),
    .A2(_07426_),
    .B1(_07400_),
    .B2(_07402_),
    .C1(_07424_),
    .Y(_07429_));
 sky130_fd_sc_hd__o211ai_2 _17636_ (.A1(_07423_),
    .A2(_07427_),
    .B1(_07401_),
    .C1(_07403_),
    .Y(_07430_));
 sky130_fd_sc_hd__o22ai_4 _17637_ (.A1(_07400_),
    .A2(_07402_),
    .B1(_07423_),
    .B2(_07427_),
    .Y(_07431_));
 sky130_fd_sc_hd__o2111ai_4 _17638_ (.A1(_07417_),
    .A2(_07426_),
    .B1(_07424_),
    .C1(_07401_),
    .D1(_07403_),
    .Y(_07433_));
 sky130_fd_sc_hd__nand2_1 _17639_ (.A(_07431_),
    .B(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__a22o_1 _17640_ (.A1(_07148_),
    .A2(_07144_),
    .B1(_07175_),
    .B2(_07173_),
    .X(_07435_));
 sky130_fd_sc_hd__a31o_1 _17641_ (.A1(_07149_),
    .A2(_07177_),
    .A3(_07179_),
    .B1(_07150_),
    .X(_07436_));
 sky130_fd_sc_hd__and4_2 _17642_ (.A(_07151_),
    .B(_07431_),
    .C(_07433_),
    .D(_07435_),
    .X(_07437_));
 sky130_fd_sc_hd__nand4_4 _17643_ (.A(_07151_),
    .B(_07431_),
    .C(_07433_),
    .D(_07435_),
    .Y(_07438_));
 sky130_fd_sc_hd__o2111ai_4 _17644_ (.A1(_07181_),
    .A2(_07150_),
    .B1(_07149_),
    .C1(_07430_),
    .D1(_07429_),
    .Y(_07439_));
 sky130_fd_sc_hd__nand2_1 _17645_ (.A(_07438_),
    .B(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__a22oi_2 _17646_ (.A1(_07384_),
    .A2(_07386_),
    .B1(_07438_),
    .B2(_07439_),
    .Y(_07441_));
 sky130_fd_sc_hd__o21ai_4 _17647_ (.A1(_07383_),
    .A2(_07385_),
    .B1(_07440_),
    .Y(_07442_));
 sky130_fd_sc_hd__nand3_4 _17648_ (.A(_07384_),
    .B(_07386_),
    .C(_07439_),
    .Y(_07444_));
 sky130_fd_sc_hd__and4_1 _17649_ (.A(_07384_),
    .B(_07386_),
    .C(_07438_),
    .D(_07439_),
    .X(_07445_));
 sky130_fd_sc_hd__nand4_1 _17650_ (.A(_07384_),
    .B(_07386_),
    .C(_07438_),
    .D(_07439_),
    .Y(_07446_));
 sky130_fd_sc_hd__o21a_1 _17651_ (.A1(_07437_),
    .A2(_07444_),
    .B1(_07442_),
    .X(_07447_));
 sky130_fd_sc_hd__o211a_1 _17652_ (.A1(_07437_),
    .A2(_07444_),
    .B1(_07442_),
    .C1(_07347_),
    .X(_07448_));
 sky130_fd_sc_hd__o211ai_4 _17653_ (.A1(_07437_),
    .A2(_07444_),
    .B1(_07442_),
    .C1(_07347_),
    .Y(_07449_));
 sky130_fd_sc_hd__a21oi_2 _17654_ (.A1(_07442_),
    .A2(_07446_),
    .B1(_07347_),
    .Y(_07450_));
 sky130_fd_sc_hd__o2bb2ai_4 _17655_ (.A1_N(_07188_),
    .A2_N(_07346_),
    .B1(_07441_),
    .B2(_07445_),
    .Y(_07451_));
 sky130_fd_sc_hd__a31oi_1 _17656_ (.A1(_06803_),
    .A2(_07117_),
    .A3(_07118_),
    .B1(_07115_),
    .Y(_07452_));
 sky130_fd_sc_hd__a31o_1 _17657_ (.A1(_06803_),
    .A2(_07117_),
    .A3(_07118_),
    .B1(_07115_),
    .X(_07453_));
 sky130_fd_sc_hd__o21ai_1 _17658_ (.A1(_07096_),
    .A2(_07097_),
    .B1(_07101_),
    .Y(_07455_));
 sky130_fd_sc_hd__o22a_1 _17659_ (.A1(_06805_),
    .A2(_07099_),
    .B1(_07096_),
    .B2(_07097_),
    .X(_07456_));
 sky130_fd_sc_hd__nand2_1 _17660_ (.A(net41),
    .B(net10),
    .Y(_07457_));
 sky130_fd_sc_hd__a22oi_4 _17661_ (.A1(net40),
    .A2(net11),
    .B1(net13),
    .B2(net39),
    .Y(_07458_));
 sky130_fd_sc_hd__a22o_1 _17662_ (.A1(net40),
    .A2(net11),
    .B1(net13),
    .B2(net39),
    .X(_07459_));
 sky130_fd_sc_hd__and4_1 _17663_ (.A(net39),
    .B(net40),
    .C(net11),
    .D(net13),
    .X(_07460_));
 sky130_fd_sc_hd__nand4_4 _17664_ (.A(net39),
    .B(net40),
    .C(net11),
    .D(net13),
    .Y(_07461_));
 sky130_fd_sc_hd__o211ai_1 _17665_ (.A1(_02010_),
    .A2(_02021_),
    .B1(_07459_),
    .C1(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__o21bai_1 _17666_ (.A1(_07458_),
    .A2(_07460_),
    .B1_N(_07457_),
    .Y(_07463_));
 sky130_fd_sc_hd__a22o_1 _17667_ (.A1(net41),
    .A2(net10),
    .B1(_07459_),
    .B2(_07461_),
    .X(_07464_));
 sky130_fd_sc_hd__and4_1 _17668_ (.A(_07459_),
    .B(_07461_),
    .C(net41),
    .D(net10),
    .X(_07465_));
 sky130_fd_sc_hd__nand4_1 _17669_ (.A(_07459_),
    .B(_07461_),
    .C(net41),
    .D(net10),
    .Y(_07466_));
 sky130_fd_sc_hd__nand3_2 _17670_ (.A(_07456_),
    .B(_07462_),
    .C(_07463_),
    .Y(_07467_));
 sky130_fd_sc_hd__nand2_1 _17671_ (.A(_07464_),
    .B(_07455_),
    .Y(_07468_));
 sky130_fd_sc_hd__nand3_1 _17672_ (.A(_07464_),
    .B(_07466_),
    .C(_07455_),
    .Y(_07469_));
 sky130_fd_sc_hd__o21a_1 _17673_ (.A1(_01999_),
    .A2(_02010_),
    .B1(_07252_),
    .X(_07470_));
 sky130_fd_sc_hd__a31o_1 _17674_ (.A1(_07250_),
    .A2(net41),
    .A3(net9),
    .B1(_07251_),
    .X(_07471_));
 sky130_fd_sc_hd__o2bb2ai_2 _17675_ (.A1_N(_07467_),
    .A2_N(_07469_),
    .B1(_07470_),
    .B2(_07249_),
    .Y(_07472_));
 sky130_fd_sc_hd__nand3_2 _17676_ (.A(_07467_),
    .B(_07469_),
    .C(_07471_),
    .Y(_07473_));
 sky130_fd_sc_hd__o21ai_1 _17677_ (.A1(_07243_),
    .A2(_07260_),
    .B1(_07259_),
    .Y(_07474_));
 sky130_fd_sc_hd__a21oi_1 _17678_ (.A1(_07472_),
    .A2(_07473_),
    .B1(_07474_),
    .Y(_07476_));
 sky130_fd_sc_hd__a21o_1 _17679_ (.A1(_07472_),
    .A2(_07473_),
    .B1(_07474_),
    .X(_07477_));
 sky130_fd_sc_hd__o211a_1 _17680_ (.A1(_07258_),
    .A2(_07262_),
    .B1(_07472_),
    .C1(_07473_),
    .X(_07478_));
 sky130_fd_sc_hd__o211ai_2 _17681_ (.A1(_07258_),
    .A2(_07262_),
    .B1(_07472_),
    .C1(_07473_),
    .Y(_07479_));
 sky130_fd_sc_hd__o21a_2 _17682_ (.A1(_07209_),
    .A2(_07210_),
    .B1(_07214_),
    .X(_07480_));
 sky130_fd_sc_hd__and2_1 _17683_ (.A(net7),
    .B(net45),
    .X(_07481_));
 sky130_fd_sc_hd__nand2_2 _17684_ (.A(net9),
    .B(net42),
    .Y(_07482_));
 sky130_fd_sc_hd__and4_1 _17685_ (.A(net8),
    .B(net9),
    .C(net42),
    .D(net43),
    .X(_07483_));
 sky130_fd_sc_hd__nand4_2 _17686_ (.A(net8),
    .B(net9),
    .C(net42),
    .D(net43),
    .Y(_07484_));
 sky130_fd_sc_hd__a22oi_1 _17687_ (.A1(net9),
    .A2(net42),
    .B1(net43),
    .B2(net8),
    .Y(_07485_));
 sky130_fd_sc_hd__a22o_4 _17688_ (.A1(net9),
    .A2(net42),
    .B1(net43),
    .B2(net8),
    .X(_07487_));
 sky130_fd_sc_hd__o211ai_4 _17689_ (.A1(_01977_),
    .A2(_02054_),
    .B1(_07484_),
    .C1(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__o21ai_2 _17690_ (.A1(_07483_),
    .A2(_07485_),
    .B1(_07481_),
    .Y(_07489_));
 sky130_fd_sc_hd__a22o_1 _17691_ (.A1(net7),
    .A2(net45),
    .B1(_07484_),
    .B2(_07487_),
    .X(_07490_));
 sky130_fd_sc_hd__nand4_1 _17692_ (.A(_07487_),
    .B(net45),
    .C(net7),
    .D(_07484_),
    .Y(_07491_));
 sky130_fd_sc_hd__nand3_1 _17693_ (.A(_07480_),
    .B(_07488_),
    .C(_07489_),
    .Y(_07492_));
 sky130_fd_sc_hd__a21oi_2 _17694_ (.A1(_07488_),
    .A2(_07489_),
    .B1(_07480_),
    .Y(_07493_));
 sky130_fd_sc_hd__nand3b_1 _17695_ (.A_N(_07480_),
    .B(_07490_),
    .C(_07491_),
    .Y(_07494_));
 sky130_fd_sc_hd__and2_1 _17696_ (.A(net4),
    .B(net48),
    .X(_07495_));
 sky130_fd_sc_hd__nand2_1 _17697_ (.A(net4),
    .B(net48),
    .Y(_07496_));
 sky130_fd_sc_hd__nand2_1 _17698_ (.A(net6),
    .B(net47),
    .Y(_07498_));
 sky130_fd_sc_hd__nand4_4 _17699_ (.A(net5),
    .B(net6),
    .C(net46),
    .D(net47),
    .Y(_07499_));
 sky130_fd_sc_hd__a22o_2 _17700_ (.A1(net6),
    .A2(net46),
    .B1(net47),
    .B2(net5),
    .X(_07500_));
 sky130_fd_sc_hd__and3_1 _17701_ (.A(_07496_),
    .B(_07499_),
    .C(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__o211ai_4 _17702_ (.A1(_01945_),
    .A2(_02109_),
    .B1(_07499_),
    .C1(_07500_),
    .Y(_07502_));
 sky130_fd_sc_hd__a21oi_1 _17703_ (.A1(_07499_),
    .A2(_07500_),
    .B1(_07496_),
    .Y(_07503_));
 sky130_fd_sc_hd__a21o_1 _17704_ (.A1(_07499_),
    .A2(_07500_),
    .B1(_07496_),
    .X(_07504_));
 sky130_fd_sc_hd__nand2_1 _17705_ (.A(_07502_),
    .B(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__o2bb2ai_1 _17706_ (.A1_N(_07492_),
    .A2_N(_07494_),
    .B1(_07501_),
    .B2(_07503_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand4_1 _17707_ (.A(_07492_),
    .B(_07494_),
    .C(_07502_),
    .D(_07504_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand2_1 _17708_ (.A(_07506_),
    .B(_07507_),
    .Y(_07509_));
 sky130_fd_sc_hd__o21bai_1 _17709_ (.A1(_07476_),
    .A2(_07478_),
    .B1_N(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand3_1 _17710_ (.A(_07477_),
    .B(_07479_),
    .C(_07509_),
    .Y(_07511_));
 sky130_fd_sc_hd__nand4_2 _17711_ (.A(_07477_),
    .B(_07479_),
    .C(_07506_),
    .D(_07507_),
    .Y(_07512_));
 sky130_fd_sc_hd__o21ai_1 _17712_ (.A1(_07476_),
    .A2(_07478_),
    .B1(_07509_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand2_1 _17713_ (.A(_07510_),
    .B(_07511_),
    .Y(_07514_));
 sky130_fd_sc_hd__nand3_2 _17714_ (.A(_07453_),
    .B(_07512_),
    .C(_07513_),
    .Y(_07515_));
 sky130_fd_sc_hd__a22oi_2 _17715_ (.A1(_07117_),
    .A2(_07123_),
    .B1(_07512_),
    .B2(_07513_),
    .Y(_07516_));
 sky130_fd_sc_hd__nand3_2 _17716_ (.A(_07510_),
    .B(_07511_),
    .C(_07452_),
    .Y(_07517_));
 sky130_fd_sc_hd__o21ai_4 _17717_ (.A1(_07239_),
    .A2(_07270_),
    .B1(_07269_),
    .Y(_07518_));
 sky130_fd_sc_hd__a21oi_4 _17718_ (.A1(_07515_),
    .A2(_07517_),
    .B1(_07518_),
    .Y(_07520_));
 sky130_fd_sc_hd__a21o_1 _17719_ (.A1(_07515_),
    .A2(_07517_),
    .B1(_07518_),
    .X(_07521_));
 sky130_fd_sc_hd__nand2_1 _17720_ (.A(_07515_),
    .B(_07518_),
    .Y(_07522_));
 sky130_fd_sc_hd__and3_2 _17721_ (.A(_07515_),
    .B(_07517_),
    .C(_07518_),
    .X(_07523_));
 sky130_fd_sc_hd__nor2_1 _17722_ (.A(_07520_),
    .B(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__o21ai_2 _17723_ (.A1(_07448_),
    .A2(_07450_),
    .B1(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__o211ai_4 _17724_ (.A1(_07520_),
    .A2(_07523_),
    .B1(_07449_),
    .C1(_07451_),
    .Y(_07526_));
 sky130_fd_sc_hd__o2bb2ai_2 _17725_ (.A1_N(_07449_),
    .A2_N(_07451_),
    .B1(_07520_),
    .B2(_07523_),
    .Y(_07527_));
 sky130_fd_sc_hd__o211ai_2 _17726_ (.A1(_07516_),
    .A2(_07522_),
    .B1(_07521_),
    .C1(_07449_),
    .Y(_07528_));
 sky130_fd_sc_hd__a22oi_4 _17727_ (.A1(_07195_),
    .A2(_07199_),
    .B1(_07286_),
    .B2(_07203_),
    .Y(_07529_));
 sky130_fd_sc_hd__o221a_2 _17728_ (.A1(_07450_),
    .A2(_07528_),
    .B1(_07200_),
    .B2(_07291_),
    .C1(_07527_),
    .X(_07531_));
 sky130_fd_sc_hd__o221ai_4 _17729_ (.A1(_07450_),
    .A2(_07528_),
    .B1(_07200_),
    .B2(_07291_),
    .C1(_07527_),
    .Y(_07532_));
 sky130_fd_sc_hd__nand3_4 _17730_ (.A(_07525_),
    .B(_07529_),
    .C(_07526_),
    .Y(_07533_));
 sky130_fd_sc_hd__a31oi_2 _17731_ (.A1(_07272_),
    .A2(_07273_),
    .A3(_07207_),
    .B1(_07204_),
    .Y(_07534_));
 sky130_fd_sc_hd__o21ai_2 _17732_ (.A1(_07205_),
    .A2(_07277_),
    .B1(_07276_),
    .Y(_07535_));
 sky130_fd_sc_hd__o21ai_2 _17733_ (.A1(_06980_),
    .A2(_06997_),
    .B1(_07000_),
    .Y(_07536_));
 sky130_fd_sc_hd__nand2_1 _17734_ (.A(net31),
    .B(net53),
    .Y(_07537_));
 sky130_fd_sc_hd__and4_1 _17735_ (.A(net30),
    .B(net31),
    .C(net52),
    .D(net53),
    .X(_07538_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(net31),
    .B(net52),
    .Y(_07539_));
 sky130_fd_sc_hd__a22o_1 _17737_ (.A1(net31),
    .A2(net52),
    .B1(net53),
    .B2(net30),
    .X(_07540_));
 sky130_fd_sc_hd__o2bb2ai_1 _17738_ (.A1_N(_06986_),
    .A2_N(_07539_),
    .B1(_07537_),
    .B2(_06987_),
    .Y(_07542_));
 sky130_fd_sc_hd__o21ai_1 _17739_ (.A1(_01857_),
    .A2(_02207_),
    .B1(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__o2111a_1 _17740_ (.A1(_06987_),
    .A2(_07537_),
    .B1(net29),
    .C1(net54),
    .D1(_07540_),
    .X(_07544_));
 sky130_fd_sc_hd__o2111ai_2 _17741_ (.A1(_06987_),
    .A2(_07537_),
    .B1(net29),
    .C1(net54),
    .D1(_07540_),
    .Y(_07545_));
 sky130_fd_sc_hd__o22ai_2 _17742_ (.A1(_06612_),
    .A2(_06986_),
    .B1(_06985_),
    .B2(_06989_),
    .Y(_07546_));
 sky130_fd_sc_hd__a21o_1 _17743_ (.A1(_07543_),
    .A2(_07545_),
    .B1(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__nand2_1 _17744_ (.A(_07543_),
    .B(_07546_),
    .Y(_07548_));
 sky130_fd_sc_hd__nand3_2 _17745_ (.A(_07543_),
    .B(_07545_),
    .C(_07546_),
    .Y(_07549_));
 sky130_fd_sc_hd__nand2_1 _17746_ (.A(net28),
    .B(net56),
    .Y(_07550_));
 sky130_fd_sc_hd__nand2_1 _17747_ (.A(_01769_),
    .B(net57),
    .Y(_07551_));
 sky130_fd_sc_hd__and4_1 _17748_ (.A(_01769_),
    .B(net56),
    .C(net57),
    .D(net28),
    .X(_07553_));
 sky130_fd_sc_hd__o22a_1 _17749_ (.A1(net27),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01748_),
    .X(_07554_));
 sky130_fd_sc_hd__nor2_2 _17750_ (.A(_07553_),
    .B(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__a21oi_1 _17751_ (.A1(_07547_),
    .A2(_07549_),
    .B1(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__a21o_1 _17752_ (.A1(_07547_),
    .A2(_07549_),
    .B1(_07555_),
    .X(_07557_));
 sky130_fd_sc_hd__and3_1 _17753_ (.A(_07547_),
    .B(_07549_),
    .C(_07555_),
    .X(_07558_));
 sky130_fd_sc_hd__o211ai_4 _17754_ (.A1(_07544_),
    .A2(_07548_),
    .B1(_07555_),
    .C1(_07547_),
    .Y(_07559_));
 sky130_fd_sc_hd__nand2_1 _17755_ (.A(_07557_),
    .B(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__nand3_2 _17756_ (.A(_07536_),
    .B(_07557_),
    .C(_07559_),
    .Y(_07561_));
 sky130_fd_sc_hd__o21bai_2 _17757_ (.A1(_07556_),
    .A2(_07558_),
    .B1_N(_07536_),
    .Y(_07562_));
 sky130_fd_sc_hd__a21oi_1 _17758_ (.A1(_07000_),
    .A2(_07560_),
    .B1(_06979_),
    .Y(_07564_));
 sky130_fd_sc_hd__nand3_2 _17759_ (.A(_07562_),
    .B(_06978_),
    .C(_07561_),
    .Y(_07565_));
 sky130_fd_sc_hd__a21oi_1 _17760_ (.A1(_07561_),
    .A2(_07562_),
    .B1(_06978_),
    .Y(_07566_));
 sky130_fd_sc_hd__o2bb2ai_2 _17761_ (.A1_N(_07561_),
    .A2_N(_07562_),
    .B1(_02240_),
    .B2(_06977_),
    .Y(_07567_));
 sky130_fd_sc_hd__a21oi_1 _17762_ (.A1(_07561_),
    .A2(_07564_),
    .B1(_07566_),
    .Y(_07568_));
 sky130_fd_sc_hd__nand2_1 _17763_ (.A(_07565_),
    .B(_07567_),
    .Y(_07569_));
 sky130_fd_sc_hd__o21ai_2 _17764_ (.A1(_07222_),
    .A2(_07225_),
    .B1(_07223_),
    .Y(_07570_));
 sky130_fd_sc_hd__nand2_1 _17765_ (.A(net32),
    .B(net51),
    .Y(_07571_));
 sky130_fd_sc_hd__a22oi_4 _17766_ (.A1(net3),
    .A2(net49),
    .B1(net50),
    .B2(net2),
    .Y(_07572_));
 sky130_fd_sc_hd__a22o_1 _17767_ (.A1(net3),
    .A2(net49),
    .B1(net50),
    .B2(net2),
    .X(_07573_));
 sky130_fd_sc_hd__and4_1 _17768_ (.A(net2),
    .B(net3),
    .C(net49),
    .D(net50),
    .X(_07575_));
 sky130_fd_sc_hd__nand4_4 _17769_ (.A(net2),
    .B(net3),
    .C(net49),
    .D(net50),
    .Y(_07576_));
 sky130_fd_sc_hd__o211ai_2 _17770_ (.A1(_01912_),
    .A2(_02152_),
    .B1(_07573_),
    .C1(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__o21bai_2 _17771_ (.A1(_07572_),
    .A2(_07575_),
    .B1_N(_07571_),
    .Y(_07578_));
 sky130_fd_sc_hd__a22o_1 _17772_ (.A1(net32),
    .A2(net51),
    .B1(_07573_),
    .B2(_07576_),
    .X(_07579_));
 sky130_fd_sc_hd__nand4_2 _17773_ (.A(_07573_),
    .B(_07576_),
    .C(net32),
    .D(net51),
    .Y(_07580_));
 sky130_fd_sc_hd__nand3b_4 _17774_ (.A_N(_07570_),
    .B(_07577_),
    .C(_07578_),
    .Y(_07581_));
 sky130_fd_sc_hd__and3_1 _17775_ (.A(_07579_),
    .B(_07580_),
    .C(_07570_),
    .X(_07582_));
 sky130_fd_sc_hd__nand3_4 _17776_ (.A(_07579_),
    .B(_07580_),
    .C(_07570_),
    .Y(_07583_));
 sky130_fd_sc_hd__o21a_1 _17777_ (.A1(_01879_),
    .A2(_02152_),
    .B1(_07032_),
    .X(_07584_));
 sky130_fd_sc_hd__and3_1 _17778_ (.A(_07030_),
    .B(net51),
    .C(net31),
    .X(_07586_));
 sky130_fd_sc_hd__a31o_1 _17779_ (.A1(_07030_),
    .A2(net51),
    .A3(net31),
    .B1(_07031_),
    .X(_07587_));
 sky130_fd_sc_hd__o2bb2ai_1 _17780_ (.A1_N(_07581_),
    .A2_N(_07583_),
    .B1(_07584_),
    .B2(_07029_),
    .Y(_07588_));
 sky130_fd_sc_hd__o21ai_4 _17781_ (.A1(_07031_),
    .A2(_07586_),
    .B1(_07581_),
    .Y(_07589_));
 sky130_fd_sc_hd__o2bb2ai_2 _17782_ (.A1_N(_07581_),
    .A2_N(_07583_),
    .B1(_07586_),
    .B2(_07031_),
    .Y(_07590_));
 sky130_fd_sc_hd__o2111ai_4 _17783_ (.A1(_07028_),
    .A2(_07029_),
    .B1(_07032_),
    .C1(_07581_),
    .D1(_07583_),
    .Y(_07591_));
 sky130_fd_sc_hd__a2bb2oi_2 _17784_ (.A1_N(_07219_),
    .A2_N(_07217_),
    .B1(_07218_),
    .B2(_07232_),
    .Y(_07592_));
 sky130_fd_sc_hd__o2bb2ai_2 _17785_ (.A1_N(_07218_),
    .A2_N(_07232_),
    .B1(_07219_),
    .B2(_07217_),
    .Y(_07593_));
 sky130_fd_sc_hd__nand3_4 _17786_ (.A(_07590_),
    .B(_07592_),
    .C(_07591_),
    .Y(_07594_));
 sky130_fd_sc_hd__a21oi_1 _17787_ (.A1(_07590_),
    .A2(_07591_),
    .B1(_07592_),
    .Y(_07595_));
 sky130_fd_sc_hd__o211ai_4 _17788_ (.A1(_07582_),
    .A2(_07589_),
    .B1(_07593_),
    .C1(_07588_),
    .Y(_07597_));
 sky130_fd_sc_hd__o311a_1 _17789_ (.A1(_01868_),
    .A2(_02152_),
    .A3(_06657_),
    .B1(_06660_),
    .C1(_07039_),
    .X(_07598_));
 sky130_fd_sc_hd__o31a_1 _17790_ (.A1(_06659_),
    .A2(_07024_),
    .A3(_07038_),
    .B1(_07041_),
    .X(_07599_));
 sky130_fd_sc_hd__o2bb2ai_4 _17791_ (.A1_N(_07594_),
    .A2_N(_07597_),
    .B1(_07598_),
    .B2(_07040_),
    .Y(_07600_));
 sky130_fd_sc_hd__nand3_4 _17792_ (.A(_07594_),
    .B(_07597_),
    .C(_07599_),
    .Y(_07601_));
 sky130_fd_sc_hd__a32oi_4 _17793_ (.A1(_07021_),
    .A2(_07044_),
    .A3(_07045_),
    .B1(_07047_),
    .B2(_07020_),
    .Y(_07602_));
 sky130_fd_sc_hd__a21oi_4 _17794_ (.A1(_07600_),
    .A2(_07601_),
    .B1(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__a21o_1 _17795_ (.A1(_07600_),
    .A2(_07601_),
    .B1(_07602_),
    .X(_07604_));
 sky130_fd_sc_hd__o211a_2 _17796_ (.A1(_07046_),
    .A2(_07051_),
    .B1(_07600_),
    .C1(_07601_),
    .X(_07605_));
 sky130_fd_sc_hd__o211ai_4 _17797_ (.A1(_07046_),
    .A2(_07051_),
    .B1(_07600_),
    .C1(_07601_),
    .Y(_07606_));
 sky130_fd_sc_hd__nand3_1 _17798_ (.A(_07569_),
    .B(_07604_),
    .C(_07606_),
    .Y(_07608_));
 sky130_fd_sc_hd__o21ai_2 _17799_ (.A1(_07603_),
    .A2(_07605_),
    .B1(_07568_),
    .Y(_07609_));
 sky130_fd_sc_hd__nand4_4 _17800_ (.A(_07565_),
    .B(_07567_),
    .C(_07604_),
    .D(_07606_),
    .Y(_07610_));
 sky130_fd_sc_hd__o21ai_2 _17801_ (.A1(_07603_),
    .A2(_07605_),
    .B1(_07569_),
    .Y(_07611_));
 sky130_fd_sc_hd__and3_1 _17802_ (.A(_07535_),
    .B(_07610_),
    .C(_07611_),
    .X(_07612_));
 sky130_fd_sc_hd__nand3_4 _17803_ (.A(_07535_),
    .B(_07610_),
    .C(_07611_),
    .Y(_07613_));
 sky130_fd_sc_hd__o211ai_4 _17804_ (.A1(_07277_),
    .A2(_07534_),
    .B1(_07608_),
    .C1(_07609_),
    .Y(_07614_));
 sky130_fd_sc_hd__a31o_1 _17805_ (.A1(_07017_),
    .A2(_07052_),
    .A3(_07053_),
    .B1(_07061_),
    .X(_07615_));
 sky130_fd_sc_hd__and4_1 _17806_ (.A(_07057_),
    .B(_07062_),
    .C(_07613_),
    .D(_07614_),
    .X(_07616_));
 sky130_fd_sc_hd__nand4_2 _17807_ (.A(_07057_),
    .B(_07062_),
    .C(_07613_),
    .D(_07614_),
    .Y(_07617_));
 sky130_fd_sc_hd__a22oi_2 _17808_ (.A1(_07057_),
    .A2(_07062_),
    .B1(_07613_),
    .B2(_07614_),
    .Y(_07619_));
 sky130_fd_sc_hd__a22o_1 _17809_ (.A1(_07057_),
    .A2(_07062_),
    .B1(_07613_),
    .B2(_07614_),
    .X(_07620_));
 sky130_fd_sc_hd__a21oi_4 _17810_ (.A1(_07613_),
    .A2(_07614_),
    .B1(_07615_),
    .Y(_07621_));
 sky130_fd_sc_hd__o21a_1 _17811_ (.A1(_07056_),
    .A2(_07061_),
    .B1(_07614_),
    .X(_07622_));
 sky130_fd_sc_hd__and3_1 _17812_ (.A(_07613_),
    .B(_07614_),
    .C(_07615_),
    .X(_07623_));
 sky130_fd_sc_hd__a21oi_2 _17813_ (.A1(_07622_),
    .A2(_07613_),
    .B1(_07621_),
    .Y(_07624_));
 sky130_fd_sc_hd__a32oi_2 _17814_ (.A1(_07525_),
    .A2(_07529_),
    .A3(_07526_),
    .B1(_07620_),
    .B2(_07617_),
    .Y(_07625_));
 sky130_fd_sc_hd__a32o_1 _17815_ (.A1(_07525_),
    .A2(_07529_),
    .A3(_07526_),
    .B1(_07620_),
    .B2(_07617_),
    .X(_07626_));
 sky130_fd_sc_hd__nand3_2 _17816_ (.A(_07532_),
    .B(_07533_),
    .C(_07624_),
    .Y(_07627_));
 sky130_fd_sc_hd__o2bb2ai_2 _17817_ (.A1_N(_07532_),
    .A2_N(_07533_),
    .B1(_07621_),
    .B2(_07623_),
    .Y(_07628_));
 sky130_fd_sc_hd__o2bb2ai_4 _17818_ (.A1_N(_07532_),
    .A2_N(_07533_),
    .B1(_07616_),
    .B2(_07619_),
    .Y(_07630_));
 sky130_fd_sc_hd__o211ai_4 _17819_ (.A1(_07621_),
    .A2(_07623_),
    .B1(_07532_),
    .C1(_07533_),
    .Y(_07631_));
 sky130_fd_sc_hd__a22oi_1 _17820_ (.A1(_07302_),
    .A2(_07305_),
    .B1(_07630_),
    .B2(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__nand3_4 _17821_ (.A(_07345_),
    .B(_07627_),
    .C(_07628_),
    .Y(_07633_));
 sky130_fd_sc_hd__a21oi_2 _17822_ (.A1(_07627_),
    .A2(_07628_),
    .B1(_07345_),
    .Y(_07634_));
 sky130_fd_sc_hd__nand3_4 _17823_ (.A(_07343_),
    .B(_07630_),
    .C(_07631_),
    .Y(_07635_));
 sky130_fd_sc_hd__o31a_1 _17824_ (.A1(_07063_),
    .A2(_07064_),
    .A3(_06974_),
    .B1(_06970_),
    .X(_07636_));
 sky130_fd_sc_hd__a31o_2 _17825_ (.A1(_06779_),
    .A2(_06782_),
    .A3(_07066_),
    .B1(_07636_),
    .X(_07637_));
 sky130_fd_sc_hd__o2bb2ai_2 _17826_ (.A1_N(_07633_),
    .A2_N(_07635_),
    .B1(_07636_),
    .B2(_07069_),
    .Y(_07638_));
 sky130_fd_sc_hd__o211ai_4 _17827_ (.A1(_07067_),
    .A2(_07074_),
    .B1(_07633_),
    .C1(_07635_),
    .Y(_07639_));
 sky130_fd_sc_hd__o22ai_2 _17828_ (.A1(_07067_),
    .A2(_07074_),
    .B1(_07632_),
    .B2(_07634_),
    .Y(_07641_));
 sky130_fd_sc_hd__o2111ai_4 _17829_ (.A1(_07069_),
    .A2(_06970_),
    .B1(_07068_),
    .C1(_07633_),
    .D1(_07635_),
    .Y(_07642_));
 sky130_fd_sc_hd__a22oi_4 _17830_ (.A1(_07311_),
    .A2(_07313_),
    .B1(_07638_),
    .B2(_07639_),
    .Y(_07643_));
 sky130_fd_sc_hd__nand4_4 _17831_ (.A(_07309_),
    .B(_07314_),
    .C(_07641_),
    .D(_07642_),
    .Y(_07644_));
 sky130_fd_sc_hd__a21oi_1 _17832_ (.A1(_07641_),
    .A2(_07642_),
    .B1(_07316_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand4_2 _17833_ (.A(_07311_),
    .B(_07313_),
    .C(_07638_),
    .D(_07639_),
    .Y(_07646_));
 sky130_fd_sc_hd__o21ai_1 _17834_ (.A1(_06628_),
    .A2(_07007_),
    .B1(_07008_),
    .Y(_07647_));
 sky130_fd_sc_hd__o22ai_2 _17835_ (.A1(_07007_),
    .A2(_07009_),
    .B1(_07643_),
    .B2(_07645_),
    .Y(_07648_));
 sky130_fd_sc_hd__nand3_1 _17836_ (.A(_07644_),
    .B(_07646_),
    .C(_07647_),
    .Y(_07649_));
 sky130_fd_sc_hd__o21ai_1 _17837_ (.A1(_07643_),
    .A2(_07645_),
    .B1(_07647_),
    .Y(_07650_));
 sky130_fd_sc_hd__o2111ai_1 _17838_ (.A1(_06628_),
    .A2(_07007_),
    .B1(_07008_),
    .C1(_07644_),
    .D1(_07646_),
    .Y(_07652_));
 sky130_fd_sc_hd__a21oi_1 _17839_ (.A1(_07320_),
    .A2(_07326_),
    .B1(_07322_),
    .Y(_07653_));
 sky130_fd_sc_hd__o2bb2ai_1 _17840_ (.A1_N(_07320_),
    .A2_N(_07326_),
    .B1(_07321_),
    .B2(_07315_),
    .Y(_07654_));
 sky130_fd_sc_hd__a21oi_1 _17841_ (.A1(_07648_),
    .A2(_07649_),
    .B1(_07654_),
    .Y(_07655_));
 sky130_fd_sc_hd__nand3_1 _17842_ (.A(_07653_),
    .B(_07652_),
    .C(_07650_),
    .Y(_07656_));
 sky130_fd_sc_hd__o211a_1 _17843_ (.A1(_07322_),
    .A2(_07330_),
    .B1(_07648_),
    .C1(_07649_),
    .X(_07657_));
 sky130_fd_sc_hd__o211ai_1 _17844_ (.A1(_07322_),
    .A2(_07330_),
    .B1(_07648_),
    .C1(_07649_),
    .Y(_07658_));
 sky130_fd_sc_hd__nor2_1 _17845_ (.A(_07655_),
    .B(_07657_),
    .Y(_07659_));
 sky130_fd_sc_hd__a2bb2o_1 _17846_ (.A1_N(_07339_),
    .A2_N(_07342_),
    .B1(_07332_),
    .B2(_07336_),
    .X(_07660_));
 sky130_fd_sc_hd__xor2_1 _17847_ (.A(_07659_),
    .B(_07660_),
    .X(net93));
 sky130_fd_sc_hd__a32oi_4 _17848_ (.A1(_07343_),
    .A2(_07630_),
    .A3(_07631_),
    .B1(_07633_),
    .B2(_07637_),
    .Y(_07662_));
 sky130_fd_sc_hd__a31o_1 _17849_ (.A1(_07535_),
    .A2(_07610_),
    .A3(_07611_),
    .B1(_07615_),
    .X(_07663_));
 sky130_fd_sc_hd__a31o_1 _17850_ (.A1(_07535_),
    .A2(_07610_),
    .A3(_07611_),
    .B1(_07622_),
    .X(_07664_));
 sky130_fd_sc_hd__inv_2 _17851_ (.A(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__o21ai_1 _17852_ (.A1(_07621_),
    .A2(_07623_),
    .B1(_07532_),
    .Y(_07666_));
 sky130_fd_sc_hd__o21ai_4 _17853_ (.A1(_07520_),
    .A2(_07523_),
    .B1(_07449_),
    .Y(_07667_));
 sky130_fd_sc_hd__o21ai_4 _17854_ (.A1(_07347_),
    .A2(_07447_),
    .B1(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__o21ai_2 _17855_ (.A1(_07434_),
    .A2(_07436_),
    .B1(_07444_),
    .Y(_07669_));
 sky130_fd_sc_hd__a21oi_2 _17856_ (.A1(_07424_),
    .A2(_07428_),
    .B1(_07402_),
    .Y(_07670_));
 sky130_fd_sc_hd__a31o_1 _17857_ (.A1(_07401_),
    .A2(_07424_),
    .A3(_07428_),
    .B1(_07402_),
    .X(_07671_));
 sky130_fd_sc_hd__a31oi_2 _17858_ (.A1(_07392_),
    .A2(_07394_),
    .A3(_07129_),
    .B1(_06880_),
    .Y(_07673_));
 sky130_fd_sc_hd__a31o_1 _17859_ (.A1(_07392_),
    .A2(_07394_),
    .A3(_07129_),
    .B1(_06880_),
    .X(_07674_));
 sky130_fd_sc_hd__nand2_1 _17860_ (.A(net60),
    .B(net25),
    .Y(_07675_));
 sky130_fd_sc_hd__a22oi_1 _17861_ (.A1(net60),
    .A2(net25),
    .B1(_07134_),
    .B2(_07389_),
    .Y(_07676_));
 sky130_fd_sc_hd__o2bb2ai_4 _17862_ (.A1_N(_07134_),
    .A2_N(_07389_),
    .B1(_01835_),
    .B2(_02251_),
    .Y(_07677_));
 sky130_fd_sc_hd__and3_1 _17863_ (.A(_07389_),
    .B(net60),
    .C(_07134_),
    .X(_07678_));
 sky130_fd_sc_hd__nand3_4 _17864_ (.A(_07389_),
    .B(net60),
    .C(_07134_),
    .Y(_07679_));
 sky130_fd_sc_hd__o31a_1 _17865_ (.A1(_01835_),
    .A2(_07133_),
    .A3(_07387_),
    .B1(_07677_),
    .X(_07680_));
 sky130_fd_sc_hd__a22oi_4 _17866_ (.A1(_06881_),
    .A2(_07128_),
    .B1(_07677_),
    .B2(_07679_),
    .Y(_07681_));
 sky130_fd_sc_hd__a22o_4 _17867_ (.A1(_06881_),
    .A2(_07128_),
    .B1(_07677_),
    .B2(_07679_),
    .X(_07682_));
 sky130_fd_sc_hd__o311a_1 _17868_ (.A1(_01835_),
    .A2(_07133_),
    .A3(_07387_),
    .B1(_07129_),
    .C1(_07677_),
    .X(_07684_));
 sky130_fd_sc_hd__o211ai_4 _17869_ (.A1(_01835_),
    .A2(_07390_),
    .B1(_07677_),
    .C1(_07129_),
    .Y(_07685_));
 sky130_fd_sc_hd__o21ai_4 _17870_ (.A1(_07681_),
    .A2(_07684_),
    .B1(_07673_),
    .Y(_07686_));
 sky130_fd_sc_hd__inv_2 _17871_ (.A(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__a21oi_1 _17872_ (.A1(_06881_),
    .A2(_07397_),
    .B1(_07681_),
    .Y(_07688_));
 sky130_fd_sc_hd__nand3_4 _17873_ (.A(_07674_),
    .B(_07682_),
    .C(_07685_),
    .Y(_07689_));
 sky130_fd_sc_hd__o21a_1 _17874_ (.A1(_01890_),
    .A2(_02163_),
    .B1(_07411_),
    .X(_07690_));
 sky130_fd_sc_hd__and3_1 _17875_ (.A(_07408_),
    .B(net20),
    .C(net63),
    .X(_07691_));
 sky130_fd_sc_hd__a31o_1 _17876_ (.A1(_07408_),
    .A2(net20),
    .A3(net63),
    .B1(_07409_),
    .X(_07692_));
 sky130_fd_sc_hd__o31a_1 _17877_ (.A1(_01890_),
    .A2(_02163_),
    .A3(_07407_),
    .B1(_07411_),
    .X(_07693_));
 sky130_fd_sc_hd__a31oi_4 _17878_ (.A1(net58),
    .A2(net59),
    .A3(net25),
    .B1(net24),
    .Y(_07695_));
 sky130_fd_sc_hd__a31oi_2 _17879_ (.A1(net58),
    .A2(net59),
    .A3(net25),
    .B1(net60),
    .Y(_07696_));
 sky130_fd_sc_hd__a31o_1 _17880_ (.A1(net58),
    .A2(net59),
    .A3(net25),
    .B1(net60),
    .X(_07697_));
 sky130_fd_sc_hd__a21oi_4 _17881_ (.A1(_01835_),
    .A2(_07134_),
    .B1(_07387_),
    .Y(_07698_));
 sky130_fd_sc_hd__a21o_4 _17882_ (.A1(_01835_),
    .A2(_07134_),
    .B1(_07387_),
    .X(_07699_));
 sky130_fd_sc_hd__o2111a_1 _17883_ (.A1(net58),
    .A2(net59),
    .B1(net60),
    .C1(net24),
    .D1(net25),
    .X(_07700_));
 sky130_fd_sc_hd__nand4_4 _17884_ (.A(net61),
    .B(net62),
    .C(net22),
    .D(net24),
    .Y(_07701_));
 sky130_fd_sc_hd__a22oi_4 _17885_ (.A1(net62),
    .A2(net22),
    .B1(net24),
    .B2(net61),
    .Y(_07702_));
 sky130_fd_sc_hd__a22o_1 _17886_ (.A1(net62),
    .A2(net22),
    .B1(net24),
    .B2(net61),
    .X(_07703_));
 sky130_fd_sc_hd__nand4_4 _17887_ (.A(_07703_),
    .B(net21),
    .C(net63),
    .D(_07701_),
    .Y(_07704_));
 sky130_fd_sc_hd__o2bb2ai_4 _17888_ (.A1_N(_07701_),
    .A2_N(_07703_),
    .B1(_01890_),
    .B2(_02185_),
    .Y(_07706_));
 sky130_fd_sc_hd__o211a_4 _17889_ (.A1(_07133_),
    .A2(_07700_),
    .B1(_07704_),
    .C1(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__o2111ai_4 _17890_ (.A1(net24),
    .A2(_07133_),
    .B1(_07698_),
    .C1(_07704_),
    .D1(_07706_),
    .Y(_07708_));
 sky130_fd_sc_hd__a2bb2oi_4 _17891_ (.A1_N(_07695_),
    .A2_N(_07699_),
    .B1(_07704_),
    .B2(_07706_),
    .Y(_07709_));
 sky130_fd_sc_hd__o2bb2ai_4 _17892_ (.A1_N(_07704_),
    .A2_N(_07706_),
    .B1(_07695_),
    .B2(_07699_),
    .Y(_07710_));
 sky130_fd_sc_hd__o21ai_1 _17893_ (.A1(_07707_),
    .A2(_07709_),
    .B1(_07692_),
    .Y(_07711_));
 sky130_fd_sc_hd__o2111ai_1 _17894_ (.A1(_07406_),
    .A2(_07407_),
    .B1(_07411_),
    .C1(_07708_),
    .D1(_07710_),
    .Y(_07712_));
 sky130_fd_sc_hd__o21ai_2 _17895_ (.A1(_07409_),
    .A2(_07691_),
    .B1(_07710_),
    .Y(_07713_));
 sky130_fd_sc_hd__o211ai_4 _17896_ (.A1(_07409_),
    .A2(_07691_),
    .B1(_07708_),
    .C1(_07710_),
    .Y(_07714_));
 sky130_fd_sc_hd__o22ai_4 _17897_ (.A1(_07407_),
    .A2(_07690_),
    .B1(_07707_),
    .B2(_07709_),
    .Y(_07715_));
 sky130_fd_sc_hd__a22oi_4 _17898_ (.A1(_07686_),
    .A2(_07689_),
    .B1(_07714_),
    .B2(_07715_),
    .Y(_07717_));
 sky130_fd_sc_hd__a22o_1 _17899_ (.A1(_07686_),
    .A2(_07689_),
    .B1(_07714_),
    .B2(_07715_),
    .X(_07718_));
 sky130_fd_sc_hd__o2111a_1 _17900_ (.A1(_07707_),
    .A2(_07713_),
    .B1(_07715_),
    .C1(_07689_),
    .D1(_07686_),
    .X(_07719_));
 sky130_fd_sc_hd__o2111ai_4 _17901_ (.A1(_07707_),
    .A2(_07713_),
    .B1(_07715_),
    .C1(_07689_),
    .D1(_07686_),
    .Y(_07720_));
 sky130_fd_sc_hd__nand3_4 _17902_ (.A(_07671_),
    .B(_07718_),
    .C(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__o22a_1 _17903_ (.A1(_07400_),
    .A2(_07670_),
    .B1(_07717_),
    .B2(_07719_),
    .X(_07722_));
 sky130_fd_sc_hd__o22ai_4 _17904_ (.A1(_07400_),
    .A2(_07670_),
    .B1(_07717_),
    .B2(_07719_),
    .Y(_07723_));
 sky130_fd_sc_hd__a21oi_2 _17905_ (.A1(_07416_),
    .A2(_07420_),
    .B1(_07417_),
    .Y(_07724_));
 sky130_fd_sc_hd__a31o_1 _17906_ (.A1(_07404_),
    .A2(_07414_),
    .A3(_07415_),
    .B1(_07425_),
    .X(_07725_));
 sky130_fd_sc_hd__o21ai_4 _17907_ (.A1(_07349_),
    .A2(_07350_),
    .B1(_07353_),
    .Y(_07726_));
 sky130_fd_sc_hd__nand2_1 _17908_ (.A(net35),
    .B(net18),
    .Y(_07728_));
 sky130_fd_sc_hd__and4_1 _17909_ (.A(net64),
    .B(net34),
    .C(net19),
    .D(net20),
    .X(_07729_));
 sky130_fd_sc_hd__nand4_4 _17910_ (.A(net64),
    .B(net34),
    .C(net19),
    .D(net20),
    .Y(_07730_));
 sky130_fd_sc_hd__a22oi_2 _17911_ (.A1(net34),
    .A2(net19),
    .B1(net20),
    .B2(net64),
    .Y(_07731_));
 sky130_fd_sc_hd__a22o_1 _17912_ (.A1(net34),
    .A2(net19),
    .B1(net20),
    .B2(net64),
    .X(_07732_));
 sky130_fd_sc_hd__o211ai_2 _17913_ (.A1(_01934_),
    .A2(_02131_),
    .B1(_07730_),
    .C1(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__o21bai_2 _17914_ (.A1(_07729_),
    .A2(_07731_),
    .B1_N(_07728_),
    .Y(_07734_));
 sky130_fd_sc_hd__a22o_2 _17915_ (.A1(net35),
    .A2(net18),
    .B1(_07730_),
    .B2(_07732_),
    .X(_07735_));
 sky130_fd_sc_hd__nand4_4 _17916_ (.A(_07732_),
    .B(net18),
    .C(net35),
    .D(_07730_),
    .Y(_07736_));
 sky130_fd_sc_hd__nand3b_4 _17917_ (.A_N(_07726_),
    .B(_07733_),
    .C(_07734_),
    .Y(_07737_));
 sky130_fd_sc_hd__nand3_4 _17918_ (.A(_07735_),
    .B(_07736_),
    .C(_07726_),
    .Y(_07739_));
 sky130_fd_sc_hd__nand2_1 _17919_ (.A(net38),
    .B(net15),
    .Y(_07740_));
 sky130_fd_sc_hd__nand2_1 _17920_ (.A(net36),
    .B(net17),
    .Y(_07741_));
 sky130_fd_sc_hd__a22oi_4 _17921_ (.A1(net37),
    .A2(net16),
    .B1(net17),
    .B2(net36),
    .Y(_07742_));
 sky130_fd_sc_hd__nand2_1 _17922_ (.A(net37),
    .B(net17),
    .Y(_07743_));
 sky130_fd_sc_hd__and4_2 _17923_ (.A(net36),
    .B(net37),
    .C(net16),
    .D(net17),
    .X(_07744_));
 sky130_fd_sc_hd__o2bb2a_1 _17924_ (.A1_N(net38),
    .A2_N(net15),
    .B1(_07742_),
    .B2(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__o21ai_2 _17925_ (.A1(_07742_),
    .A2(_07744_),
    .B1(_07740_),
    .Y(_07746_));
 sky130_fd_sc_hd__a41o_1 _17926_ (.A1(net36),
    .A2(net37),
    .A3(net16),
    .A4(net17),
    .B1(_07740_),
    .X(_07747_));
 sky130_fd_sc_hd__nor2_1 _17927_ (.A(_07742_),
    .B(_07747_),
    .Y(_07748_));
 sky130_fd_sc_hd__o21ai_1 _17928_ (.A1(_07742_),
    .A2(_07747_),
    .B1(_07746_),
    .Y(_07750_));
 sky130_fd_sc_hd__o21a_1 _17929_ (.A1(_07742_),
    .A2(_07747_),
    .B1(_07746_),
    .X(_07751_));
 sky130_fd_sc_hd__o2111ai_4 _17930_ (.A1(_07742_),
    .A2(_07747_),
    .B1(_07746_),
    .C1(_07737_),
    .D1(_07739_),
    .Y(_07752_));
 sky130_fd_sc_hd__a21o_1 _17931_ (.A1(_07737_),
    .A2(_07739_),
    .B1(_07751_),
    .X(_07753_));
 sky130_fd_sc_hd__o211ai_4 _17932_ (.A1(_07745_),
    .A2(_07748_),
    .B1(_07737_),
    .C1(_07739_),
    .Y(_07754_));
 sky130_fd_sc_hd__a21o_1 _17933_ (.A1(_07737_),
    .A2(_07739_),
    .B1(_07750_),
    .X(_07755_));
 sky130_fd_sc_hd__and3_2 _17934_ (.A(_07755_),
    .B(_07724_),
    .C(_07754_),
    .X(_07756_));
 sky130_fd_sc_hd__nand3_2 _17935_ (.A(_07755_),
    .B(_07724_),
    .C(_07754_),
    .Y(_07757_));
 sky130_fd_sc_hd__o211ai_4 _17936_ (.A1(_07417_),
    .A2(_07425_),
    .B1(_07752_),
    .C1(_07753_),
    .Y(_07758_));
 sky130_fd_sc_hd__a32oi_4 _17937_ (.A1(_07348_),
    .A2(_07357_),
    .A3(_07358_),
    .B1(_07359_),
    .B2(_07370_),
    .Y(_07759_));
 sky130_fd_sc_hd__a32o_1 _17938_ (.A1(_07348_),
    .A2(_07357_),
    .A3(_07358_),
    .B1(_07359_),
    .B2(_07370_),
    .X(_07761_));
 sky130_fd_sc_hd__a21o_1 _17939_ (.A1(_07757_),
    .A2(_07758_),
    .B1(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__nand3_1 _17940_ (.A(_07757_),
    .B(_07758_),
    .C(_07761_),
    .Y(_07763_));
 sky130_fd_sc_hd__and3_1 _17941_ (.A(_07757_),
    .B(_07758_),
    .C(_07759_),
    .X(_07764_));
 sky130_fd_sc_hd__nand4_2 _17942_ (.A(_07360_),
    .B(_07374_),
    .C(_07757_),
    .D(_07758_),
    .Y(_07765_));
 sky130_fd_sc_hd__a21oi_1 _17943_ (.A1(_07757_),
    .A2(_07758_),
    .B1(_07759_),
    .Y(_07766_));
 sky130_fd_sc_hd__a22o_1 _17944_ (.A1(_07360_),
    .A2(_07374_),
    .B1(_07757_),
    .B2(_07758_),
    .X(_07767_));
 sky130_fd_sc_hd__nand4_2 _17945_ (.A(_07721_),
    .B(_07723_),
    .C(_07765_),
    .D(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__o2bb2ai_2 _17946_ (.A1_N(_07721_),
    .A2_N(_07723_),
    .B1(_07764_),
    .B2(_07766_),
    .Y(_07769_));
 sky130_fd_sc_hd__a22o_1 _17947_ (.A1(_07721_),
    .A2(_07723_),
    .B1(_07762_),
    .B2(_07763_),
    .X(_07770_));
 sky130_fd_sc_hd__nand3_1 _17948_ (.A(_07721_),
    .B(_07762_),
    .C(_07763_),
    .Y(_07772_));
 sky130_fd_sc_hd__o2111ai_4 _17949_ (.A1(_07434_),
    .A2(_07436_),
    .B1(_07444_),
    .C1(_07768_),
    .D1(_07769_),
    .Y(_07773_));
 sky130_fd_sc_hd__a22oi_2 _17950_ (.A1(_07438_),
    .A2(_07444_),
    .B1(_07768_),
    .B2(_07769_),
    .Y(_07774_));
 sky130_fd_sc_hd__o211ai_4 _17951_ (.A1(_07772_),
    .A2(_07722_),
    .B1(_07669_),
    .C1(_07770_),
    .Y(_07775_));
 sky130_fd_sc_hd__a21boi_2 _17952_ (.A1(_07380_),
    .A2(_07382_),
    .B1_N(_07381_),
    .Y(_07776_));
 sky130_fd_sc_hd__o21ai_2 _17953_ (.A1(_07376_),
    .A2(_07379_),
    .B1(_07384_),
    .Y(_07777_));
 sky130_fd_sc_hd__a41o_2 _17954_ (.A1(net8),
    .A2(net9),
    .A3(net42),
    .A4(net43),
    .B1(_07481_),
    .X(_07778_));
 sky130_fd_sc_hd__a31o_1 _17955_ (.A1(_07487_),
    .A2(net45),
    .A3(net7),
    .B1(_07483_),
    .X(_07779_));
 sky130_fd_sc_hd__and2_1 _17956_ (.A(net8),
    .B(net45),
    .X(_07780_));
 sky130_fd_sc_hd__nand2_2 _17957_ (.A(net10),
    .B(net43),
    .Y(_07781_));
 sky130_fd_sc_hd__nand4_1 _17958_ (.A(net9),
    .B(net10),
    .C(net42),
    .D(net43),
    .Y(_07783_));
 sky130_fd_sc_hd__a22o_2 _17959_ (.A1(net10),
    .A2(net42),
    .B1(net43),
    .B2(net9),
    .X(_07784_));
 sky130_fd_sc_hd__a2bb2oi_1 _17960_ (.A1_N(_01988_),
    .A2_N(_02054_),
    .B1(_07783_),
    .B2(_07784_),
    .Y(_07785_));
 sky130_fd_sc_hd__a22o_1 _17961_ (.A1(net8),
    .A2(net45),
    .B1(_07783_),
    .B2(_07784_),
    .X(_07786_));
 sky130_fd_sc_hd__o211a_2 _17962_ (.A1(_07482_),
    .A2(_07781_),
    .B1(_07780_),
    .C1(_07784_),
    .X(_07787_));
 sky130_fd_sc_hd__o2111ai_4 _17963_ (.A1(_07482_),
    .A2(_07781_),
    .B1(net8),
    .C1(net45),
    .D1(_07784_),
    .Y(_07788_));
 sky130_fd_sc_hd__o2bb2ai_4 _17964_ (.A1_N(_07487_),
    .A2_N(_07778_),
    .B1(_07785_),
    .B2(_07787_),
    .Y(_07789_));
 sky130_fd_sc_hd__nand2_1 _17965_ (.A(_07779_),
    .B(_07786_),
    .Y(_07790_));
 sky130_fd_sc_hd__nand4_4 _17966_ (.A(_07487_),
    .B(_07778_),
    .C(_07786_),
    .D(_07788_),
    .Y(_07791_));
 sky130_fd_sc_hd__inv_2 _17967_ (.A(_07791_),
    .Y(_07792_));
 sky130_fd_sc_hd__nand2_1 _17968_ (.A(net7),
    .B(net46),
    .Y(_07794_));
 sky130_fd_sc_hd__a22oi_2 _17969_ (.A1(net7),
    .A2(net46),
    .B1(net47),
    .B2(net6),
    .Y(_07795_));
 sky130_fd_sc_hd__a22o_1 _17970_ (.A1(net7),
    .A2(net46),
    .B1(net47),
    .B2(net6),
    .X(_07796_));
 sky130_fd_sc_hd__and4_2 _17971_ (.A(net6),
    .B(net7),
    .C(net46),
    .D(net47),
    .X(_07797_));
 sky130_fd_sc_hd__nand4_2 _17972_ (.A(net6),
    .B(net7),
    .C(net46),
    .D(net47),
    .Y(_07798_));
 sky130_fd_sc_hd__nand2_1 _17973_ (.A(net5),
    .B(net48),
    .Y(_07799_));
 sky130_fd_sc_hd__a22oi_4 _17974_ (.A1(net5),
    .A2(net48),
    .B1(_07796_),
    .B2(_07798_),
    .Y(_07800_));
 sky130_fd_sc_hd__nor3_2 _17975_ (.A(_07795_),
    .B(_07799_),
    .C(_07797_),
    .Y(_07801_));
 sky130_fd_sc_hd__nor2_2 _17976_ (.A(_07800_),
    .B(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__a211oi_2 _17977_ (.A1(_07789_),
    .A2(_07791_),
    .B1(_07800_),
    .C1(_07801_),
    .Y(_07803_));
 sky130_fd_sc_hd__o221a_1 _17978_ (.A1(_07800_),
    .A2(_07801_),
    .B1(_07787_),
    .B2(_07790_),
    .C1(_07789_),
    .X(_07805_));
 sky130_fd_sc_hd__o2bb2a_2 _17979_ (.A1_N(_07789_),
    .A2_N(_07791_),
    .B1(_07800_),
    .B2(_07801_),
    .X(_07806_));
 sky130_fd_sc_hd__a21o_1 _17980_ (.A1(_07789_),
    .A2(_07791_),
    .B1(_07802_),
    .X(_07807_));
 sky130_fd_sc_hd__nand2_4 _17981_ (.A(_07789_),
    .B(_07802_),
    .Y(_07808_));
 sky130_fd_sc_hd__and3_2 _17982_ (.A(_07789_),
    .B(_07791_),
    .C(_07802_),
    .X(_07809_));
 sky130_fd_sc_hd__o21ai_2 _17983_ (.A1(_07808_),
    .A2(_07792_),
    .B1(_07807_),
    .Y(_07810_));
 sky130_fd_sc_hd__o2bb2a_1 _17984_ (.A1_N(_07471_),
    .A2_N(_07467_),
    .B1(_07465_),
    .B2(_07468_),
    .X(_07811_));
 sky130_fd_sc_hd__o2bb2ai_4 _17985_ (.A1_N(_07471_),
    .A2_N(_07467_),
    .B1(_07465_),
    .B2(_07468_),
    .Y(_07812_));
 sky130_fd_sc_hd__o21a_1 _17986_ (.A1(_02010_),
    .A2(_02021_),
    .B1(_07461_),
    .X(_07813_));
 sky130_fd_sc_hd__a31o_1 _17987_ (.A1(_07459_),
    .A2(net10),
    .A3(net41),
    .B1(_07460_),
    .X(_07814_));
 sky130_fd_sc_hd__o31a_1 _17988_ (.A1(_02010_),
    .A2(_02021_),
    .A3(_07458_),
    .B1(_07461_),
    .X(_07816_));
 sky130_fd_sc_hd__a21oi_2 _17989_ (.A1(_07099_),
    .A2(_07363_),
    .B1(_07362_),
    .Y(_07817_));
 sky130_fd_sc_hd__o21ai_4 _17990_ (.A1(_07362_),
    .A2(_07364_),
    .B1(_07367_),
    .Y(_07818_));
 sky130_fd_sc_hd__nand2_1 _17991_ (.A(net41),
    .B(net11),
    .Y(_07819_));
 sky130_fd_sc_hd__and4_1 _17992_ (.A(net39),
    .B(net40),
    .C(net13),
    .D(net14),
    .X(_07820_));
 sky130_fd_sc_hd__nand4_4 _17993_ (.A(net39),
    .B(net40),
    .C(net13),
    .D(net14),
    .Y(_07821_));
 sky130_fd_sc_hd__a22o_4 _17994_ (.A1(net40),
    .A2(net13),
    .B1(net14),
    .B2(net39),
    .X(_07822_));
 sky130_fd_sc_hd__o211a_1 _17995_ (.A1(_02010_),
    .A2(_02032_),
    .B1(_07821_),
    .C1(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__a21oi_1 _17996_ (.A1(_07821_),
    .A2(_07822_),
    .B1(_07819_),
    .Y(_07824_));
 sky130_fd_sc_hd__nand4_4 _17997_ (.A(_07822_),
    .B(net11),
    .C(net41),
    .D(_07821_),
    .Y(_07825_));
 sky130_fd_sc_hd__o2bb2ai_4 _17998_ (.A1_N(_07821_),
    .A2_N(_07822_),
    .B1(_02010_),
    .B2(_02032_),
    .Y(_07827_));
 sky130_fd_sc_hd__o211a_2 _17999_ (.A1(_07365_),
    .A2(_07817_),
    .B1(_07825_),
    .C1(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__o211ai_4 _18000_ (.A1(_07365_),
    .A2(_07817_),
    .B1(_07825_),
    .C1(_07827_),
    .Y(_07829_));
 sky130_fd_sc_hd__a21oi_4 _18001_ (.A1(_07825_),
    .A2(_07827_),
    .B1(_07818_),
    .Y(_07830_));
 sky130_fd_sc_hd__o31ai_4 _18002_ (.A1(_07818_),
    .A2(_07823_),
    .A3(_07824_),
    .B1(_07814_),
    .Y(_07831_));
 sky130_fd_sc_hd__nand3b_1 _18003_ (.A_N(_07830_),
    .B(_07814_),
    .C(_07829_),
    .Y(_07832_));
 sky130_fd_sc_hd__o22ai_4 _18004_ (.A1(_07458_),
    .A2(_07813_),
    .B1(_07828_),
    .B2(_07830_),
    .Y(_07833_));
 sky130_fd_sc_hd__o21ai_1 _18005_ (.A1(_07828_),
    .A2(_07831_),
    .B1(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__o211a_4 _18006_ (.A1(_07831_),
    .A2(_07828_),
    .B1(_07812_),
    .C1(_07833_),
    .X(_07835_));
 sky130_fd_sc_hd__o211ai_4 _18007_ (.A1(_07831_),
    .A2(_07828_),
    .B1(_07812_),
    .C1(_07833_),
    .Y(_07836_));
 sky130_fd_sc_hd__a21oi_4 _18008_ (.A1(_07832_),
    .A2(_07833_),
    .B1(_07812_),
    .Y(_07838_));
 sky130_fd_sc_hd__nand2_2 _18009_ (.A(_07834_),
    .B(_07811_),
    .Y(_07839_));
 sky130_fd_sc_hd__o211ai_4 _18010_ (.A1(_07806_),
    .A2(_07809_),
    .B1(_07836_),
    .C1(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__o22ai_4 _18011_ (.A1(_07803_),
    .A2(_07805_),
    .B1(_07835_),
    .B2(_07838_),
    .Y(_07841_));
 sky130_fd_sc_hd__o211a_1 _18012_ (.A1(_07808_),
    .A2(_07792_),
    .B1(_07807_),
    .C1(_07839_),
    .X(_07842_));
 sky130_fd_sc_hd__o2111ai_4 _18013_ (.A1(_07808_),
    .A2(_07792_),
    .B1(_07807_),
    .C1(_07836_),
    .D1(_07839_),
    .Y(_07843_));
 sky130_fd_sc_hd__o22ai_4 _18014_ (.A1(_07806_),
    .A2(_07809_),
    .B1(_07835_),
    .B2(_07838_),
    .Y(_07844_));
 sky130_fd_sc_hd__nand3_4 _18015_ (.A(_07777_),
    .B(_07843_),
    .C(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__and3_1 _18016_ (.A(_07841_),
    .B(_07776_),
    .C(_07840_),
    .X(_07846_));
 sky130_fd_sc_hd__nand3_2 _18017_ (.A(_07841_),
    .B(_07776_),
    .C(_07840_),
    .Y(_07847_));
 sky130_fd_sc_hd__a21oi_2 _18018_ (.A1(_07477_),
    .A2(_07509_),
    .B1(_07478_),
    .Y(_07849_));
 sky130_fd_sc_hd__a32o_2 _18019_ (.A1(_07472_),
    .A2(_07473_),
    .A3(_07474_),
    .B1(_07477_),
    .B2(_07509_),
    .X(_07850_));
 sky130_fd_sc_hd__and3_1 _18020_ (.A(_07845_),
    .B(_07847_),
    .C(_07849_),
    .X(_07851_));
 sky130_fd_sc_hd__a21oi_1 _18021_ (.A1(_07845_),
    .A2(_07847_),
    .B1(_07849_),
    .Y(_07852_));
 sky130_fd_sc_hd__a21oi_2 _18022_ (.A1(_07845_),
    .A2(_07847_),
    .B1(_07850_),
    .Y(_07853_));
 sky130_fd_sc_hd__a21o_1 _18023_ (.A1(_07845_),
    .A2(_07847_),
    .B1(_07850_),
    .X(_07854_));
 sky130_fd_sc_hd__and3_1 _18024_ (.A(_07845_),
    .B(_07847_),
    .C(_07850_),
    .X(_07855_));
 sky130_fd_sc_hd__nand3_2 _18025_ (.A(_07845_),
    .B(_07847_),
    .C(_07850_),
    .Y(_07856_));
 sky130_fd_sc_hd__o2bb2a_1 _18026_ (.A1_N(_07773_),
    .A2_N(_07775_),
    .B1(_07853_),
    .B2(_07855_),
    .X(_07857_));
 sky130_fd_sc_hd__o2bb2ai_2 _18027_ (.A1_N(_07773_),
    .A2_N(_07775_),
    .B1(_07853_),
    .B2(_07855_),
    .Y(_07858_));
 sky130_fd_sc_hd__nand4_4 _18028_ (.A(_07773_),
    .B(_07775_),
    .C(_07854_),
    .D(_07856_),
    .Y(_07860_));
 sky130_fd_sc_hd__o2bb2ai_2 _18029_ (.A1_N(_07773_),
    .A2_N(_07775_),
    .B1(_07851_),
    .B2(_07852_),
    .Y(_07861_));
 sky130_fd_sc_hd__o211ai_4 _18030_ (.A1(_07853_),
    .A2(_07855_),
    .B1(_07773_),
    .C1(_07775_),
    .Y(_07862_));
 sky130_fd_sc_hd__o211ai_4 _18031_ (.A1(_07448_),
    .A2(_07524_),
    .B1(_07860_),
    .C1(_07451_),
    .Y(_07863_));
 sky130_fd_sc_hd__and4_1 _18032_ (.A(_07451_),
    .B(_07667_),
    .C(_07858_),
    .D(_07860_),
    .X(_07864_));
 sky130_fd_sc_hd__nand4_4 _18033_ (.A(_07451_),
    .B(_07667_),
    .C(_07858_),
    .D(_07860_),
    .Y(_07865_));
 sky130_fd_sc_hd__nand3_4 _18034_ (.A(_07668_),
    .B(_07861_),
    .C(_07862_),
    .Y(_07866_));
 sky130_fd_sc_hd__a21oi_2 _18035_ (.A1(_07515_),
    .A2(_07518_),
    .B1(_07516_),
    .Y(_07867_));
 sky130_fd_sc_hd__o21ai_2 _18036_ (.A1(_07453_),
    .A2(_07514_),
    .B1(_07522_),
    .Y(_07868_));
 sky130_fd_sc_hd__a21oi_2 _18037_ (.A1(_07594_),
    .A2(_07599_),
    .B1(_07595_),
    .Y(_07869_));
 sky130_fd_sc_hd__a21bo_2 _18038_ (.A1(_07500_),
    .A2(_07495_),
    .B1_N(_07499_),
    .X(_07871_));
 sky130_fd_sc_hd__a21boi_1 _18039_ (.A1(_07500_),
    .A2(_07495_),
    .B1_N(_07499_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_1 _18040_ (.A(net2),
    .B(net51),
    .Y(_07873_));
 sky130_fd_sc_hd__nand4_4 _18041_ (.A(net3),
    .B(net4),
    .C(net49),
    .D(net50),
    .Y(_07874_));
 sky130_fd_sc_hd__a22oi_4 _18042_ (.A1(net4),
    .A2(net49),
    .B1(net50),
    .B2(net3),
    .Y(_07875_));
 sky130_fd_sc_hd__a22o_1 _18043_ (.A1(net4),
    .A2(net49),
    .B1(net50),
    .B2(net3),
    .X(_07876_));
 sky130_fd_sc_hd__o211ai_1 _18044_ (.A1(_01901_),
    .A2(_02152_),
    .B1(_07874_),
    .C1(_07876_),
    .Y(_07877_));
 sky130_fd_sc_hd__a21o_1 _18045_ (.A1(_07874_),
    .A2(_07876_),
    .B1(_07873_),
    .X(_07878_));
 sky130_fd_sc_hd__a22o_2 _18046_ (.A1(net2),
    .A2(net51),
    .B1(_07874_),
    .B2(_07876_),
    .X(_07879_));
 sky130_fd_sc_hd__nand4_4 _18047_ (.A(_07876_),
    .B(net51),
    .C(net2),
    .D(_07874_),
    .Y(_07880_));
 sky130_fd_sc_hd__a21oi_4 _18048_ (.A1(_07879_),
    .A2(_07880_),
    .B1(_07871_),
    .Y(_07882_));
 sky130_fd_sc_hd__nand3_2 _18049_ (.A(_07872_),
    .B(_07877_),
    .C(_07878_),
    .Y(_07883_));
 sky130_fd_sc_hd__and3_2 _18050_ (.A(_07871_),
    .B(_07879_),
    .C(_07880_),
    .X(_07884_));
 sky130_fd_sc_hd__nand3_4 _18051_ (.A(_07871_),
    .B(_07879_),
    .C(_07880_),
    .Y(_07885_));
 sky130_fd_sc_hd__o21a_1 _18052_ (.A1(_01912_),
    .A2(_02152_),
    .B1(_07576_),
    .X(_07886_));
 sky130_fd_sc_hd__and3_1 _18053_ (.A(_07573_),
    .B(net51),
    .C(net32),
    .X(_07887_));
 sky130_fd_sc_hd__o2bb2ai_1 _18054_ (.A1_N(_07883_),
    .A2_N(_07885_),
    .B1(_07886_),
    .B2(_07572_),
    .Y(_07888_));
 sky130_fd_sc_hd__o21a_2 _18055_ (.A1(_07575_),
    .A2(_07887_),
    .B1(_07883_),
    .X(_07889_));
 sky130_fd_sc_hd__o211ai_2 _18056_ (.A1(_07575_),
    .A2(_07887_),
    .B1(_07885_),
    .C1(_07883_),
    .Y(_07890_));
 sky130_fd_sc_hd__o2111ai_4 _18057_ (.A1(_07571_),
    .A2(_07572_),
    .B1(_07576_),
    .C1(_07883_),
    .D1(_07885_),
    .Y(_07891_));
 sky130_fd_sc_hd__o2bb2ai_1 _18058_ (.A1_N(_07883_),
    .A2_N(_07885_),
    .B1(_07887_),
    .B2(_07575_),
    .Y(_07893_));
 sky130_fd_sc_hd__a32oi_4 _18059_ (.A1(_07480_),
    .A2(_07488_),
    .A3(_07489_),
    .B1(_07502_),
    .B2(_07504_),
    .Y(_07894_));
 sky130_fd_sc_hd__a21oi_2 _18060_ (.A1(_07492_),
    .A2(_07505_),
    .B1(_07493_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand3_4 _18061_ (.A(_07895_),
    .B(_07893_),
    .C(_07891_),
    .Y(_07896_));
 sky130_fd_sc_hd__o211ai_4 _18062_ (.A1(_07493_),
    .A2(_07894_),
    .B1(_07890_),
    .C1(_07888_),
    .Y(_07897_));
 sky130_fd_sc_hd__a21oi_2 _18063_ (.A1(_07581_),
    .A2(_07587_),
    .B1(_07582_),
    .Y(_07898_));
 sky130_fd_sc_hd__a21bo_1 _18064_ (.A1(_07896_),
    .A2(_07897_),
    .B1_N(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__nand3b_2 _18065_ (.A_N(_07898_),
    .B(_07897_),
    .C(_07896_),
    .Y(_07900_));
 sky130_fd_sc_hd__a22o_1 _18066_ (.A1(_07583_),
    .A2(_07589_),
    .B1(_07896_),
    .B2(_07897_),
    .X(_07901_));
 sky130_fd_sc_hd__nand4_2 _18067_ (.A(_07583_),
    .B(_07589_),
    .C(_07896_),
    .D(_07897_),
    .Y(_07902_));
 sky130_fd_sc_hd__nand3_4 _18068_ (.A(_07901_),
    .B(_07902_),
    .C(_07869_),
    .Y(_07904_));
 sky130_fd_sc_hd__inv_2 _18069_ (.A(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__nand3b_4 _18070_ (.A_N(_07869_),
    .B(_07899_),
    .C(_07900_),
    .Y(_07906_));
 sky130_fd_sc_hd__a2bb2oi_1 _18071_ (.A1_N(_07544_),
    .A2_N(_07548_),
    .B1(_07555_),
    .B2(_07547_),
    .Y(_07907_));
 sky130_fd_sc_hd__o22a_1 _18072_ (.A1(net28),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01857_),
    .X(_07908_));
 sky130_fd_sc_hd__a22o_1 _18073_ (.A1(net29),
    .A2(net56),
    .B1(_01748_),
    .B2(net57),
    .X(_07909_));
 sky130_fd_sc_hd__or3_4 _18074_ (.A(net28),
    .B(_01857_),
    .C(_02229_),
    .X(_07910_));
 sky130_fd_sc_hd__and4_2 _18075_ (.A(_01748_),
    .B(net29),
    .C(net56),
    .D(net57),
    .X(_07911_));
 sky130_fd_sc_hd__o21a_1 _18076_ (.A1(_02240_),
    .A2(_07910_),
    .B1(_07909_),
    .X(_07912_));
 sky130_fd_sc_hd__a31oi_2 _18077_ (.A1(_07540_),
    .A2(net54),
    .A3(net29),
    .B1(_07538_),
    .Y(_07913_));
 sky130_fd_sc_hd__a31o_1 _18078_ (.A1(_07540_),
    .A2(net54),
    .A3(net29),
    .B1(_07538_),
    .X(_07915_));
 sky130_fd_sc_hd__nand2_1 _18079_ (.A(net30),
    .B(net54),
    .Y(_07916_));
 sky130_fd_sc_hd__a22oi_1 _18080_ (.A1(net32),
    .A2(net52),
    .B1(net53),
    .B2(net31),
    .Y(_07917_));
 sky130_fd_sc_hd__a22o_1 _18081_ (.A1(net32),
    .A2(net52),
    .B1(net53),
    .B2(net31),
    .X(_07918_));
 sky130_fd_sc_hd__nand4_4 _18082_ (.A(net31),
    .B(net32),
    .C(net52),
    .D(net53),
    .Y(_07919_));
 sky130_fd_sc_hd__o211ai_2 _18083_ (.A1(_01868_),
    .A2(_02207_),
    .B1(_07918_),
    .C1(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__a21o_1 _18084_ (.A1(_07918_),
    .A2(_07919_),
    .B1(_07916_),
    .X(_07921_));
 sky130_fd_sc_hd__a22o_1 _18085_ (.A1(net30),
    .A2(net54),
    .B1(_07918_),
    .B2(_07919_),
    .X(_07922_));
 sky130_fd_sc_hd__nand4_2 _18086_ (.A(_07918_),
    .B(_07919_),
    .C(net30),
    .D(net54),
    .Y(_07923_));
 sky130_fd_sc_hd__nand3_4 _18087_ (.A(_07921_),
    .B(_07913_),
    .C(_07920_),
    .Y(_07924_));
 sky130_fd_sc_hd__nand3_4 _18088_ (.A(_07915_),
    .B(_07922_),
    .C(_07923_),
    .Y(_07926_));
 sky130_fd_sc_hd__a2bb2oi_2 _18089_ (.A1_N(_07908_),
    .A2_N(_07911_),
    .B1(_07924_),
    .B2(_07926_),
    .Y(_07927_));
 sky130_fd_sc_hd__a2bb2o_1 _18090_ (.A1_N(_07908_),
    .A2_N(_07911_),
    .B1(_07924_),
    .B2(_07926_),
    .X(_07928_));
 sky130_fd_sc_hd__o2111a_1 _18091_ (.A1(_02240_),
    .A2(_07910_),
    .B1(_07924_),
    .C1(_07926_),
    .D1(_07909_),
    .X(_07929_));
 sky130_fd_sc_hd__o2111ai_4 _18092_ (.A1(_02240_),
    .A2(_07910_),
    .B1(_07924_),
    .C1(_07926_),
    .D1(_07909_),
    .Y(_07930_));
 sky130_fd_sc_hd__o21ai_2 _18093_ (.A1(_07927_),
    .A2(_07929_),
    .B1(_07907_),
    .Y(_07931_));
 sky130_fd_sc_hd__a211oi_4 _18094_ (.A1(_07549_),
    .A2(_07559_),
    .B1(_07927_),
    .C1(_07929_),
    .Y(_07932_));
 sky130_fd_sc_hd__nand3b_2 _18095_ (.A_N(_07907_),
    .B(_07928_),
    .C(_07930_),
    .Y(_07933_));
 sky130_fd_sc_hd__o311a_1 _18096_ (.A1(net27),
    .A2(_02240_),
    .A3(_07550_),
    .B1(_07931_),
    .C1(_07933_),
    .X(_07934_));
 sky130_fd_sc_hd__a211oi_1 _18097_ (.A1(_07931_),
    .A2(_07933_),
    .B1(_07550_),
    .C1(_07551_),
    .Y(_07935_));
 sky130_fd_sc_hd__o2bb2a_1 _18098_ (.A1_N(_07931_),
    .A2_N(_07933_),
    .B1(_07550_),
    .B2(_07551_),
    .X(_07937_));
 sky130_fd_sc_hd__a2bb2o_1 _18099_ (.A1_N(_07550_),
    .A2_N(_07551_),
    .B1(_07931_),
    .B2(_07933_),
    .X(_07938_));
 sky130_fd_sc_hd__nand2_2 _18100_ (.A(_07931_),
    .B(_07553_),
    .Y(_07939_));
 sky130_fd_sc_hd__and3_1 _18101_ (.A(_07931_),
    .B(_07933_),
    .C(_07553_),
    .X(_07940_));
 sky130_fd_sc_hd__o21ai_2 _18102_ (.A1(_07932_),
    .A2(_07939_),
    .B1(_07938_),
    .Y(_07941_));
 sky130_fd_sc_hd__o2bb2ai_1 _18103_ (.A1_N(_07904_),
    .A2_N(_07906_),
    .B1(_07937_),
    .B2(_07940_),
    .Y(_07942_));
 sky130_fd_sc_hd__a31o_1 _18104_ (.A1(_07869_),
    .A2(_07901_),
    .A3(_07902_),
    .B1(_07941_),
    .X(_07943_));
 sky130_fd_sc_hd__o2111ai_4 _18105_ (.A1(_07932_),
    .A2(_07939_),
    .B1(_07938_),
    .C1(_07904_),
    .D1(_07906_),
    .Y(_07944_));
 sky130_fd_sc_hd__o2bb2ai_1 _18106_ (.A1_N(_07904_),
    .A2_N(_07906_),
    .B1(_07934_),
    .B2(_07935_),
    .Y(_07945_));
 sky130_fd_sc_hd__o211ai_2 _18107_ (.A1(_07937_),
    .A2(_07940_),
    .B1(_07904_),
    .C1(_07906_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand3_4 _18108_ (.A(_07945_),
    .B(_07946_),
    .C(_07867_),
    .Y(_07948_));
 sky130_fd_sc_hd__inv_2 _18109_ (.A(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__nand3_4 _18110_ (.A(_07868_),
    .B(_07942_),
    .C(_07944_),
    .Y(_07950_));
 sky130_fd_sc_hd__inv_2 _18111_ (.A(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__a21oi_2 _18112_ (.A1(_07565_),
    .A2(_07567_),
    .B1(_07605_),
    .Y(_07952_));
 sky130_fd_sc_hd__and3_1 _18113_ (.A(_07565_),
    .B(_07567_),
    .C(_07604_),
    .X(_07953_));
 sky130_fd_sc_hd__o21a_1 _18114_ (.A1(_07603_),
    .A2(_07569_),
    .B1(_07606_),
    .X(_07954_));
 sky130_fd_sc_hd__o211a_2 _18115_ (.A1(_07605_),
    .A2(_07953_),
    .B1(_07950_),
    .C1(_07948_),
    .X(_07955_));
 sky130_fd_sc_hd__o2bb2a_1 _18116_ (.A1_N(_07948_),
    .A2_N(_07950_),
    .B1(_07952_),
    .B2(_07603_),
    .X(_07956_));
 sky130_fd_sc_hd__o2bb2a_1 _18117_ (.A1_N(_07948_),
    .A2_N(_07950_),
    .B1(_07953_),
    .B2(_07605_),
    .X(_07957_));
 sky130_fd_sc_hd__o2bb2ai_2 _18118_ (.A1_N(_07948_),
    .A2_N(_07950_),
    .B1(_07953_),
    .B2(_07605_),
    .Y(_07959_));
 sky130_fd_sc_hd__o211ai_4 _18119_ (.A1(_07603_),
    .A2(_07952_),
    .B1(_07950_),
    .C1(_07948_),
    .Y(_07960_));
 sky130_fd_sc_hd__inv_2 _18120_ (.A(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand2_1 _18121_ (.A(_07959_),
    .B(_07960_),
    .Y(_07962_));
 sky130_fd_sc_hd__nand4_2 _18122_ (.A(_07865_),
    .B(_07866_),
    .C(_07959_),
    .D(_07960_),
    .Y(_07963_));
 sky130_fd_sc_hd__o2bb2ai_1 _18123_ (.A1_N(_07865_),
    .A2_N(_07866_),
    .B1(_07957_),
    .B2(_07961_),
    .Y(_07964_));
 sky130_fd_sc_hd__o2bb2ai_4 _18124_ (.A1_N(_07865_),
    .A2_N(_07866_),
    .B1(_07955_),
    .B2(_07956_),
    .Y(_07965_));
 sky130_fd_sc_hd__o211ai_4 _18125_ (.A1(_07857_),
    .A2(_07863_),
    .B1(_07866_),
    .C1(_07962_),
    .Y(_07966_));
 sky130_fd_sc_hd__a2bb2oi_2 _18126_ (.A1_N(_07531_),
    .A2_N(_07625_),
    .B1(_07963_),
    .B2(_07964_),
    .Y(_07967_));
 sky130_fd_sc_hd__o2111ai_4 _18127_ (.A1(_07624_),
    .A2(_07531_),
    .B1(_07533_),
    .C1(_07965_),
    .D1(_07966_),
    .Y(_07968_));
 sky130_fd_sc_hd__a22oi_4 _18128_ (.A1(_07533_),
    .A2(_07666_),
    .B1(_07965_),
    .B2(_07966_),
    .Y(_07970_));
 sky130_fd_sc_hd__nand4_2 _18129_ (.A(_07532_),
    .B(_07626_),
    .C(_07963_),
    .D(_07964_),
    .Y(_07971_));
 sky130_fd_sc_hd__o211ai_1 _18130_ (.A1(_07612_),
    .A2(_07622_),
    .B1(_07968_),
    .C1(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__o2bb2ai_1 _18131_ (.A1_N(_07614_),
    .A2_N(_07663_),
    .B1(_07967_),
    .B2(_07970_),
    .Y(_07973_));
 sky130_fd_sc_hd__o22ai_2 _18132_ (.A1(_07612_),
    .A2(_07622_),
    .B1(_07967_),
    .B2(_07970_),
    .Y(_07974_));
 sky130_fd_sc_hd__nand3_1 _18133_ (.A(_07665_),
    .B(_07968_),
    .C(_07971_),
    .Y(_07975_));
 sky130_fd_sc_hd__o2111ai_4 _18134_ (.A1(_07637_),
    .A2(_07634_),
    .B1(_07633_),
    .C1(_07975_),
    .D1(_07974_),
    .Y(_07976_));
 sky130_fd_sc_hd__nand3_1 _18135_ (.A(_07973_),
    .B(_07662_),
    .C(_07972_),
    .Y(_07977_));
 sky130_fd_sc_hd__a31o_1 _18136_ (.A1(_07536_),
    .A2(_07557_),
    .A3(_07559_),
    .B1(_07564_),
    .X(_07978_));
 sky130_fd_sc_hd__a21o_1 _18137_ (.A1(_07976_),
    .A2(_07977_),
    .B1(_07978_),
    .X(_07979_));
 sky130_fd_sc_hd__nand3_2 _18138_ (.A(_07976_),
    .B(_07977_),
    .C(_07978_),
    .Y(_07981_));
 sky130_fd_sc_hd__o211a_1 _18139_ (.A1(_06628_),
    .A2(_07007_),
    .B1(_07008_),
    .C1(_07646_),
    .X(_07982_));
 sky130_fd_sc_hd__o21ai_2 _18140_ (.A1(_07007_),
    .A2(_07009_),
    .B1(_07646_),
    .Y(_07983_));
 sky130_fd_sc_hd__o2bb2ai_2 _18141_ (.A1_N(_07979_),
    .A2_N(_07981_),
    .B1(_07982_),
    .B2(_07643_),
    .Y(_07984_));
 sky130_fd_sc_hd__nand4_4 _18142_ (.A(_07644_),
    .B(_07979_),
    .C(_07981_),
    .D(_07983_),
    .Y(_07985_));
 sky130_fd_sc_hd__nand2_1 _18143_ (.A(_07984_),
    .B(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__nand4_1 _18144_ (.A(_07335_),
    .B(_07337_),
    .C(_07656_),
    .D(_07658_),
    .Y(_07987_));
 sky130_fd_sc_hd__a31o_1 _18145_ (.A1(_07336_),
    .A2(_07656_),
    .A3(_07332_),
    .B1(_07657_),
    .X(_07988_));
 sky130_fd_sc_hd__a31oi_4 _18146_ (.A1(_07338_),
    .A2(_07340_),
    .A3(_07659_),
    .B1(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__nor2_2 _18147_ (.A(_07341_),
    .B(_07987_),
    .Y(_07990_));
 sky130_fd_sc_hd__a21boi_2 _18148_ (.A1(_06601_),
    .A2(_07990_),
    .B1_N(_07989_),
    .Y(_07992_));
 sky130_fd_sc_hd__xor2_1 _18149_ (.A(_07986_),
    .B(_07992_),
    .X(net94));
 sky130_fd_sc_hd__o21ai_2 _18150_ (.A1(_07665_),
    .A2(_07970_),
    .B1(_07968_),
    .Y(_07993_));
 sky130_fd_sc_hd__a21oi_1 _18151_ (.A1(_07971_),
    .A2(_07664_),
    .B1(_07967_),
    .Y(_07994_));
 sky130_fd_sc_hd__o22ai_2 _18152_ (.A1(_07857_),
    .A2(_07863_),
    .B1(_07955_),
    .B2(_07956_),
    .Y(_07995_));
 sky130_fd_sc_hd__a32oi_4 _18153_ (.A1(_07668_),
    .A2(_07861_),
    .A3(_07862_),
    .B1(_07959_),
    .B2(_07960_),
    .Y(_07996_));
 sky130_fd_sc_hd__a21boi_1 _18154_ (.A1(_07962_),
    .A2(_07866_),
    .B1_N(_07865_),
    .Y(_07997_));
 sky130_fd_sc_hd__o21ai_1 _18155_ (.A1(_07851_),
    .A2(_07852_),
    .B1(_07773_),
    .Y(_07998_));
 sky130_fd_sc_hd__a31oi_1 _18156_ (.A1(_07773_),
    .A2(_07854_),
    .A3(_07856_),
    .B1(_07774_),
    .Y(_07999_));
 sky130_fd_sc_hd__a31o_1 _18157_ (.A1(_07773_),
    .A2(_07854_),
    .A3(_07856_),
    .B1(_07774_),
    .X(_08000_));
 sky130_fd_sc_hd__nand3_1 _18158_ (.A(_07721_),
    .B(_07765_),
    .C(_07767_),
    .Y(_08002_));
 sky130_fd_sc_hd__a31o_1 _18159_ (.A1(_07721_),
    .A2(_07765_),
    .A3(_07767_),
    .B1(_07722_),
    .X(_08003_));
 sky130_fd_sc_hd__a211o_4 _18160_ (.A1(_07677_),
    .A2(_07679_),
    .B1(_06880_),
    .C1(_07129_),
    .X(_08004_));
 sky130_fd_sc_hd__a21oi_2 _18161_ (.A1(_07390_),
    .A2(_07675_),
    .B1(_06881_),
    .Y(_08005_));
 sky130_fd_sc_hd__and3_4 _18162_ (.A(_07677_),
    .B(_07679_),
    .C(_06880_),
    .X(_08006_));
 sky130_fd_sc_hd__or3_4 _18163_ (.A(_06881_),
    .B(_07676_),
    .C(_07678_),
    .X(_08007_));
 sky130_fd_sc_hd__a22oi_4 _18164_ (.A1(_08005_),
    .A2(_07679_),
    .B1(_07681_),
    .B2(_06881_),
    .Y(_08008_));
 sky130_fd_sc_hd__a22o_2 _18165_ (.A1(_08005_),
    .A2(_07679_),
    .B1(_07681_),
    .B2(_06881_),
    .X(_08009_));
 sky130_fd_sc_hd__nand2_1 _18166_ (.A(net63),
    .B(net22),
    .Y(_08010_));
 sky130_fd_sc_hd__a22oi_4 _18167_ (.A1(net62),
    .A2(net24),
    .B1(net25),
    .B2(net61),
    .Y(_08011_));
 sky130_fd_sc_hd__a22o_1 _18168_ (.A1(net62),
    .A2(net24),
    .B1(net25),
    .B2(net61),
    .X(_08013_));
 sky130_fd_sc_hd__and4_1 _18169_ (.A(net61),
    .B(net62),
    .C(net24),
    .D(net25),
    .X(_08014_));
 sky130_fd_sc_hd__nand4_2 _18170_ (.A(net61),
    .B(net62),
    .C(net24),
    .D(net25),
    .Y(_08015_));
 sky130_fd_sc_hd__o211ai_2 _18171_ (.A1(_01890_),
    .A2(_02196_),
    .B1(_08013_),
    .C1(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__o21bai_2 _18172_ (.A1(_08011_),
    .A2(_08014_),
    .B1_N(_08010_),
    .Y(_08017_));
 sky130_fd_sc_hd__o21ai_1 _18173_ (.A1(_08011_),
    .A2(_08014_),
    .B1(_08010_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand4_1 _18174_ (.A(_08013_),
    .B(_08015_),
    .C(net63),
    .D(net22),
    .Y(_08019_));
 sky130_fd_sc_hd__nand3_2 _18175_ (.A(_07699_),
    .B(_08016_),
    .C(_08017_),
    .Y(_08020_));
 sky130_fd_sc_hd__and3_1 _18176_ (.A(_08018_),
    .B(_08019_),
    .C(_07698_),
    .X(_08021_));
 sky130_fd_sc_hd__nand3_2 _18177_ (.A(_08018_),
    .B(_08019_),
    .C(_07698_),
    .Y(_08022_));
 sky130_fd_sc_hd__o31ai_4 _18178_ (.A1(_01890_),
    .A2(_02185_),
    .A3(_07702_),
    .B1(_07701_),
    .Y(_08024_));
 sky130_fd_sc_hd__o31a_1 _18179_ (.A1(_01890_),
    .A2(_02185_),
    .A3(_07702_),
    .B1(_07701_),
    .X(_08025_));
 sky130_fd_sc_hd__a21oi_1 _18180_ (.A1(_08020_),
    .A2(_08022_),
    .B1(_08024_),
    .Y(_08026_));
 sky130_fd_sc_hd__a21o_1 _18181_ (.A1(_08020_),
    .A2(_08022_),
    .B1(_08024_),
    .X(_08027_));
 sky130_fd_sc_hd__a31oi_2 _18182_ (.A1(_07699_),
    .A2(_08016_),
    .A3(_08017_),
    .B1(_08025_),
    .Y(_08028_));
 sky130_fd_sc_hd__and3_1 _18183_ (.A(_08020_),
    .B(_08022_),
    .C(_08024_),
    .X(_08029_));
 sky130_fd_sc_hd__nand3_2 _18184_ (.A(_08020_),
    .B(_08022_),
    .C(_08024_),
    .Y(_08030_));
 sky130_fd_sc_hd__o2bb2ai_4 _18185_ (.A1_N(_08004_),
    .A2_N(_08007_),
    .B1(_08026_),
    .B2(_08029_),
    .Y(_08031_));
 sky130_fd_sc_hd__o2111ai_4 _18186_ (.A1(_06880_),
    .A2(_07682_),
    .B1(_08007_),
    .C1(_08027_),
    .D1(_08030_),
    .Y(_08032_));
 sky130_fd_sc_hd__a22oi_2 _18187_ (.A1(_07688_),
    .A2(_07685_),
    .B1(_07715_),
    .B2(_07714_),
    .Y(_08033_));
 sky130_fd_sc_hd__nand3_2 _18188_ (.A(_07689_),
    .B(_07711_),
    .C(_07712_),
    .Y(_08035_));
 sky130_fd_sc_hd__a22oi_4 _18189_ (.A1(_08031_),
    .A2(_08032_),
    .B1(_08035_),
    .B2(_07686_),
    .Y(_08036_));
 sky130_fd_sc_hd__o2bb2ai_4 _18190_ (.A1_N(_08031_),
    .A2_N(_08032_),
    .B1(_08033_),
    .B2(_07687_),
    .Y(_08037_));
 sky130_fd_sc_hd__nand4_4 _18191_ (.A(_07686_),
    .B(_08031_),
    .C(_08032_),
    .D(_08035_),
    .Y(_08038_));
 sky130_fd_sc_hd__nor2_1 _18192_ (.A(_07728_),
    .B(_07731_),
    .Y(_08039_));
 sky130_fd_sc_hd__o21ai_2 _18193_ (.A1(_07728_),
    .A2(_07731_),
    .B1(_07730_),
    .Y(_08040_));
 sky130_fd_sc_hd__nand2_1 _18194_ (.A(net35),
    .B(net19),
    .Y(_08041_));
 sky130_fd_sc_hd__nand2_1 _18195_ (.A(net34),
    .B(net21),
    .Y(_08042_));
 sky130_fd_sc_hd__nand4_4 _18196_ (.A(net64),
    .B(net34),
    .C(net20),
    .D(net21),
    .Y(_08043_));
 sky130_fd_sc_hd__a22oi_2 _18197_ (.A1(net34),
    .A2(net20),
    .B1(net21),
    .B2(net64),
    .Y(_08044_));
 sky130_fd_sc_hd__a22o_1 _18198_ (.A1(net34),
    .A2(net20),
    .B1(net21),
    .B2(net64),
    .X(_08046_));
 sky130_fd_sc_hd__o2bb2ai_4 _18199_ (.A1_N(_08043_),
    .A2_N(_08046_),
    .B1(_01934_),
    .B2(_02142_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand4_4 _18200_ (.A(_08046_),
    .B(net19),
    .C(net35),
    .D(_08043_),
    .Y(_08048_));
 sky130_fd_sc_hd__a21oi_4 _18201_ (.A1(_08047_),
    .A2(_08048_),
    .B1(_08040_),
    .Y(_08049_));
 sky130_fd_sc_hd__a21o_2 _18202_ (.A1(_08047_),
    .A2(_08048_),
    .B1(_08040_),
    .X(_08050_));
 sky130_fd_sc_hd__nand2_1 _18203_ (.A(net38),
    .B(net16),
    .Y(_08051_));
 sky130_fd_sc_hd__a22oi_2 _18204_ (.A1(net37),
    .A2(net17),
    .B1(net18),
    .B2(net36),
    .Y(_08052_));
 sky130_fd_sc_hd__a22o_2 _18205_ (.A1(net37),
    .A2(net17),
    .B1(net18),
    .B2(net36),
    .X(_08053_));
 sky130_fd_sc_hd__nand2_1 _18206_ (.A(net37),
    .B(net18),
    .Y(_08054_));
 sky130_fd_sc_hd__nand4_4 _18207_ (.A(net36),
    .B(net37),
    .C(net17),
    .D(net18),
    .Y(_08055_));
 sky130_fd_sc_hd__a22oi_4 _18208_ (.A1(net38),
    .A2(net16),
    .B1(_08053_),
    .B2(_08055_),
    .Y(_08057_));
 sky130_fd_sc_hd__a22o_1 _18209_ (.A1(net38),
    .A2(net16),
    .B1(_08053_),
    .B2(_08055_),
    .X(_08058_));
 sky130_fd_sc_hd__o2111a_1 _18210_ (.A1(_07741_),
    .A2(_08054_),
    .B1(net38),
    .C1(net16),
    .D1(_08053_),
    .X(_08059_));
 sky130_fd_sc_hd__o2111ai_4 _18211_ (.A1(_07741_),
    .A2(_08054_),
    .B1(net38),
    .C1(net16),
    .D1(_08053_),
    .Y(_08060_));
 sky130_fd_sc_hd__nor2_2 _18212_ (.A(_08057_),
    .B(_08059_),
    .Y(_08061_));
 sky130_fd_sc_hd__o211a_2 _18213_ (.A1(_07729_),
    .A2(_08039_),
    .B1(_08047_),
    .C1(_08048_),
    .X(_08062_));
 sky130_fd_sc_hd__o211ai_2 _18214_ (.A1(_07729_),
    .A2(_08039_),
    .B1(_08047_),
    .C1(_08048_),
    .Y(_08063_));
 sky130_fd_sc_hd__a32o_2 _18215_ (.A1(_08047_),
    .A2(_08048_),
    .A3(_08040_),
    .B1(_08058_),
    .B2(_08060_),
    .X(_08064_));
 sky130_fd_sc_hd__a311o_1 _18216_ (.A1(_08040_),
    .A2(_08047_),
    .A3(_08048_),
    .B1(_08061_),
    .C1(_08049_),
    .X(_08065_));
 sky130_fd_sc_hd__o21ai_4 _18217_ (.A1(_08049_),
    .A2(_08062_),
    .B1(_08061_),
    .Y(_08066_));
 sky130_fd_sc_hd__o22ai_4 _18218_ (.A1(_08057_),
    .A2(_08059_),
    .B1(_08062_),
    .B2(_08049_),
    .Y(_08068_));
 sky130_fd_sc_hd__nand4_4 _18219_ (.A(_08050_),
    .B(_08058_),
    .C(_08060_),
    .D(_08063_),
    .Y(_08069_));
 sky130_fd_sc_hd__o21ai_4 _18220_ (.A1(_07693_),
    .A2(_07709_),
    .B1(_07708_),
    .Y(_08070_));
 sky130_fd_sc_hd__a21oi_4 _18221_ (.A1(_07710_),
    .A2(_07692_),
    .B1(_07707_),
    .Y(_08071_));
 sky130_fd_sc_hd__o211a_1 _18222_ (.A1(_08064_),
    .A2(_08049_),
    .B1(_08071_),
    .C1(_08066_),
    .X(_08072_));
 sky130_fd_sc_hd__o211ai_4 _18223_ (.A1(_08064_),
    .A2(_08049_),
    .B1(_08071_),
    .C1(_08066_),
    .Y(_08073_));
 sky130_fd_sc_hd__nand3_4 _18224_ (.A(_08068_),
    .B(_08069_),
    .C(_08070_),
    .Y(_08074_));
 sky130_fd_sc_hd__inv_2 _18225_ (.A(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__a32oi_4 _18226_ (.A1(_07726_),
    .A2(_07735_),
    .A3(_07736_),
    .B1(_07737_),
    .B2(_07751_),
    .Y(_08076_));
 sky130_fd_sc_hd__a32o_2 _18227_ (.A1(_07726_),
    .A2(_07735_),
    .A3(_07736_),
    .B1(_07737_),
    .B2(_07751_),
    .X(_08077_));
 sky130_fd_sc_hd__a21o_1 _18228_ (.A1(_08073_),
    .A2(_08074_),
    .B1(_08076_),
    .X(_08079_));
 sky130_fd_sc_hd__nand3_1 _18229_ (.A(_08073_),
    .B(_08074_),
    .C(_08076_),
    .Y(_08080_));
 sky130_fd_sc_hd__a21oi_1 _18230_ (.A1(_08073_),
    .A2(_08074_),
    .B1(_08077_),
    .Y(_08081_));
 sky130_fd_sc_hd__a21o_1 _18231_ (.A1(_08073_),
    .A2(_08074_),
    .B1(_08077_),
    .X(_08082_));
 sky130_fd_sc_hd__nand2_1 _18232_ (.A(_08073_),
    .B(_08077_),
    .Y(_08083_));
 sky130_fd_sc_hd__and3_1 _18233_ (.A(_08073_),
    .B(_08074_),
    .C(_08077_),
    .X(_08084_));
 sky130_fd_sc_hd__nand3_1 _18234_ (.A(_08073_),
    .B(_08074_),
    .C(_08077_),
    .Y(_08085_));
 sky130_fd_sc_hd__a22oi_2 _18235_ (.A1(_08037_),
    .A2(_08038_),
    .B1(_08082_),
    .B2(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__o2bb2ai_2 _18236_ (.A1_N(_08037_),
    .A2_N(_08038_),
    .B1(_08081_),
    .B2(_08084_),
    .Y(_08087_));
 sky130_fd_sc_hd__o211ai_2 _18237_ (.A1(_08083_),
    .A2(_08075_),
    .B1(_08038_),
    .C1(_08082_),
    .Y(_08088_));
 sky130_fd_sc_hd__o2111a_1 _18238_ (.A1(_08083_),
    .A2(_08075_),
    .B1(_08038_),
    .C1(_08037_),
    .D1(_08082_),
    .X(_08090_));
 sky130_fd_sc_hd__o2111ai_1 _18239_ (.A1(_08083_),
    .A2(_08075_),
    .B1(_08038_),
    .C1(_08037_),
    .D1(_08082_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand2_1 _18240_ (.A(_08087_),
    .B(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__o2111a_1 _18241_ (.A1(_08036_),
    .A2(_08088_),
    .B1(_08087_),
    .C1(_07723_),
    .D1(_08002_),
    .X(_08093_));
 sky130_fd_sc_hd__o2111ai_4 _18242_ (.A1(_08036_),
    .A2(_08088_),
    .B1(_08087_),
    .C1(_07723_),
    .D1(_08002_),
    .Y(_08094_));
 sky130_fd_sc_hd__o21ai_4 _18243_ (.A1(_08086_),
    .A2(_08090_),
    .B1(_08003_),
    .Y(_08095_));
 sky130_fd_sc_hd__a31oi_4 _18244_ (.A1(_07725_),
    .A2(_07752_),
    .A3(_07753_),
    .B1(_07761_),
    .Y(_08096_));
 sky130_fd_sc_hd__a32oi_4 _18245_ (.A1(_07724_),
    .A2(_07754_),
    .A3(_07755_),
    .B1(_07758_),
    .B2(_07759_),
    .Y(_08097_));
 sky130_fd_sc_hd__o2bb2ai_1 _18246_ (.A1_N(_07780_),
    .A2_N(_07784_),
    .B1(_07781_),
    .B2(_07482_),
    .Y(_08098_));
 sky130_fd_sc_hd__o2bb2a_1 _18247_ (.A1_N(_07780_),
    .A2_N(_07784_),
    .B1(_07781_),
    .B2(_07482_),
    .X(_08099_));
 sky130_fd_sc_hd__nand2_1 _18248_ (.A(net9),
    .B(net45),
    .Y(_08101_));
 sky130_fd_sc_hd__nand2_2 _18249_ (.A(net42),
    .B(net11),
    .Y(_08102_));
 sky130_fd_sc_hd__and4_2 _18250_ (.A(net10),
    .B(net42),
    .C(net11),
    .D(net43),
    .X(_08103_));
 sky130_fd_sc_hd__nand4_2 _18251_ (.A(net10),
    .B(net42),
    .C(net11),
    .D(net43),
    .Y(_08104_));
 sky130_fd_sc_hd__a22oi_2 _18252_ (.A1(net42),
    .A2(net11),
    .B1(net43),
    .B2(net10),
    .Y(_08105_));
 sky130_fd_sc_hd__a22o_2 _18253_ (.A1(net42),
    .A2(net11),
    .B1(net43),
    .B2(net10),
    .X(_08106_));
 sky130_fd_sc_hd__o211ai_4 _18254_ (.A1(_01999_),
    .A2(_02054_),
    .B1(_08104_),
    .C1(_08106_),
    .Y(_08107_));
 sky130_fd_sc_hd__o21bai_2 _18255_ (.A1(_08103_),
    .A2(_08105_),
    .B1_N(_08101_),
    .Y(_08108_));
 sky130_fd_sc_hd__o22ai_2 _18256_ (.A1(_01999_),
    .A2(_02054_),
    .B1(_08103_),
    .B2(_08105_),
    .Y(_08109_));
 sky130_fd_sc_hd__and4_1 _18257_ (.A(_08106_),
    .B(net45),
    .C(net9),
    .D(_08104_),
    .X(_08110_));
 sky130_fd_sc_hd__nand4_1 _18258_ (.A(_08106_),
    .B(net45),
    .C(net9),
    .D(_08104_),
    .Y(_08112_));
 sky130_fd_sc_hd__nand3_2 _18259_ (.A(_08099_),
    .B(_08107_),
    .C(_08108_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand2_1 _18260_ (.A(_08109_),
    .B(_08098_),
    .Y(_08114_));
 sky130_fd_sc_hd__and3_2 _18261_ (.A(_08109_),
    .B(_08112_),
    .C(_08098_),
    .X(_08115_));
 sky130_fd_sc_hd__nand3_1 _18262_ (.A(_08109_),
    .B(_08112_),
    .C(_08098_),
    .Y(_08116_));
 sky130_fd_sc_hd__nand2_1 _18263_ (.A(net8),
    .B(net46),
    .Y(_08117_));
 sky130_fd_sc_hd__a22oi_2 _18264_ (.A1(net8),
    .A2(net46),
    .B1(net47),
    .B2(net7),
    .Y(_08118_));
 sky130_fd_sc_hd__a22o_1 _18265_ (.A1(net8),
    .A2(net46),
    .B1(net47),
    .B2(net7),
    .X(_08119_));
 sky130_fd_sc_hd__nand2_1 _18266_ (.A(net8),
    .B(net47),
    .Y(_08120_));
 sky130_fd_sc_hd__and4_1 _18267_ (.A(net7),
    .B(net8),
    .C(net46),
    .D(net47),
    .X(_08121_));
 sky130_fd_sc_hd__nand4_2 _18268_ (.A(net7),
    .B(net8),
    .C(net46),
    .D(net47),
    .Y(_08123_));
 sky130_fd_sc_hd__nand2_1 _18269_ (.A(net6),
    .B(net48),
    .Y(_08124_));
 sky130_fd_sc_hd__a22oi_2 _18270_ (.A1(net6),
    .A2(net48),
    .B1(_08119_),
    .B2(_08123_),
    .Y(_08125_));
 sky130_fd_sc_hd__o22ai_1 _18271_ (.A1(_01966_),
    .A2(_02109_),
    .B1(_08118_),
    .B2(_08121_),
    .Y(_08126_));
 sky130_fd_sc_hd__o2111a_1 _18272_ (.A1(_07794_),
    .A2(_08120_),
    .B1(net6),
    .C1(net48),
    .D1(_08119_),
    .X(_08127_));
 sky130_fd_sc_hd__o2111ai_1 _18273_ (.A1(_07794_),
    .A2(_08120_),
    .B1(net6),
    .C1(net48),
    .D1(_08119_),
    .Y(_08128_));
 sky130_fd_sc_hd__nor2_1 _18274_ (.A(_08125_),
    .B(_08127_),
    .Y(_08129_));
 sky130_fd_sc_hd__nand2_1 _18275_ (.A(_08126_),
    .B(_08128_),
    .Y(_08130_));
 sky130_fd_sc_hd__a21oi_2 _18276_ (.A1(_08113_),
    .A2(_08116_),
    .B1(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__o221a_1 _18277_ (.A1(_08125_),
    .A2(_08127_),
    .B1(_08110_),
    .B2(_08114_),
    .C1(_08113_),
    .X(_08132_));
 sky130_fd_sc_hd__o2bb2a_2 _18278_ (.A1_N(_08113_),
    .A2_N(_08116_),
    .B1(_08125_),
    .B2(_08127_),
    .X(_08134_));
 sky130_fd_sc_hd__a31oi_4 _18279_ (.A1(_08099_),
    .A2(_08107_),
    .A3(_08108_),
    .B1(_08130_),
    .Y(_08135_));
 sky130_fd_sc_hd__and3_1 _18280_ (.A(_08113_),
    .B(_08116_),
    .C(_08129_),
    .X(_08136_));
 sky130_fd_sc_hd__o311a_1 _18281_ (.A1(_02010_),
    .A2(_02021_),
    .A3(_07458_),
    .B1(_07461_),
    .C1(_07829_),
    .X(_08137_));
 sky130_fd_sc_hd__o21ai_1 _18282_ (.A1(_07816_),
    .A2(_07830_),
    .B1(_07829_),
    .Y(_08138_));
 sky130_fd_sc_hd__o31a_1 _18283_ (.A1(_07458_),
    .A2(_07813_),
    .A3(_07830_),
    .B1(_07829_),
    .X(_08139_));
 sky130_fd_sc_hd__o21ai_2 _18284_ (.A1(_02010_),
    .A2(_02032_),
    .B1(_07821_),
    .Y(_08140_));
 sky130_fd_sc_hd__and3_1 _18285_ (.A(_07822_),
    .B(net11),
    .C(net41),
    .X(_08141_));
 sky130_fd_sc_hd__a31o_1 _18286_ (.A1(_07822_),
    .A2(net11),
    .A3(net41),
    .B1(_07820_),
    .X(_08142_));
 sky130_fd_sc_hd__nand2_1 _18287_ (.A(_07822_),
    .B(_08140_),
    .Y(_08143_));
 sky130_fd_sc_hd__nor2_1 _18288_ (.A(_07740_),
    .B(_07742_),
    .Y(_08145_));
 sky130_fd_sc_hd__o22a_1 _18289_ (.A1(_07363_),
    .A2(_07743_),
    .B1(_07740_),
    .B2(_07742_),
    .X(_08146_));
 sky130_fd_sc_hd__nand2_1 _18290_ (.A(net41),
    .B(net13),
    .Y(_08147_));
 sky130_fd_sc_hd__a22oi_4 _18291_ (.A1(net40),
    .A2(net14),
    .B1(net15),
    .B2(net39),
    .Y(_08148_));
 sky130_fd_sc_hd__a22o_1 _18292_ (.A1(net40),
    .A2(net14),
    .B1(net15),
    .B2(net39),
    .X(_08149_));
 sky130_fd_sc_hd__and4_2 _18293_ (.A(net39),
    .B(net40),
    .C(net14),
    .D(net15),
    .X(_08150_));
 sky130_fd_sc_hd__nand4_4 _18294_ (.A(net39),
    .B(net40),
    .C(net14),
    .D(net15),
    .Y(_08151_));
 sky130_fd_sc_hd__o211ai_4 _18295_ (.A1(_02010_),
    .A2(_02043_),
    .B1(_08149_),
    .C1(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__o21bai_4 _18296_ (.A1(_08148_),
    .A2(_08150_),
    .B1_N(_08147_),
    .Y(_08153_));
 sky130_fd_sc_hd__nand4_2 _18297_ (.A(_08149_),
    .B(_08151_),
    .C(net41),
    .D(net13),
    .Y(_08154_));
 sky130_fd_sc_hd__o21ai_1 _18298_ (.A1(_08148_),
    .A2(_08150_),
    .B1(_08147_),
    .Y(_08156_));
 sky130_fd_sc_hd__a2bb2oi_2 _18299_ (.A1_N(_07744_),
    .A2_N(_08145_),
    .B1(_08152_),
    .B2(_08153_),
    .Y(_08157_));
 sky130_fd_sc_hd__o211ai_4 _18300_ (.A1(_07744_),
    .A2(_08145_),
    .B1(_08154_),
    .C1(_08156_),
    .Y(_08158_));
 sky130_fd_sc_hd__nand3_2 _18301_ (.A(_08146_),
    .B(_08152_),
    .C(_08153_),
    .Y(_08159_));
 sky130_fd_sc_hd__a31oi_4 _18302_ (.A1(_08146_),
    .A2(_08152_),
    .A3(_08153_),
    .B1(_08143_),
    .Y(_08160_));
 sky130_fd_sc_hd__a31o_1 _18303_ (.A1(_08146_),
    .A2(_08152_),
    .A3(_08153_),
    .B1(_08143_),
    .X(_08161_));
 sky130_fd_sc_hd__o211a_1 _18304_ (.A1(_07820_),
    .A2(_08141_),
    .B1(_08158_),
    .C1(_08159_),
    .X(_08162_));
 sky130_fd_sc_hd__a22oi_4 _18305_ (.A1(_07822_),
    .A2(_08140_),
    .B1(_08158_),
    .B2(_08159_),
    .Y(_08163_));
 sky130_fd_sc_hd__a22o_1 _18306_ (.A1(_07822_),
    .A2(_08140_),
    .B1(_08158_),
    .B2(_08159_),
    .X(_08164_));
 sky130_fd_sc_hd__a221oi_4 _18307_ (.A1(_08160_),
    .A2(_08158_),
    .B1(_07831_),
    .B2(_07829_),
    .C1(_08163_),
    .Y(_08165_));
 sky130_fd_sc_hd__o211ai_2 _18308_ (.A1(_08157_),
    .A2(_08161_),
    .B1(_08138_),
    .C1(_08164_),
    .Y(_08167_));
 sky130_fd_sc_hd__o22a_2 _18309_ (.A1(_07830_),
    .A2(_08137_),
    .B1(_08162_),
    .B2(_08163_),
    .X(_08168_));
 sky130_fd_sc_hd__o22ai_4 _18310_ (.A1(_07830_),
    .A2(_08137_),
    .B1(_08162_),
    .B2(_08163_),
    .Y(_08169_));
 sky130_fd_sc_hd__o21ai_2 _18311_ (.A1(_08131_),
    .A2(_08132_),
    .B1(_08169_),
    .Y(_08170_));
 sky130_fd_sc_hd__o211a_1 _18312_ (.A1(_08131_),
    .A2(_08132_),
    .B1(_08167_),
    .C1(_08169_),
    .X(_08171_));
 sky130_fd_sc_hd__o211ai_1 _18313_ (.A1(_08131_),
    .A2(_08132_),
    .B1(_08167_),
    .C1(_08169_),
    .Y(_08172_));
 sky130_fd_sc_hd__a2bb2oi_1 _18314_ (.A1_N(_08134_),
    .A2_N(_08136_),
    .B1(_08167_),
    .B2(_08169_),
    .Y(_08173_));
 sky130_fd_sc_hd__o22ai_4 _18315_ (.A1(_08134_),
    .A2(_08136_),
    .B1(_08165_),
    .B2(_08168_),
    .Y(_08174_));
 sky130_fd_sc_hd__a2bb2oi_2 _18316_ (.A1_N(_07756_),
    .A2_N(_08096_),
    .B1(_08172_),
    .B2(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__o22ai_4 _18317_ (.A1(_07756_),
    .A2(_08096_),
    .B1(_08171_),
    .B2(_08173_),
    .Y(_08176_));
 sky130_fd_sc_hd__o211a_2 _18318_ (.A1(_08165_),
    .A2(_08170_),
    .B1(_08097_),
    .C1(_08174_),
    .X(_08178_));
 sky130_fd_sc_hd__o211ai_4 _18319_ (.A1(_08165_),
    .A2(_08170_),
    .B1(_08097_),
    .C1(_08174_),
    .Y(_08179_));
 sky130_fd_sc_hd__o31a_1 _18320_ (.A1(_07803_),
    .A2(_07805_),
    .A3(_07835_),
    .B1(_07839_),
    .X(_08180_));
 sky130_fd_sc_hd__o31a_1 _18321_ (.A1(_07806_),
    .A2(_07809_),
    .A3(_07838_),
    .B1(_07836_),
    .X(_08181_));
 sky130_fd_sc_hd__and3_1 _18322_ (.A(_08176_),
    .B(_08179_),
    .C(_08180_),
    .X(_08182_));
 sky130_fd_sc_hd__o211ai_4 _18323_ (.A1(_07835_),
    .A2(_07842_),
    .B1(_08176_),
    .C1(_08179_),
    .Y(_08183_));
 sky130_fd_sc_hd__o221a_1 _18324_ (.A1(_07810_),
    .A2(_07838_),
    .B1(_08175_),
    .B2(_08178_),
    .C1(_07836_),
    .X(_08184_));
 sky130_fd_sc_hd__o21ai_2 _18325_ (.A1(_08175_),
    .A2(_08178_),
    .B1(_08181_),
    .Y(_08185_));
 sky130_fd_sc_hd__and3_1 _18326_ (.A(_08176_),
    .B(_08179_),
    .C(_08181_),
    .X(_08186_));
 sky130_fd_sc_hd__o2111ai_4 _18327_ (.A1(_07810_),
    .A2(_07838_),
    .B1(_08176_),
    .C1(_08179_),
    .D1(_07836_),
    .Y(_08187_));
 sky130_fd_sc_hd__o22a_1 _18328_ (.A1(_07835_),
    .A2(_07842_),
    .B1(_08175_),
    .B2(_08178_),
    .X(_08189_));
 sky130_fd_sc_hd__o22ai_2 _18329_ (.A1(_07835_),
    .A2(_07842_),
    .B1(_08175_),
    .B2(_08178_),
    .Y(_08190_));
 sky130_fd_sc_hd__nand4_2 _18330_ (.A(_08094_),
    .B(_08095_),
    .C(_08187_),
    .D(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__o2bb2ai_2 _18331_ (.A1_N(_08094_),
    .A2_N(_08095_),
    .B1(_08186_),
    .B2(_08189_),
    .Y(_08192_));
 sky130_fd_sc_hd__o2bb2ai_2 _18332_ (.A1_N(_08094_),
    .A2_N(_08095_),
    .B1(_08182_),
    .B2(_08184_),
    .Y(_08193_));
 sky130_fd_sc_hd__nand4_4 _18333_ (.A(_08094_),
    .B(_08095_),
    .C(_08183_),
    .D(_08185_),
    .Y(_08194_));
 sky130_fd_sc_hd__nand3_2 _18334_ (.A(_08000_),
    .B(_08193_),
    .C(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__and3_1 _18335_ (.A(_07999_),
    .B(_08191_),
    .C(_08192_),
    .X(_08196_));
 sky130_fd_sc_hd__nand4_4 _18336_ (.A(_07775_),
    .B(_07998_),
    .C(_08191_),
    .D(_08192_),
    .Y(_08197_));
 sky130_fd_sc_hd__a31oi_2 _18337_ (.A1(_07777_),
    .A2(_07843_),
    .A3(_07844_),
    .B1(_07850_),
    .Y(_08198_));
 sky130_fd_sc_hd__a32oi_4 _18338_ (.A1(_07776_),
    .A2(_07840_),
    .A3(_07841_),
    .B1(_07845_),
    .B2(_07849_),
    .Y(_08200_));
 sky130_fd_sc_hd__a21boi_2 _18339_ (.A1(_07912_),
    .A2(_07924_),
    .B1_N(_07926_),
    .Y(_08201_));
 sky130_fd_sc_hd__o21ai_2 _18340_ (.A1(_07916_),
    .A2(_07917_),
    .B1(_07919_),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_1 _18341_ (.A(net31),
    .B(net54),
    .Y(_08203_));
 sky130_fd_sc_hd__a22oi_1 _18342_ (.A1(net2),
    .A2(net52),
    .B1(net53),
    .B2(net32),
    .Y(_08204_));
 sky130_fd_sc_hd__a22o_1 _18343_ (.A1(net2),
    .A2(net52),
    .B1(net53),
    .B2(net32),
    .X(_08205_));
 sky130_fd_sc_hd__nand4_4 _18344_ (.A(net2),
    .B(net32),
    .C(net52),
    .D(net53),
    .Y(_08206_));
 sky130_fd_sc_hd__o211ai_1 _18345_ (.A1(_01879_),
    .A2(_02207_),
    .B1(_08205_),
    .C1(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__a21o_1 _18346_ (.A1(_08205_),
    .A2(_08206_),
    .B1(_08203_),
    .X(_08208_));
 sky130_fd_sc_hd__a22o_1 _18347_ (.A1(net31),
    .A2(net54),
    .B1(_08205_),
    .B2(_08206_),
    .X(_08209_));
 sky130_fd_sc_hd__nand4_1 _18348_ (.A(_08205_),
    .B(_08206_),
    .C(net31),
    .D(net54),
    .Y(_08211_));
 sky130_fd_sc_hd__nand3b_2 _18349_ (.A_N(_08202_),
    .B(_08207_),
    .C(_08208_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand3_2 _18350_ (.A(_08209_),
    .B(_08211_),
    .C(_08202_),
    .Y(_08213_));
 sky130_fd_sc_hd__nand2_1 _18351_ (.A(net30),
    .B(net56),
    .Y(_08214_));
 sky130_fd_sc_hd__and4_1 _18352_ (.A(_01857_),
    .B(net30),
    .C(net56),
    .D(net57),
    .X(_08215_));
 sky130_fd_sc_hd__or4_2 _18353_ (.A(net29),
    .B(_01868_),
    .C(_02229_),
    .D(_02240_),
    .X(_08216_));
 sky130_fd_sc_hd__o22a_1 _18354_ (.A1(net29),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01868_),
    .X(_08217_));
 sky130_fd_sc_hd__nor2_1 _18355_ (.A(_08215_),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__and3_2 _18356_ (.A(_08212_),
    .B(_08213_),
    .C(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__a21oi_4 _18357_ (.A1(_08212_),
    .A2(_08213_),
    .B1(_08218_),
    .Y(_08220_));
 sky130_fd_sc_hd__o21a_1 _18358_ (.A1(_08219_),
    .A2(_08220_),
    .B1(_08201_),
    .X(_08222_));
 sky130_fd_sc_hd__o21ai_2 _18359_ (.A1(_08219_),
    .A2(_08220_),
    .B1(_08201_),
    .Y(_08223_));
 sky130_fd_sc_hd__a211oi_4 _18360_ (.A1(_07926_),
    .A2(_07930_),
    .B1(_08219_),
    .C1(_08220_),
    .Y(_08224_));
 sky130_fd_sc_hd__o22a_1 _18361_ (.A1(_02240_),
    .A2(_07910_),
    .B1(_08222_),
    .B2(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__o22ai_2 _18362_ (.A1(_02240_),
    .A2(_07910_),
    .B1(_08222_),
    .B2(_08224_),
    .Y(_08226_));
 sky130_fd_sc_hd__nand2_2 _18363_ (.A(_08223_),
    .B(_07911_),
    .Y(_08227_));
 sky130_fd_sc_hd__nor2_1 _18364_ (.A(_08224_),
    .B(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__nor3_1 _18365_ (.A(_07911_),
    .B(_08222_),
    .C(_08224_),
    .Y(_08229_));
 sky130_fd_sc_hd__o21a_1 _18366_ (.A1(_08222_),
    .A2(_08224_),
    .B1(_07911_),
    .X(_08230_));
 sky130_fd_sc_hd__o21ai_1 _18367_ (.A1(_08224_),
    .A2(_08227_),
    .B1(_08226_),
    .Y(_08231_));
 sky130_fd_sc_hd__nand2_2 _18368_ (.A(_07897_),
    .B(_07898_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand2_1 _18369_ (.A(_07896_),
    .B(_08233_),
    .Y(_08234_));
 sky130_fd_sc_hd__o311a_2 _18370_ (.A1(_01912_),
    .A2(_02152_),
    .A3(_07572_),
    .B1(_07576_),
    .C1(_07885_),
    .X(_08235_));
 sky130_fd_sc_hd__o31a_2 _18371_ (.A1(_07572_),
    .A2(_07882_),
    .A3(_07886_),
    .B1(_07885_),
    .X(_08236_));
 sky130_fd_sc_hd__a32o_2 _18372_ (.A1(_07779_),
    .A2(_07786_),
    .A3(_07788_),
    .B1(_07789_),
    .B2(_07802_),
    .X(_08237_));
 sky130_fd_sc_hd__o21a_1 _18373_ (.A1(_01901_),
    .A2(_02152_),
    .B1(_07874_),
    .X(_08238_));
 sky130_fd_sc_hd__o31a_2 _18374_ (.A1(_01901_),
    .A2(_02152_),
    .A3(_07875_),
    .B1(_07874_),
    .X(_08239_));
 sky130_fd_sc_hd__a21oi_2 _18375_ (.A1(_07498_),
    .A2(_07794_),
    .B1(_07799_),
    .Y(_08240_));
 sky130_fd_sc_hd__a31o_1 _18376_ (.A1(_07796_),
    .A2(net48),
    .A3(net5),
    .B1(_07797_),
    .X(_08241_));
 sky130_fd_sc_hd__o31a_1 _18377_ (.A1(_01956_),
    .A2(_02109_),
    .A3(_07795_),
    .B1(_07798_),
    .X(_08242_));
 sky130_fd_sc_hd__nor2_1 _18378_ (.A(_01923_),
    .B(_02152_),
    .Y(_08244_));
 sky130_fd_sc_hd__a22oi_4 _18379_ (.A1(net5),
    .A2(net49),
    .B1(net50),
    .B2(net4),
    .Y(_08245_));
 sky130_fd_sc_hd__a22o_1 _18380_ (.A1(net5),
    .A2(net49),
    .B1(net50),
    .B2(net4),
    .X(_08246_));
 sky130_fd_sc_hd__and4_2 _18381_ (.A(net4),
    .B(net5),
    .C(net49),
    .D(net50),
    .X(_08247_));
 sky130_fd_sc_hd__nand4_4 _18382_ (.A(net4),
    .B(net5),
    .C(net49),
    .D(net50),
    .Y(_08248_));
 sky130_fd_sc_hd__o211ai_2 _18383_ (.A1(_01923_),
    .A2(_02152_),
    .B1(_08246_),
    .C1(_08248_),
    .Y(_08249_));
 sky130_fd_sc_hd__o21ai_2 _18384_ (.A1(_08245_),
    .A2(_08247_),
    .B1(_08244_),
    .Y(_08250_));
 sky130_fd_sc_hd__nand4_4 _18385_ (.A(_08246_),
    .B(_08248_),
    .C(net3),
    .D(net51),
    .Y(_08251_));
 sky130_fd_sc_hd__o22ai_4 _18386_ (.A1(_01923_),
    .A2(_02152_),
    .B1(_08245_),
    .B2(_08247_),
    .Y(_08252_));
 sky130_fd_sc_hd__o211a_2 _18387_ (.A1(_07797_),
    .A2(_08240_),
    .B1(_08251_),
    .C1(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__o211ai_4 _18388_ (.A1(_07797_),
    .A2(_08240_),
    .B1(_08251_),
    .C1(_08252_),
    .Y(_08255_));
 sky130_fd_sc_hd__a21oi_4 _18389_ (.A1(_08251_),
    .A2(_08252_),
    .B1(_08241_),
    .Y(_08256_));
 sky130_fd_sc_hd__nand3_1 _18390_ (.A(_08242_),
    .B(_08249_),
    .C(_08250_),
    .Y(_08257_));
 sky130_fd_sc_hd__a31oi_4 _18391_ (.A1(_08242_),
    .A2(_08249_),
    .A3(_08250_),
    .B1(_08239_),
    .Y(_08258_));
 sky130_fd_sc_hd__nor3_2 _18392_ (.A(_08239_),
    .B(_08253_),
    .C(_08256_),
    .Y(_08259_));
 sky130_fd_sc_hd__nand2_2 _18393_ (.A(_08258_),
    .B(_08255_),
    .Y(_08260_));
 sky130_fd_sc_hd__a2bb2oi_4 _18394_ (.A1_N(_07875_),
    .A2_N(_08238_),
    .B1(_08255_),
    .B2(_08257_),
    .Y(_08261_));
 sky130_fd_sc_hd__o22ai_4 _18395_ (.A1(_07875_),
    .A2(_08238_),
    .B1(_08253_),
    .B2(_08256_),
    .Y(_08262_));
 sky130_fd_sc_hd__a21oi_1 _18396_ (.A1(_08255_),
    .A2(_08258_),
    .B1(_08261_),
    .Y(_08263_));
 sky130_fd_sc_hd__a221oi_4 _18397_ (.A1(_08258_),
    .A2(_08255_),
    .B1(_07808_),
    .B2(_07791_),
    .C1(_08261_),
    .Y(_08264_));
 sky130_fd_sc_hd__nand3_4 _18398_ (.A(_08237_),
    .B(_08260_),
    .C(_08262_),
    .Y(_08266_));
 sky130_fd_sc_hd__a21oi_4 _18399_ (.A1(_08260_),
    .A2(_08262_),
    .B1(_08237_),
    .Y(_08267_));
 sky130_fd_sc_hd__o221ai_4 _18400_ (.A1(_07790_),
    .A2(_07787_),
    .B1(_08261_),
    .B2(_08259_),
    .C1(_07808_),
    .Y(_08268_));
 sky130_fd_sc_hd__o22ai_4 _18401_ (.A1(_07882_),
    .A2(_08235_),
    .B1(_08264_),
    .B2(_08267_),
    .Y(_08269_));
 sky130_fd_sc_hd__o22ai_2 _18402_ (.A1(_07884_),
    .A2(_07889_),
    .B1(_08237_),
    .B2(_08263_),
    .Y(_08270_));
 sky130_fd_sc_hd__o211ai_4 _18403_ (.A1(_07884_),
    .A2(_07889_),
    .B1(_08266_),
    .C1(_08268_),
    .Y(_08271_));
 sky130_fd_sc_hd__o22ai_4 _18404_ (.A1(_07884_),
    .A2(_07889_),
    .B1(_08264_),
    .B2(_08267_),
    .Y(_08272_));
 sky130_fd_sc_hd__o211ai_4 _18405_ (.A1(_07882_),
    .A2(_08235_),
    .B1(_08266_),
    .C1(_08268_),
    .Y(_08273_));
 sky130_fd_sc_hd__a22oi_4 _18406_ (.A1(_07896_),
    .A2(_08233_),
    .B1(_08269_),
    .B2(_08271_),
    .Y(_08274_));
 sky130_fd_sc_hd__nand4_4 _18407_ (.A(_07897_),
    .B(_07900_),
    .C(_08272_),
    .D(_08273_),
    .Y(_08275_));
 sky130_fd_sc_hd__a21oi_2 _18408_ (.A1(_08272_),
    .A2(_08273_),
    .B1(_08234_),
    .Y(_08277_));
 sky130_fd_sc_hd__nand4_4 _18409_ (.A(_07896_),
    .B(_08233_),
    .C(_08269_),
    .D(_08271_),
    .Y(_08278_));
 sky130_fd_sc_hd__o211a_1 _18410_ (.A1(_08229_),
    .A2(_08230_),
    .B1(_08275_),
    .C1(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__o2111ai_4 _18411_ (.A1(_08227_),
    .A2(_08224_),
    .B1(_08226_),
    .C1(_08275_),
    .D1(_08278_),
    .Y(_08280_));
 sky130_fd_sc_hd__o22ai_2 _18412_ (.A1(_08225_),
    .A2(_08228_),
    .B1(_08274_),
    .B2(_08277_),
    .Y(_08281_));
 sky130_fd_sc_hd__nand3_1 _18413_ (.A(_08231_),
    .B(_08275_),
    .C(_08278_),
    .Y(_08282_));
 sky130_fd_sc_hd__o22ai_2 _18414_ (.A1(_08229_),
    .A2(_08230_),
    .B1(_08274_),
    .B2(_08277_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand3_4 _18415_ (.A(_08281_),
    .B(_08200_),
    .C(_08280_),
    .Y(_08284_));
 sky130_fd_sc_hd__o211ai_4 _18416_ (.A1(_07846_),
    .A2(_08198_),
    .B1(_08282_),
    .C1(_08283_),
    .Y(_08285_));
 sky130_fd_sc_hd__inv_2 _18417_ (.A(_08285_),
    .Y(_08286_));
 sky130_fd_sc_hd__o21a_1 _18418_ (.A1(_07937_),
    .A2(_07940_),
    .B1(_07906_),
    .X(_08288_));
 sky130_fd_sc_hd__o21ai_1 _18419_ (.A1(_07905_),
    .A2(_07941_),
    .B1(_07906_),
    .Y(_08289_));
 sky130_fd_sc_hd__a22oi_1 _18420_ (.A1(_07906_),
    .A2(_07943_),
    .B1(_08284_),
    .B2(_08285_),
    .Y(_08290_));
 sky130_fd_sc_hd__a22o_1 _18421_ (.A1(_07906_),
    .A2(_07943_),
    .B1(_08284_),
    .B2(_08285_),
    .X(_08291_));
 sky130_fd_sc_hd__o211a_1 _18422_ (.A1(_07905_),
    .A2(_08288_),
    .B1(_08285_),
    .C1(_08284_),
    .X(_08292_));
 sky130_fd_sc_hd__o2111ai_2 _18423_ (.A1(_07905_),
    .A2(_07941_),
    .B1(_08284_),
    .C1(_08285_),
    .D1(_07906_),
    .Y(_08293_));
 sky130_fd_sc_hd__o2bb2a_1 _18424_ (.A1_N(_08284_),
    .A2_N(_08285_),
    .B1(_08288_),
    .B2(_07905_),
    .X(_08294_));
 sky130_fd_sc_hd__o2bb2ai_2 _18425_ (.A1_N(_08284_),
    .A2_N(_08285_),
    .B1(_08288_),
    .B2(_07905_),
    .Y(_08295_));
 sky130_fd_sc_hd__and3_1 _18426_ (.A(_08289_),
    .B(_08285_),
    .C(_08284_),
    .X(_08296_));
 sky130_fd_sc_hd__nand3_2 _18427_ (.A(_08289_),
    .B(_08285_),
    .C(_08284_),
    .Y(_08297_));
 sky130_fd_sc_hd__nand4_2 _18428_ (.A(_08195_),
    .B(_08197_),
    .C(_08291_),
    .D(_08293_),
    .Y(_08299_));
 sky130_fd_sc_hd__o2bb2ai_1 _18429_ (.A1_N(_08195_),
    .A2_N(_08197_),
    .B1(_08290_),
    .B2(_08292_),
    .Y(_08300_));
 sky130_fd_sc_hd__o2bb2ai_2 _18430_ (.A1_N(_08195_),
    .A2_N(_08197_),
    .B1(_08294_),
    .B2(_08296_),
    .Y(_08301_));
 sky130_fd_sc_hd__nand4_2 _18431_ (.A(_08195_),
    .B(_08197_),
    .C(_08295_),
    .D(_08297_),
    .Y(_08302_));
 sky130_fd_sc_hd__a2bb2oi_2 _18432_ (.A1_N(_07864_),
    .A2_N(_07996_),
    .B1(_08299_),
    .B2(_08300_),
    .Y(_08303_));
 sky130_fd_sc_hd__o211ai_2 _18433_ (.A1(_07864_),
    .A2(_07996_),
    .B1(_08301_),
    .C1(_08302_),
    .Y(_08304_));
 sky130_fd_sc_hd__a22oi_4 _18434_ (.A1(_07866_),
    .A2(_07995_),
    .B1(_08301_),
    .B2(_08302_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand3_2 _18435_ (.A(_07997_),
    .B(_08299_),
    .C(_08300_),
    .Y(_08306_));
 sky130_fd_sc_hd__o211a_1 _18436_ (.A1(_07569_),
    .A2(_07603_),
    .B1(_07606_),
    .C1(_07950_),
    .X(_08307_));
 sky130_fd_sc_hd__o22ai_1 _18437_ (.A1(_07951_),
    .A2(_07955_),
    .B1(_08303_),
    .B2(_08305_),
    .Y(_08308_));
 sky130_fd_sc_hd__o2111ai_1 _18438_ (.A1(_07954_),
    .A2(_07949_),
    .B1(_07950_),
    .C1(_08304_),
    .D1(_08306_),
    .Y(_08310_));
 sky130_fd_sc_hd__o2bb2ai_1 _18439_ (.A1_N(_08304_),
    .A2_N(_08306_),
    .B1(_08307_),
    .B2(_07949_),
    .Y(_08311_));
 sky130_fd_sc_hd__o21ai_1 _18440_ (.A1(_07951_),
    .A2(_07955_),
    .B1(_08306_),
    .Y(_08312_));
 sky130_fd_sc_hd__nand3_2 _18441_ (.A(_07994_),
    .B(_08308_),
    .C(_08310_),
    .Y(_08313_));
 sky130_fd_sc_hd__o211ai_4 _18442_ (.A1(_08303_),
    .A2(_08312_),
    .B1(_08311_),
    .C1(_07993_),
    .Y(_08314_));
 sky130_fd_sc_hd__a21o_1 _18443_ (.A1(_07553_),
    .A2(_07931_),
    .B1(_07932_),
    .X(_08315_));
 sky130_fd_sc_hd__a21o_1 _18444_ (.A1(_08313_),
    .A2(_08314_),
    .B1(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__nand3_2 _18445_ (.A(_08313_),
    .B(_08314_),
    .C(_08315_),
    .Y(_08317_));
 sky130_fd_sc_hd__a22o_1 _18446_ (.A1(_07933_),
    .A2(_07939_),
    .B1(_08313_),
    .B2(_08314_),
    .X(_08318_));
 sky130_fd_sc_hd__nand4_1 _18447_ (.A(_07933_),
    .B(_07939_),
    .C(_08313_),
    .D(_08314_),
    .Y(_08319_));
 sky130_fd_sc_hd__a31o_1 _18448_ (.A1(_07973_),
    .A2(_07662_),
    .A3(_07972_),
    .B1(_07978_),
    .X(_08321_));
 sky130_fd_sc_hd__nand4_1 _18449_ (.A(_07977_),
    .B(_07981_),
    .C(_08318_),
    .D(_08319_),
    .Y(_08322_));
 sky130_fd_sc_hd__nand4_2 _18450_ (.A(_07976_),
    .B(_08316_),
    .C(_08317_),
    .D(_08321_),
    .Y(_08323_));
 sky130_fd_sc_hd__and2_1 _18451_ (.A(_08322_),
    .B(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__nand2_1 _18452_ (.A(_07992_),
    .B(_07985_),
    .Y(_08325_));
 sky130_fd_sc_hd__nand2_1 _18453_ (.A(_07984_),
    .B(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__xnor2_1 _18454_ (.A(_08324_),
    .B(_08326_),
    .Y(net95));
 sky130_fd_sc_hd__a22oi_2 _18455_ (.A1(_08003_),
    .A2(_08092_),
    .B1(_08187_),
    .B2(_08190_),
    .Y(_08327_));
 sky130_fd_sc_hd__a31oi_2 _18456_ (.A1(_08095_),
    .A2(_08183_),
    .A3(_08185_),
    .B1(_08093_),
    .Y(_08328_));
 sky130_fd_sc_hd__a31o_1 _18457_ (.A1(_08013_),
    .A2(net22),
    .A3(net63),
    .B1(_08014_),
    .X(_08329_));
 sky130_fd_sc_hd__o31a_1 _18458_ (.A1(_01890_),
    .A2(_02196_),
    .A3(_08011_),
    .B1(_08015_),
    .X(_08331_));
 sky130_fd_sc_hd__o21ai_4 _18459_ (.A1(net61),
    .A2(net62),
    .B1(net25),
    .Y(_08332_));
 sky130_fd_sc_hd__o21a_2 _18460_ (.A1(net61),
    .A2(net62),
    .B1(net25),
    .X(_08333_));
 sky130_fd_sc_hd__and3_4 _18461_ (.A(net61),
    .B(net62),
    .C(net25),
    .X(_08334_));
 sky130_fd_sc_hd__nand3_4 _18462_ (.A(net61),
    .B(net62),
    .C(net25),
    .Y(_08335_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(net63),
    .B(net24),
    .Y(_08336_));
 sky130_fd_sc_hd__o211ai_4 _18464_ (.A1(_01890_),
    .A2(_02218_),
    .B1(_08333_),
    .C1(_08335_),
    .Y(_08337_));
 sky130_fd_sc_hd__o21bai_2 _18465_ (.A1(_08332_),
    .A2(_08334_),
    .B1_N(_08336_),
    .Y(_08338_));
 sky130_fd_sc_hd__nand4_2 _18466_ (.A(_08333_),
    .B(_08335_),
    .C(net63),
    .D(net24),
    .Y(_08339_));
 sky130_fd_sc_hd__o22ai_2 _18467_ (.A1(_01890_),
    .A2(_02218_),
    .B1(_08332_),
    .B2(_08334_),
    .Y(_08340_));
 sky130_fd_sc_hd__and3_2 _18468_ (.A(_08340_),
    .B(_07698_),
    .C(_08339_),
    .X(_08342_));
 sky130_fd_sc_hd__o2111ai_4 _18469_ (.A1(net60),
    .A2(_07133_),
    .B1(_07389_),
    .C1(_08339_),
    .D1(_08340_),
    .Y(_08343_));
 sky130_fd_sc_hd__nand3_2 _18470_ (.A(_07699_),
    .B(_08337_),
    .C(_08338_),
    .Y(_08344_));
 sky130_fd_sc_hd__a31oi_4 _18471_ (.A1(_07699_),
    .A2(_08337_),
    .A3(_08338_),
    .B1(_08331_),
    .Y(_08345_));
 sky130_fd_sc_hd__nand3_1 _18472_ (.A(_08344_),
    .B(_08329_),
    .C(_08343_),
    .Y(_08346_));
 sky130_fd_sc_hd__a21oi_1 _18473_ (.A1(_08343_),
    .A2(_08344_),
    .B1(_08329_),
    .Y(_08347_));
 sky130_fd_sc_hd__a21o_1 _18474_ (.A1(_08343_),
    .A2(_08344_),
    .B1(_08329_),
    .X(_08348_));
 sky130_fd_sc_hd__o2111a_1 _18475_ (.A1(_08010_),
    .A2(_08011_),
    .B1(_08015_),
    .C1(_08343_),
    .D1(_08344_),
    .X(_08349_));
 sky130_fd_sc_hd__a21oi_1 _18476_ (.A1(_08343_),
    .A2(_08344_),
    .B1(_08331_),
    .Y(_08350_));
 sky130_fd_sc_hd__a21oi_1 _18477_ (.A1(_08343_),
    .A2(_08345_),
    .B1(_08347_),
    .Y(_08351_));
 sky130_fd_sc_hd__o21ai_1 _18478_ (.A1(_06880_),
    .A2(_07682_),
    .B1(_08346_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand3_4 _18479_ (.A(_08348_),
    .B(_08008_),
    .C(_08346_),
    .Y(_08354_));
 sky130_fd_sc_hd__o31ai_4 _18480_ (.A1(_08008_),
    .A2(_08349_),
    .A3(_08350_),
    .B1(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__a31oi_4 _18481_ (.A1(_08027_),
    .A2(_08030_),
    .A3(_08008_),
    .B1(_08006_),
    .Y(_08356_));
 sky130_fd_sc_hd__a31o_1 _18482_ (.A1(_08027_),
    .A2(_08030_),
    .A3(_08008_),
    .B1(_08006_),
    .X(_08357_));
 sky130_fd_sc_hd__o311a_2 _18483_ (.A1(_06881_),
    .A2(_07676_),
    .A3(_07678_),
    .B1(_08032_),
    .C1(_08355_),
    .X(_08358_));
 sky130_fd_sc_hd__nand2_2 _18484_ (.A(_08355_),
    .B(_08356_),
    .Y(_08359_));
 sky130_fd_sc_hd__o211ai_4 _18485_ (.A1(_08008_),
    .A2(_08351_),
    .B1(_08354_),
    .C1(_08357_),
    .Y(_08360_));
 sky130_fd_sc_hd__a21boi_2 _18486_ (.A1(_08020_),
    .A2(_08024_),
    .B1_N(_08022_),
    .Y(_08361_));
 sky130_fd_sc_hd__o21ai_4 _18487_ (.A1(_08041_),
    .A2(_08044_),
    .B1(_08043_),
    .Y(_08362_));
 sky130_fd_sc_hd__nand2_2 _18488_ (.A(net35),
    .B(net20),
    .Y(_08364_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(net64),
    .B(net22),
    .Y(_08365_));
 sky130_fd_sc_hd__a22oi_4 _18490_ (.A1(net34),
    .A2(net21),
    .B1(net22),
    .B2(net64),
    .Y(_08366_));
 sky130_fd_sc_hd__a22o_1 _18491_ (.A1(net34),
    .A2(net21),
    .B1(net22),
    .B2(net64),
    .X(_08367_));
 sky130_fd_sc_hd__and4_2 _18492_ (.A(net64),
    .B(net34),
    .C(net21),
    .D(net22),
    .X(_08368_));
 sky130_fd_sc_hd__nand4_4 _18493_ (.A(net64),
    .B(net34),
    .C(net21),
    .D(net22),
    .Y(_08369_));
 sky130_fd_sc_hd__o211ai_2 _18494_ (.A1(_01934_),
    .A2(_02163_),
    .B1(_08367_),
    .C1(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__o21bai_1 _18495_ (.A1(_08366_),
    .A2(_08368_),
    .B1_N(_08364_),
    .Y(_08371_));
 sky130_fd_sc_hd__nand4_4 _18496_ (.A(_08367_),
    .B(_08369_),
    .C(net35),
    .D(net20),
    .Y(_08372_));
 sky130_fd_sc_hd__o21ai_4 _18497_ (.A1(_08366_),
    .A2(_08368_),
    .B1(_08364_),
    .Y(_08373_));
 sky130_fd_sc_hd__nand3_4 _18498_ (.A(_08373_),
    .B(_08362_),
    .C(_08372_),
    .Y(_08375_));
 sky130_fd_sc_hd__nand3b_4 _18499_ (.A_N(_08362_),
    .B(_08370_),
    .C(_08371_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand2_1 _18500_ (.A(net38),
    .B(net17),
    .Y(_08377_));
 sky130_fd_sc_hd__and4_2 _18501_ (.A(net36),
    .B(net37),
    .C(net18),
    .D(net19),
    .X(_08378_));
 sky130_fd_sc_hd__nand4_4 _18502_ (.A(net36),
    .B(net37),
    .C(net18),
    .D(net19),
    .Y(_08379_));
 sky130_fd_sc_hd__a22oi_4 _18503_ (.A1(net37),
    .A2(net18),
    .B1(net19),
    .B2(net36),
    .Y(_08380_));
 sky130_fd_sc_hd__a22o_1 _18504_ (.A1(net37),
    .A2(net18),
    .B1(net19),
    .B2(net36),
    .X(_08381_));
 sky130_fd_sc_hd__and3_1 _18505_ (.A(_08377_),
    .B(_08379_),
    .C(_08381_),
    .X(_08382_));
 sky130_fd_sc_hd__o211a_1 _18506_ (.A1(_08378_),
    .A2(_08380_),
    .B1(net38),
    .C1(net17),
    .X(_08383_));
 sky130_fd_sc_hd__a22oi_4 _18507_ (.A1(net38),
    .A2(net17),
    .B1(_08379_),
    .B2(_08381_),
    .Y(_08384_));
 sky130_fd_sc_hd__and4_1 _18508_ (.A(_08381_),
    .B(net17),
    .C(net38),
    .D(_08379_),
    .X(_08386_));
 sky130_fd_sc_hd__nor2_1 _18509_ (.A(_08384_),
    .B(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__o2bb2ai_2 _18510_ (.A1_N(_08375_),
    .A2_N(_08376_),
    .B1(_08382_),
    .B2(_08383_),
    .Y(_08388_));
 sky130_fd_sc_hd__o211ai_4 _18511_ (.A1(_08384_),
    .A2(_08386_),
    .B1(_08375_),
    .C1(_08376_),
    .Y(_08389_));
 sky130_fd_sc_hd__o2bb2ai_2 _18512_ (.A1_N(_08375_),
    .A2_N(_08376_),
    .B1(_08384_),
    .B2(_08386_),
    .Y(_08390_));
 sky130_fd_sc_hd__o211ai_2 _18513_ (.A1(_08382_),
    .A2(_08383_),
    .B1(_08375_),
    .C1(_08376_),
    .Y(_08391_));
 sky130_fd_sc_hd__nand3_2 _18514_ (.A(_08361_),
    .B(_08388_),
    .C(_08389_),
    .Y(_08392_));
 sky130_fd_sc_hd__o211a_2 _18515_ (.A1(_08021_),
    .A2(_08028_),
    .B1(_08390_),
    .C1(_08391_),
    .X(_08393_));
 sky130_fd_sc_hd__o211ai_4 _18516_ (.A1(_08021_),
    .A2(_08028_),
    .B1(_08390_),
    .C1(_08391_),
    .Y(_08394_));
 sky130_fd_sc_hd__a21oi_2 _18517_ (.A1(_08050_),
    .A2(_08061_),
    .B1(_08062_),
    .Y(_08395_));
 sky130_fd_sc_hd__a22oi_4 _18518_ (.A1(_08050_),
    .A2(_08064_),
    .B1(_08392_),
    .B2(_08394_),
    .Y(_08397_));
 sky130_fd_sc_hd__a22o_1 _18519_ (.A1(_08050_),
    .A2(_08064_),
    .B1(_08392_),
    .B2(_08394_),
    .X(_08398_));
 sky130_fd_sc_hd__a31oi_4 _18520_ (.A1(_08361_),
    .A2(_08388_),
    .A3(_08389_),
    .B1(_08395_),
    .Y(_08399_));
 sky130_fd_sc_hd__and3b_1 _18521_ (.A_N(_08395_),
    .B(_08394_),
    .C(_08392_),
    .X(_08400_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(_08399_),
    .B(_08394_),
    .Y(_08401_));
 sky130_fd_sc_hd__o2bb2ai_4 _18523_ (.A1_N(_08359_),
    .A2_N(_08360_),
    .B1(_08397_),
    .B2(_08400_),
    .Y(_08402_));
 sky130_fd_sc_hd__nand4_4 _18524_ (.A(_08359_),
    .B(_08360_),
    .C(_08398_),
    .D(_08401_),
    .Y(_08403_));
 sky130_fd_sc_hd__a21boi_1 _18525_ (.A1(_08082_),
    .A2(_08085_),
    .B1_N(_08038_),
    .Y(_08404_));
 sky130_fd_sc_hd__a31oi_4 _18526_ (.A1(_08038_),
    .A2(_08079_),
    .A3(_08080_),
    .B1(_08036_),
    .Y(_08405_));
 sky130_fd_sc_hd__a21oi_4 _18527_ (.A1(_08402_),
    .A2(_08403_),
    .B1(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__o2bb2ai_2 _18528_ (.A1_N(_08402_),
    .A2_N(_08403_),
    .B1(_08404_),
    .B2(_08036_),
    .Y(_08408_));
 sky130_fd_sc_hd__nand3_4 _18529_ (.A(_08405_),
    .B(_08403_),
    .C(_08402_),
    .Y(_08409_));
 sky130_fd_sc_hd__nand2_1 _18530_ (.A(_08408_),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__o21ai_2 _18531_ (.A1(_08051_),
    .A2(_08052_),
    .B1(_08055_),
    .Y(_08411_));
 sky130_fd_sc_hd__o22a_1 _18532_ (.A1(_07741_),
    .A2(_08054_),
    .B1(_08051_),
    .B2(_08052_),
    .X(_08412_));
 sky130_fd_sc_hd__nor2_1 _18533_ (.A(_02010_),
    .B(_02065_),
    .Y(_08413_));
 sky130_fd_sc_hd__a22oi_4 _18534_ (.A1(net40),
    .A2(net15),
    .B1(net16),
    .B2(net39),
    .Y(_08414_));
 sky130_fd_sc_hd__a22o_1 _18535_ (.A1(net40),
    .A2(net15),
    .B1(net16),
    .B2(net39),
    .X(_08415_));
 sky130_fd_sc_hd__and4_1 _18536_ (.A(net39),
    .B(net40),
    .C(net15),
    .D(net16),
    .X(_08416_));
 sky130_fd_sc_hd__nand4_4 _18537_ (.A(net39),
    .B(net40),
    .C(net15),
    .D(net16),
    .Y(_08417_));
 sky130_fd_sc_hd__o211ai_4 _18538_ (.A1(_02010_),
    .A2(_02065_),
    .B1(_08415_),
    .C1(_08417_),
    .Y(_08419_));
 sky130_fd_sc_hd__o21ai_2 _18539_ (.A1(_08414_),
    .A2(_08416_),
    .B1(_08413_),
    .Y(_08420_));
 sky130_fd_sc_hd__a22o_1 _18540_ (.A1(net41),
    .A2(net14),
    .B1(_08415_),
    .B2(_08417_),
    .X(_08421_));
 sky130_fd_sc_hd__nand4_2 _18541_ (.A(_08415_),
    .B(_08417_),
    .C(net41),
    .D(net14),
    .Y(_08422_));
 sky130_fd_sc_hd__nand3_4 _18542_ (.A(_08412_),
    .B(_08419_),
    .C(_08420_),
    .Y(_08423_));
 sky130_fd_sc_hd__and3_1 _18543_ (.A(_08421_),
    .B(_08422_),
    .C(_08411_),
    .X(_08424_));
 sky130_fd_sc_hd__nand3_4 _18544_ (.A(_08421_),
    .B(_08422_),
    .C(_08411_),
    .Y(_08425_));
 sky130_fd_sc_hd__o21a_1 _18545_ (.A1(_02010_),
    .A2(_02043_),
    .B1(_08151_),
    .X(_08426_));
 sky130_fd_sc_hd__and3_1 _18546_ (.A(_08149_),
    .B(net13),
    .C(net41),
    .X(_08427_));
 sky130_fd_sc_hd__o31a_1 _18547_ (.A1(_02010_),
    .A2(_02043_),
    .A3(_08148_),
    .B1(_08151_),
    .X(_08428_));
 sky130_fd_sc_hd__a31oi_2 _18548_ (.A1(_08412_),
    .A2(_08419_),
    .A3(_08420_),
    .B1(_08428_),
    .Y(_08430_));
 sky130_fd_sc_hd__o211ai_2 _18549_ (.A1(_08150_),
    .A2(_08427_),
    .B1(_08425_),
    .C1(_08423_),
    .Y(_08431_));
 sky130_fd_sc_hd__o2bb2ai_1 _18550_ (.A1_N(_08423_),
    .A2_N(_08425_),
    .B1(_08426_),
    .B2(_08148_),
    .Y(_08432_));
 sky130_fd_sc_hd__o2bb2ai_2 _18551_ (.A1_N(_08423_),
    .A2_N(_08425_),
    .B1(_08427_),
    .B2(_08150_),
    .Y(_08433_));
 sky130_fd_sc_hd__o2111ai_4 _18552_ (.A1(_08147_),
    .A2(_08148_),
    .B1(_08151_),
    .C1(_08423_),
    .D1(_08425_),
    .Y(_08434_));
 sky130_fd_sc_hd__a21oi_1 _18553_ (.A1(_08159_),
    .A2(_08142_),
    .B1(_08157_),
    .Y(_08435_));
 sky130_fd_sc_hd__and3_2 _18554_ (.A(_08433_),
    .B(_08435_),
    .C(_08434_),
    .X(_08436_));
 sky130_fd_sc_hd__nand3_4 _18555_ (.A(_08433_),
    .B(_08435_),
    .C(_08434_),
    .Y(_08437_));
 sky130_fd_sc_hd__o211ai_4 _18556_ (.A1(_08157_),
    .A2(_08160_),
    .B1(_08431_),
    .C1(_08432_),
    .Y(_08438_));
 sky130_fd_sc_hd__o21ai_1 _18557_ (.A1(_07781_),
    .A2(_08102_),
    .B1(_08101_),
    .Y(_08439_));
 sky130_fd_sc_hd__a21oi_1 _18558_ (.A1(_07781_),
    .A2(_08102_),
    .B1(_08101_),
    .Y(_08441_));
 sky130_fd_sc_hd__nand2_1 _18559_ (.A(net43),
    .B(net13),
    .Y(_08442_));
 sky130_fd_sc_hd__and4_1 _18560_ (.A(net42),
    .B(net11),
    .C(net43),
    .D(net13),
    .X(_08443_));
 sky130_fd_sc_hd__nand4_1 _18561_ (.A(net42),
    .B(net11),
    .C(net43),
    .D(net13),
    .Y(_08444_));
 sky130_fd_sc_hd__a22o_2 _18562_ (.A1(net11),
    .A2(net43),
    .B1(net13),
    .B2(net42),
    .X(_08445_));
 sky130_fd_sc_hd__a2bb2oi_1 _18563_ (.A1_N(_02021_),
    .A2_N(_02054_),
    .B1(_08444_),
    .B2(_08445_),
    .Y(_08446_));
 sky130_fd_sc_hd__o2bb2ai_2 _18564_ (.A1_N(_08444_),
    .A2_N(_08445_),
    .B1(_02021_),
    .B2(_02054_),
    .Y(_08447_));
 sky130_fd_sc_hd__o2111a_2 _18565_ (.A1(_08102_),
    .A2(_08442_),
    .B1(net10),
    .C1(net45),
    .D1(_08445_),
    .X(_08448_));
 sky130_fd_sc_hd__o2111ai_4 _18566_ (.A1(_08102_),
    .A2(_08442_),
    .B1(net10),
    .C1(net45),
    .D1(_08445_),
    .Y(_08449_));
 sky130_fd_sc_hd__a22oi_2 _18567_ (.A1(_08106_),
    .A2(_08439_),
    .B1(_08447_),
    .B2(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__o2bb2ai_2 _18568_ (.A1_N(_08106_),
    .A2_N(_08439_),
    .B1(_08446_),
    .B2(_08448_),
    .Y(_08452_));
 sky130_fd_sc_hd__o21ai_2 _18569_ (.A1(_08103_),
    .A2(_08441_),
    .B1(_08447_),
    .Y(_08453_));
 sky130_fd_sc_hd__o211ai_2 _18570_ (.A1(_08103_),
    .A2(_08441_),
    .B1(_08447_),
    .C1(_08449_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand2_1 _18571_ (.A(net9),
    .B(net46),
    .Y(_08455_));
 sky130_fd_sc_hd__a22oi_1 _18572_ (.A1(net9),
    .A2(net46),
    .B1(net47),
    .B2(net8),
    .Y(_08456_));
 sky130_fd_sc_hd__nand2_1 _18573_ (.A(_08120_),
    .B(_08455_),
    .Y(_08457_));
 sky130_fd_sc_hd__nand2_2 _18574_ (.A(net9),
    .B(net47),
    .Y(_08458_));
 sky130_fd_sc_hd__nand4_2 _18575_ (.A(net8),
    .B(net9),
    .C(net46),
    .D(net47),
    .Y(_08459_));
 sky130_fd_sc_hd__nand2_1 _18576_ (.A(net7),
    .B(net48),
    .Y(_08460_));
 sky130_fd_sc_hd__a22oi_2 _18577_ (.A1(net7),
    .A2(net48),
    .B1(_08457_),
    .B2(_08459_),
    .Y(_08461_));
 sky130_fd_sc_hd__a22o_1 _18578_ (.A1(net7),
    .A2(net48),
    .B1(_08457_),
    .B2(_08459_),
    .X(_08463_));
 sky130_fd_sc_hd__o2111a_1 _18579_ (.A1(_08117_),
    .A2(_08458_),
    .B1(net7),
    .C1(net48),
    .D1(_08457_),
    .X(_08464_));
 sky130_fd_sc_hd__o2111ai_1 _18580_ (.A1(_08117_),
    .A2(_08458_),
    .B1(net7),
    .C1(net48),
    .D1(_08457_),
    .Y(_08465_));
 sky130_fd_sc_hd__nor2_1 _18581_ (.A(_08461_),
    .B(_08464_),
    .Y(_08466_));
 sky130_fd_sc_hd__nand2_1 _18582_ (.A(_08463_),
    .B(_08465_),
    .Y(_08467_));
 sky130_fd_sc_hd__a21oi_2 _18583_ (.A1(_08452_),
    .A2(_08454_),
    .B1(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__o221a_2 _18584_ (.A1(_08461_),
    .A2(_08464_),
    .B1(_08448_),
    .B2(_08453_),
    .C1(_08452_),
    .X(_08469_));
 sky130_fd_sc_hd__o2bb2a_1 _18585_ (.A1_N(_08452_),
    .A2_N(_08454_),
    .B1(_08461_),
    .B2(_08464_),
    .X(_08470_));
 sky130_fd_sc_hd__and3_1 _18586_ (.A(_08452_),
    .B(_08466_),
    .C(_08454_),
    .X(_08471_));
 sky130_fd_sc_hd__nor2_2 _18587_ (.A(_08468_),
    .B(_08469_),
    .Y(_08472_));
 sky130_fd_sc_hd__o2bb2ai_1 _18588_ (.A1_N(_08437_),
    .A2_N(_08438_),
    .B1(_08470_),
    .B2(_08471_),
    .Y(_08474_));
 sky130_fd_sc_hd__o211ai_2 _18589_ (.A1(_08468_),
    .A2(_08469_),
    .B1(_08437_),
    .C1(_08438_),
    .Y(_08475_));
 sky130_fd_sc_hd__o211ai_4 _18590_ (.A1(_08470_),
    .A2(_08471_),
    .B1(_08437_),
    .C1(_08438_),
    .Y(_08476_));
 sky130_fd_sc_hd__o2bb2ai_2 _18591_ (.A1_N(_08437_),
    .A2_N(_08438_),
    .B1(_08468_),
    .B2(_08469_),
    .Y(_08477_));
 sky130_fd_sc_hd__a31oi_4 _18592_ (.A1(_08068_),
    .A2(_08070_),
    .A3(_08069_),
    .B1(_08077_),
    .Y(_08478_));
 sky130_fd_sc_hd__a32oi_4 _18593_ (.A1(_08065_),
    .A2(_08066_),
    .A3(_08071_),
    .B1(_08074_),
    .B2(_08076_),
    .Y(_08479_));
 sky130_fd_sc_hd__o211a_1 _18594_ (.A1(_08072_),
    .A2(_08478_),
    .B1(_08477_),
    .C1(_08476_),
    .X(_08480_));
 sky130_fd_sc_hd__o211ai_4 _18595_ (.A1(_08072_),
    .A2(_08478_),
    .B1(_08477_),
    .C1(_08476_),
    .Y(_08481_));
 sky130_fd_sc_hd__nand3_4 _18596_ (.A(_08479_),
    .B(_08475_),
    .C(_08474_),
    .Y(_08482_));
 sky130_fd_sc_hd__o32a_2 _18597_ (.A1(_08162_),
    .A2(_08163_),
    .A3(_08139_),
    .B1(_08136_),
    .B2(_08134_),
    .X(_08483_));
 sky130_fd_sc_hd__o31a_1 _18598_ (.A1(_08131_),
    .A2(_08132_),
    .A3(_08165_),
    .B1(_08169_),
    .X(_08485_));
 sky130_fd_sc_hd__o31a_1 _18599_ (.A1(_08139_),
    .A2(_08162_),
    .A3(_08163_),
    .B1(_08170_),
    .X(_08486_));
 sky130_fd_sc_hd__o2bb2ai_2 _18600_ (.A1_N(_08481_),
    .A2_N(_08482_),
    .B1(_08483_),
    .B2(_08168_),
    .Y(_08487_));
 sky130_fd_sc_hd__nand3_2 _18601_ (.A(_08481_),
    .B(_08485_),
    .C(_08482_),
    .Y(_08488_));
 sky130_fd_sc_hd__a21oi_1 _18602_ (.A1(_08481_),
    .A2(_08482_),
    .B1(_08486_),
    .Y(_08489_));
 sky130_fd_sc_hd__a22o_1 _18603_ (.A1(_08167_),
    .A2(_08170_),
    .B1(_08481_),
    .B2(_08482_),
    .X(_08490_));
 sky130_fd_sc_hd__o211a_1 _18604_ (.A1(_08168_),
    .A2(_08483_),
    .B1(_08482_),
    .C1(_08481_),
    .X(_08491_));
 sky130_fd_sc_hd__o211ai_2 _18605_ (.A1(_08168_),
    .A2(_08483_),
    .B1(_08482_),
    .C1(_08481_),
    .Y(_08492_));
 sky130_fd_sc_hd__nand2_1 _18606_ (.A(_08487_),
    .B(_08488_),
    .Y(_08493_));
 sky130_fd_sc_hd__nand4_2 _18607_ (.A(_08408_),
    .B(_08409_),
    .C(_08490_),
    .D(_08492_),
    .Y(_08494_));
 sky130_fd_sc_hd__o2bb2ai_1 _18608_ (.A1_N(_08408_),
    .A2_N(_08409_),
    .B1(_08489_),
    .B2(_08491_),
    .Y(_08496_));
 sky130_fd_sc_hd__nand2_1 _18609_ (.A(_08410_),
    .B(_08493_),
    .Y(_08497_));
 sky130_fd_sc_hd__o21ai_1 _18610_ (.A1(_08489_),
    .A2(_08491_),
    .B1(_08409_),
    .Y(_08498_));
 sky130_fd_sc_hd__o221ai_4 _18611_ (.A1(_08406_),
    .A2(_08498_),
    .B1(_08093_),
    .B2(_08327_),
    .C1(_08497_),
    .Y(_08499_));
 sky130_fd_sc_hd__nand3_4 _18612_ (.A(_08328_),
    .B(_08494_),
    .C(_08496_),
    .Y(_08500_));
 sky130_fd_sc_hd__o21ai_2 _18613_ (.A1(_08225_),
    .A2(_08228_),
    .B1(_08278_),
    .Y(_08501_));
 sky130_fd_sc_hd__o21a_1 _18614_ (.A1(_08274_),
    .A2(_08231_),
    .B1(_08278_),
    .X(_08502_));
 sky130_fd_sc_hd__o21ai_2 _18615_ (.A1(_08181_),
    .A2(_08175_),
    .B1(_08179_),
    .Y(_08503_));
 sky130_fd_sc_hd__a21oi_2 _18616_ (.A1(_08176_),
    .A2(_08180_),
    .B1(_08178_),
    .Y(_08504_));
 sky130_fd_sc_hd__o21ai_1 _18617_ (.A1(_08203_),
    .A2(_08204_),
    .B1(_08206_),
    .Y(_08505_));
 sky130_fd_sc_hd__o21a_1 _18618_ (.A1(_08203_),
    .A2(_08204_),
    .B1(_08206_),
    .X(_08507_));
 sky130_fd_sc_hd__nand2_1 _18619_ (.A(net32),
    .B(net54),
    .Y(_08508_));
 sky130_fd_sc_hd__nand2_1 _18620_ (.A(net3),
    .B(net52),
    .Y(_08509_));
 sky130_fd_sc_hd__a22oi_1 _18621_ (.A1(net3),
    .A2(net52),
    .B1(net53),
    .B2(net2),
    .Y(_08510_));
 sky130_fd_sc_hd__a22o_1 _18622_ (.A1(net3),
    .A2(net52),
    .B1(net53),
    .B2(net2),
    .X(_08511_));
 sky130_fd_sc_hd__and4_1 _18623_ (.A(net2),
    .B(net3),
    .C(net52),
    .D(net53),
    .X(_08512_));
 sky130_fd_sc_hd__nand4_1 _18624_ (.A(net2),
    .B(net3),
    .C(net52),
    .D(net53),
    .Y(_08513_));
 sky130_fd_sc_hd__o211ai_1 _18625_ (.A1(_01912_),
    .A2(_02207_),
    .B1(_08511_),
    .C1(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__o21bai_1 _18626_ (.A1(_08510_),
    .A2(_08512_),
    .B1_N(_08508_),
    .Y(_08515_));
 sky130_fd_sc_hd__nand4_1 _18627_ (.A(_08511_),
    .B(_08513_),
    .C(net32),
    .D(net54),
    .Y(_08516_));
 sky130_fd_sc_hd__o21ai_1 _18628_ (.A1(_08510_),
    .A2(_08512_),
    .B1(_08508_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand3_2 _18629_ (.A(_08518_),
    .B(_08505_),
    .C(_08516_),
    .Y(_08519_));
 sky130_fd_sc_hd__nand3_2 _18630_ (.A(_08507_),
    .B(_08514_),
    .C(_08515_),
    .Y(_08520_));
 sky130_fd_sc_hd__and4_2 _18631_ (.A(_01868_),
    .B(net31),
    .C(net56),
    .D(net57),
    .X(_08521_));
 sky130_fd_sc_hd__o22a_1 _18632_ (.A1(net30),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01879_),
    .X(_08522_));
 sky130_fd_sc_hd__o211a_1 _18633_ (.A1(_01879_),
    .A2(_02229_),
    .B1(net57),
    .C1(_01868_),
    .X(_08523_));
 sky130_fd_sc_hd__o211a_1 _18634_ (.A1(net30),
    .A2(_02240_),
    .B1(net56),
    .C1(net31),
    .X(_08524_));
 sky130_fd_sc_hd__o2bb2ai_2 _18635_ (.A1_N(_08519_),
    .A2_N(_08520_),
    .B1(_08521_),
    .B2(_08522_),
    .Y(_08525_));
 sky130_fd_sc_hd__o211ai_4 _18636_ (.A1(_08523_),
    .A2(_08524_),
    .B1(_08519_),
    .C1(_08520_),
    .Y(_08526_));
 sky130_fd_sc_hd__nand2_1 _18637_ (.A(_08525_),
    .B(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__a21boi_2 _18638_ (.A1(_08212_),
    .A2(_08218_),
    .B1_N(_08213_),
    .Y(_08529_));
 sky130_fd_sc_hd__nand2_1 _18639_ (.A(_08527_),
    .B(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__nand3b_4 _18640_ (.A_N(_08529_),
    .B(_08526_),
    .C(_08525_),
    .Y(_08531_));
 sky130_fd_sc_hd__inv_2 _18641_ (.A(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__a21o_1 _18642_ (.A1(_08530_),
    .A2(_08531_),
    .B1(_08215_),
    .X(_08533_));
 sky130_fd_sc_hd__a21o_1 _18643_ (.A1(_08527_),
    .A2(_08529_),
    .B1(_08216_),
    .X(_08534_));
 sky130_fd_sc_hd__o311a_2 _18644_ (.A1(net29),
    .A2(_02240_),
    .A3(_08214_),
    .B1(_08530_),
    .C1(_08531_),
    .X(_08535_));
 sky130_fd_sc_hd__nand3_1 _18645_ (.A(_08216_),
    .B(_08530_),
    .C(_08531_),
    .Y(_08536_));
 sky130_fd_sc_hd__a21oi_2 _18646_ (.A1(_08530_),
    .A2(_08531_),
    .B1(_08216_),
    .Y(_08537_));
 sky130_fd_sc_hd__a21o_1 _18647_ (.A1(_08530_),
    .A2(_08531_),
    .B1(_08216_),
    .X(_08538_));
 sky130_fd_sc_hd__o21ai_2 _18648_ (.A1(_08534_),
    .A2(_08532_),
    .B1(_08533_),
    .Y(_08540_));
 sky130_fd_sc_hd__o21ai_4 _18649_ (.A1(_08236_),
    .A2(_08267_),
    .B1(_08266_),
    .Y(_08541_));
 sky130_fd_sc_hd__a31o_1 _18650_ (.A1(_08241_),
    .A2(_08251_),
    .A3(_08252_),
    .B1(_08258_),
    .X(_08542_));
 sky130_fd_sc_hd__o21ai_2 _18651_ (.A1(_08124_),
    .A2(_08118_),
    .B1(_08123_),
    .Y(_08543_));
 sky130_fd_sc_hd__o22a_1 _18652_ (.A1(_07794_),
    .A2(_08120_),
    .B1(_08124_),
    .B2(_08118_),
    .X(_08544_));
 sky130_fd_sc_hd__nand2_1 _18653_ (.A(net4),
    .B(net51),
    .Y(_08545_));
 sky130_fd_sc_hd__a22oi_4 _18654_ (.A1(net6),
    .A2(net49),
    .B1(net50),
    .B2(net5),
    .Y(_08546_));
 sky130_fd_sc_hd__a22o_1 _18655_ (.A1(net6),
    .A2(net49),
    .B1(net50),
    .B2(net5),
    .X(_08547_));
 sky130_fd_sc_hd__and4_1 _18656_ (.A(net5),
    .B(net6),
    .C(net49),
    .D(net50),
    .X(_08548_));
 sky130_fd_sc_hd__nand4_4 _18657_ (.A(net5),
    .B(net6),
    .C(net49),
    .D(net50),
    .Y(_08549_));
 sky130_fd_sc_hd__o211ai_2 _18658_ (.A1(_01945_),
    .A2(_02152_),
    .B1(_08547_),
    .C1(_08549_),
    .Y(_08551_));
 sky130_fd_sc_hd__o21bai_2 _18659_ (.A1(_08546_),
    .A2(_08548_),
    .B1_N(_08545_),
    .Y(_08552_));
 sky130_fd_sc_hd__a22o_1 _18660_ (.A1(net4),
    .A2(net51),
    .B1(_08547_),
    .B2(_08549_),
    .X(_08553_));
 sky130_fd_sc_hd__nand4_2 _18661_ (.A(_08547_),
    .B(_08549_),
    .C(net4),
    .D(net51),
    .Y(_08554_));
 sky130_fd_sc_hd__and3_2 _18662_ (.A(_08544_),
    .B(_08551_),
    .C(_08552_),
    .X(_08555_));
 sky130_fd_sc_hd__nand3_4 _18663_ (.A(_08544_),
    .B(_08551_),
    .C(_08552_),
    .Y(_08556_));
 sky130_fd_sc_hd__nand3_4 _18664_ (.A(_08553_),
    .B(_08554_),
    .C(_08543_),
    .Y(_08557_));
 sky130_fd_sc_hd__o21a_1 _18665_ (.A1(_01923_),
    .A2(_02152_),
    .B1(_08248_),
    .X(_08558_));
 sky130_fd_sc_hd__and3_1 _18666_ (.A(_08246_),
    .B(net51),
    .C(net3),
    .X(_08559_));
 sky130_fd_sc_hd__o31a_1 _18667_ (.A1(_01923_),
    .A2(_02152_),
    .A3(_08245_),
    .B1(_08248_),
    .X(_08560_));
 sky130_fd_sc_hd__o2bb2ai_2 _18668_ (.A1_N(_08556_),
    .A2_N(_08557_),
    .B1(_08558_),
    .B2(_08245_),
    .Y(_08562_));
 sky130_fd_sc_hd__o211a_2 _18669_ (.A1(_08247_),
    .A2(_08559_),
    .B1(_08557_),
    .C1(_08556_),
    .X(_08563_));
 sky130_fd_sc_hd__o211ai_2 _18670_ (.A1(_08247_),
    .A2(_08559_),
    .B1(_08557_),
    .C1(_08556_),
    .Y(_08564_));
 sky130_fd_sc_hd__o2bb2ai_1 _18671_ (.A1_N(_08556_),
    .A2_N(_08557_),
    .B1(_08559_),
    .B2(_08247_),
    .Y(_08565_));
 sky130_fd_sc_hd__o211ai_2 _18672_ (.A1(_08245_),
    .A2(_08558_),
    .B1(_08557_),
    .C1(_08556_),
    .Y(_08566_));
 sky130_fd_sc_hd__a2bb2oi_1 _18673_ (.A1_N(_08110_),
    .A2_N(_08114_),
    .B1(_08129_),
    .B2(_08113_),
    .Y(_08567_));
 sky130_fd_sc_hd__nand3_4 _18674_ (.A(_08567_),
    .B(_08566_),
    .C(_08565_),
    .Y(_08568_));
 sky130_fd_sc_hd__o21ai_4 _18675_ (.A1(_08115_),
    .A2(_08135_),
    .B1(_08562_),
    .Y(_08569_));
 sky130_fd_sc_hd__o211ai_4 _18676_ (.A1(_08115_),
    .A2(_08135_),
    .B1(_08562_),
    .C1(_08564_),
    .Y(_08570_));
 sky130_fd_sc_hd__a21o_1 _18677_ (.A1(_08568_),
    .A2(_08570_),
    .B1(_08542_),
    .X(_08571_));
 sky130_fd_sc_hd__o221ai_4 _18678_ (.A1(_08253_),
    .A2(_08259_),
    .B1(_08563_),
    .B2(_08569_),
    .C1(_08568_),
    .Y(_08573_));
 sky130_fd_sc_hd__a22o_1 _18679_ (.A1(_08255_),
    .A2(_08260_),
    .B1(_08568_),
    .B2(_08570_),
    .X(_08574_));
 sky130_fd_sc_hd__o2111ai_4 _18680_ (.A1(_08256_),
    .A2(_08239_),
    .B1(_08255_),
    .C1(_08568_),
    .D1(_08570_),
    .Y(_08575_));
 sky130_fd_sc_hd__a22oi_4 _18681_ (.A1(_08266_),
    .A2(_08270_),
    .B1(_08574_),
    .B2(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand3_4 _18682_ (.A(_08541_),
    .B(_08571_),
    .C(_08573_),
    .Y(_08577_));
 sky130_fd_sc_hd__a21oi_4 _18683_ (.A1(_08571_),
    .A2(_08573_),
    .B1(_08541_),
    .Y(_08578_));
 sky130_fd_sc_hd__o2111ai_4 _18684_ (.A1(_08267_),
    .A2(_08236_),
    .B1(_08266_),
    .C1(_08574_),
    .D1(_08575_),
    .Y(_08579_));
 sky130_fd_sc_hd__nand4_2 _18685_ (.A(_08536_),
    .B(_08538_),
    .C(_08577_),
    .D(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__o22ai_4 _18686_ (.A1(_08535_),
    .A2(_08537_),
    .B1(_08576_),
    .B2(_08578_),
    .Y(_08581_));
 sky130_fd_sc_hd__o211a_2 _18687_ (.A1(_08534_),
    .A2(_08532_),
    .B1(_08533_),
    .C1(_08579_),
    .X(_08582_));
 sky130_fd_sc_hd__o21ai_2 _18688_ (.A1(_08535_),
    .A2(_08537_),
    .B1(_08579_),
    .Y(_08584_));
 sky130_fd_sc_hd__o21ai_2 _18689_ (.A1(_08576_),
    .A2(_08578_),
    .B1(_08540_),
    .Y(_08585_));
 sky130_fd_sc_hd__o211a_1 _18690_ (.A1(_08576_),
    .A2(_08584_),
    .B1(_08503_),
    .C1(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__o211ai_4 _18691_ (.A1(_08576_),
    .A2(_08584_),
    .B1(_08503_),
    .C1(_08585_),
    .Y(_08587_));
 sky130_fd_sc_hd__and3_1 _18692_ (.A(_08504_),
    .B(_08580_),
    .C(_08581_),
    .X(_08588_));
 sky130_fd_sc_hd__nand3_4 _18693_ (.A(_08504_),
    .B(_08580_),
    .C(_08581_),
    .Y(_08589_));
 sky130_fd_sc_hd__a22oi_4 _18694_ (.A1(_08275_),
    .A2(_08501_),
    .B1(_08587_),
    .B2(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__a22o_1 _18695_ (.A1(_08275_),
    .A2(_08501_),
    .B1(_08587_),
    .B2(_08589_),
    .X(_08591_));
 sky130_fd_sc_hd__a31o_1 _18696_ (.A1(_08504_),
    .A2(_08580_),
    .A3(_08581_),
    .B1(_08502_),
    .X(_08592_));
 sky130_fd_sc_hd__inv_2 _18697_ (.A(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__o211a_1 _18698_ (.A1(_08277_),
    .A2(_08279_),
    .B1(_08587_),
    .C1(_08589_),
    .X(_08595_));
 sky130_fd_sc_hd__o211ai_2 _18699_ (.A1(_08277_),
    .A2(_08279_),
    .B1(_08587_),
    .C1(_08589_),
    .Y(_08596_));
 sky130_fd_sc_hd__a21oi_1 _18700_ (.A1(_08587_),
    .A2(_08589_),
    .B1(_08502_),
    .Y(_08597_));
 sky130_fd_sc_hd__and3_1 _18701_ (.A(_08502_),
    .B(_08587_),
    .C(_08589_),
    .X(_08598_));
 sky130_fd_sc_hd__o211ai_2 _18702_ (.A1(_08590_),
    .A2(_08595_),
    .B1(_08499_),
    .C1(_08500_),
    .Y(_08599_));
 sky130_fd_sc_hd__o2bb2ai_1 _18703_ (.A1_N(_08499_),
    .A2_N(_08500_),
    .B1(_08597_),
    .B2(_08598_),
    .Y(_08600_));
 sky130_fd_sc_hd__o2bb2a_2 _18704_ (.A1_N(_08499_),
    .A2_N(_08500_),
    .B1(_08590_),
    .B2(_08595_),
    .X(_08601_));
 sky130_fd_sc_hd__o2bb2ai_1 _18705_ (.A1_N(_08499_),
    .A2_N(_08500_),
    .B1(_08590_),
    .B2(_08595_),
    .Y(_08602_));
 sky130_fd_sc_hd__nand4_2 _18706_ (.A(_08499_),
    .B(_08500_),
    .C(_08591_),
    .D(_08596_),
    .Y(_08603_));
 sky130_fd_sc_hd__a32oi_4 _18707_ (.A1(_08000_),
    .A2(_08193_),
    .A3(_08194_),
    .B1(_08295_),
    .B2(_08297_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand3_1 _18708_ (.A(_08195_),
    .B(_08291_),
    .C(_08293_),
    .Y(_08606_));
 sky130_fd_sc_hd__o211ai_4 _18709_ (.A1(_08196_),
    .A2(_08604_),
    .B1(_08600_),
    .C1(_08599_),
    .Y(_08607_));
 sky130_fd_sc_hd__nand3_2 _18710_ (.A(_08197_),
    .B(_08603_),
    .C(_08606_),
    .Y(_08608_));
 sky130_fd_sc_hd__nand4_2 _18711_ (.A(_08197_),
    .B(_08602_),
    .C(_08603_),
    .D(_08606_),
    .Y(_08609_));
 sky130_fd_sc_hd__and3_1 _18712_ (.A(_07906_),
    .B(_07943_),
    .C(_08284_),
    .X(_08610_));
 sky130_fd_sc_hd__a31o_1 _18713_ (.A1(_08200_),
    .A2(_08280_),
    .A3(_08281_),
    .B1(_08296_),
    .X(_08611_));
 sky130_fd_sc_hd__o211ai_4 _18714_ (.A1(_08601_),
    .A2(_08608_),
    .B1(_08611_),
    .C1(_08607_),
    .Y(_08612_));
 sky130_fd_sc_hd__o2bb2ai_4 _18715_ (.A1_N(_08607_),
    .A2_N(_08609_),
    .B1(_08610_),
    .B2(_08286_),
    .Y(_08613_));
 sky130_fd_sc_hd__o211a_1 _18716_ (.A1(_07954_),
    .A2(_07949_),
    .B1(_07950_),
    .C1(_08304_),
    .X(_08614_));
 sky130_fd_sc_hd__o21ai_1 _18717_ (.A1(_07949_),
    .A2(_08307_),
    .B1(_08304_),
    .Y(_08615_));
 sky130_fd_sc_hd__o2bb2ai_4 _18718_ (.A1_N(_08612_),
    .A2_N(_08613_),
    .B1(_08614_),
    .B2(_08305_),
    .Y(_08617_));
 sky130_fd_sc_hd__nand4_4 _18719_ (.A(_08306_),
    .B(_08612_),
    .C(_08613_),
    .D(_08615_),
    .Y(_08618_));
 sky130_fd_sc_hd__o31a_1 _18720_ (.A1(_08201_),
    .A2(_08219_),
    .A3(_08220_),
    .B1(_08227_),
    .X(_08619_));
 sky130_fd_sc_hd__a21o_1 _18721_ (.A1(_08617_),
    .A2(_08618_),
    .B1(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__nand3_1 _18722_ (.A(_08617_),
    .B(_08618_),
    .C(_08619_),
    .Y(_08621_));
 sky130_fd_sc_hd__a21bo_1 _18723_ (.A1(_08617_),
    .A2(_08618_),
    .B1_N(_08619_),
    .X(_08622_));
 sky130_fd_sc_hd__o2111ai_4 _18724_ (.A1(_07911_),
    .A2(_08224_),
    .B1(_08617_),
    .C1(_08618_),
    .D1(_08223_),
    .Y(_08623_));
 sky130_fd_sc_hd__nand2_1 _18725_ (.A(_08314_),
    .B(_08317_),
    .Y(_08624_));
 sky130_fd_sc_hd__nand4_1 _18726_ (.A(_08314_),
    .B(_08317_),
    .C(_08620_),
    .D(_08621_),
    .Y(_08625_));
 sky130_fd_sc_hd__nand3_1 _18727_ (.A(_08624_),
    .B(_08623_),
    .C(_08622_),
    .Y(_08626_));
 sky130_fd_sc_hd__inv_2 _18728_ (.A(_08626_),
    .Y(_08628_));
 sky130_fd_sc_hd__and2_1 _18729_ (.A(_08625_),
    .B(_08626_),
    .X(_08629_));
 sky130_fd_sc_hd__a21boi_2 _18730_ (.A1(_07985_),
    .A2(_08323_),
    .B1_N(_08322_),
    .Y(_08630_));
 sky130_fd_sc_hd__nand4_1 _18731_ (.A(_07984_),
    .B(_07985_),
    .C(_08322_),
    .D(_08323_),
    .Y(_08631_));
 sky130_fd_sc_hd__o21bai_1 _18732_ (.A1(_08631_),
    .A2(_07992_),
    .B1_N(_08630_),
    .Y(_08632_));
 sky130_fd_sc_hd__xor2_1 _18733_ (.A(_08629_),
    .B(_08632_),
    .X(net96));
 sky130_fd_sc_hd__a21o_1 _18734_ (.A1(_08632_),
    .A2(_08629_),
    .B1(_08628_),
    .X(_08633_));
 sky130_fd_sc_hd__o21ai_2 _18735_ (.A1(_08590_),
    .A2(_08595_),
    .B1(_08499_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand3_2 _18736_ (.A(_08500_),
    .B(_08591_),
    .C(_08596_),
    .Y(_08635_));
 sky130_fd_sc_hd__a32oi_4 _18737_ (.A1(_08405_),
    .A2(_08403_),
    .A3(_08402_),
    .B1(_08488_),
    .B2(_08487_),
    .Y(_08636_));
 sky130_fd_sc_hd__o21ai_1 _18738_ (.A1(_08489_),
    .A2(_08491_),
    .B1(_08408_),
    .Y(_08638_));
 sky130_fd_sc_hd__a31oi_2 _18739_ (.A1(_08409_),
    .A2(_08490_),
    .A3(_08492_),
    .B1(_08406_),
    .Y(_08639_));
 sky130_fd_sc_hd__a2bb2oi_2 _18740_ (.A1_N(_08356_),
    .A2_N(_08355_),
    .B1(_08401_),
    .B2(_08398_),
    .Y(_08640_));
 sky130_fd_sc_hd__o22ai_2 _18741_ (.A1(_08355_),
    .A2(_08356_),
    .B1(_08397_),
    .B2(_08400_),
    .Y(_08641_));
 sky130_fd_sc_hd__o21ai_2 _18742_ (.A1(_08347_),
    .A2(_08353_),
    .B1(_08007_),
    .Y(_08642_));
 sky130_fd_sc_hd__a22oi_4 _18743_ (.A1(net63),
    .A2(net25),
    .B1(_08333_),
    .B2(_08335_),
    .Y(_08643_));
 sky130_fd_sc_hd__o22ai_4 _18744_ (.A1(_01890_),
    .A2(_02251_),
    .B1(_08332_),
    .B2(_08334_),
    .Y(_08644_));
 sky130_fd_sc_hd__o211a_1 _18745_ (.A1(net61),
    .A2(net62),
    .B1(net63),
    .C1(net25),
    .X(_08645_));
 sky130_fd_sc_hd__o211ai_4 _18746_ (.A1(net61),
    .A2(net62),
    .B1(net63),
    .C1(net25),
    .Y(_08646_));
 sky130_fd_sc_hd__o2111a_4 _18747_ (.A1(net61),
    .A2(net62),
    .B1(net63),
    .C1(net25),
    .D1(_08335_),
    .X(_08647_));
 sky130_fd_sc_hd__o2111ai_4 _18748_ (.A1(net61),
    .A2(net62),
    .B1(net63),
    .C1(net25),
    .D1(_08335_),
    .Y(_08649_));
 sky130_fd_sc_hd__a21oi_2 _18749_ (.A1(_08335_),
    .A2(_08645_),
    .B1(_08643_),
    .Y(_08650_));
 sky130_fd_sc_hd__a22oi_4 _18750_ (.A1(_07389_),
    .A2(_07697_),
    .B1(_08644_),
    .B2(_08649_),
    .Y(_08651_));
 sky130_fd_sc_hd__o22ai_4 _18751_ (.A1(_07387_),
    .A2(_07696_),
    .B1(_08643_),
    .B2(_08647_),
    .Y(_08652_));
 sky130_fd_sc_hd__nand2_4 _18752_ (.A(_08644_),
    .B(_07698_),
    .Y(_08653_));
 sky130_fd_sc_hd__o211a_4 _18753_ (.A1(_08334_),
    .A2(_08646_),
    .B1(_07698_),
    .C1(_08644_),
    .X(_08654_));
 sky130_fd_sc_hd__o2111ai_2 _18754_ (.A1(net60),
    .A2(_07133_),
    .B1(_07389_),
    .C1(_08644_),
    .D1(_08649_),
    .Y(_08655_));
 sky130_fd_sc_hd__a31o_2 _18755_ (.A1(_08333_),
    .A2(net24),
    .A3(net63),
    .B1(_08334_),
    .X(_08656_));
 sky130_fd_sc_hd__o31a_1 _18756_ (.A1(_01890_),
    .A2(_02218_),
    .A3(_08332_),
    .B1(_08335_),
    .X(_08657_));
 sky130_fd_sc_hd__o21ai_1 _18757_ (.A1(_08651_),
    .A2(_08654_),
    .B1(_08656_),
    .Y(_08658_));
 sky130_fd_sc_hd__o2111ai_2 _18758_ (.A1(_08336_),
    .A2(_08332_),
    .B1(_08335_),
    .C1(_08652_),
    .D1(_08655_),
    .Y(_08660_));
 sky130_fd_sc_hd__o21ai_2 _18759_ (.A1(_08651_),
    .A2(_08654_),
    .B1(_08657_),
    .Y(_08661_));
 sky130_fd_sc_hd__o211ai_4 _18760_ (.A1(_08647_),
    .A2(_08653_),
    .B1(_08656_),
    .C1(_08652_),
    .Y(_08662_));
 sky130_fd_sc_hd__nand3_1 _18761_ (.A(_08009_),
    .B(_08661_),
    .C(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__nand3_1 _18762_ (.A(_08658_),
    .B(_08660_),
    .C(_08008_),
    .Y(_08664_));
 sky130_fd_sc_hd__nand3_1 _18763_ (.A(_08009_),
    .B(_08658_),
    .C(_08660_),
    .Y(_08665_));
 sky130_fd_sc_hd__o2111ai_4 _18764_ (.A1(_06880_),
    .A2(_07682_),
    .B1(_08007_),
    .C1(_08661_),
    .D1(_08662_),
    .Y(_08666_));
 sky130_fd_sc_hd__nand4_4 _18765_ (.A(_08007_),
    .B(_08354_),
    .C(_08663_),
    .D(_08664_),
    .Y(_08667_));
 sky130_fd_sc_hd__and3_1 _18766_ (.A(_08642_),
    .B(_08665_),
    .C(_08666_),
    .X(_08668_));
 sky130_fd_sc_hd__nand3_4 _18767_ (.A(_08642_),
    .B(_08665_),
    .C(_08666_),
    .Y(_08669_));
 sky130_fd_sc_hd__and2_1 _18768_ (.A(net38),
    .B(net18),
    .X(_08671_));
 sky130_fd_sc_hd__a22oi_4 _18769_ (.A1(net37),
    .A2(net19),
    .B1(net20),
    .B2(net36),
    .Y(_08672_));
 sky130_fd_sc_hd__a22o_1 _18770_ (.A1(net37),
    .A2(net19),
    .B1(net20),
    .B2(net36),
    .X(_08673_));
 sky130_fd_sc_hd__and4_2 _18771_ (.A(net36),
    .B(net37),
    .C(net19),
    .D(net20),
    .X(_08674_));
 sky130_fd_sc_hd__a211oi_4 _18772_ (.A1(net38),
    .A2(net18),
    .B1(_08672_),
    .C1(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__o211a_1 _18773_ (.A1(_08672_),
    .A2(_08674_),
    .B1(net38),
    .C1(net18),
    .X(_08676_));
 sky130_fd_sc_hd__o2bb2a_1 _18774_ (.A1_N(net38),
    .A2_N(net18),
    .B1(_08672_),
    .B2(_08674_),
    .X(_08677_));
 sky130_fd_sc_hd__and4b_1 _18775_ (.A_N(_08674_),
    .B(net18),
    .C(net38),
    .D(_08673_),
    .X(_08678_));
 sky130_fd_sc_hd__a21oi_2 _18776_ (.A1(_08042_),
    .A2(_08365_),
    .B1(_08364_),
    .Y(_08679_));
 sky130_fd_sc_hd__a31o_1 _18777_ (.A1(_08367_),
    .A2(net20),
    .A3(net35),
    .B1(_08368_),
    .X(_08680_));
 sky130_fd_sc_hd__o31a_1 _18778_ (.A1(_01934_),
    .A2(_02163_),
    .A3(_08366_),
    .B1(_08369_),
    .X(_08682_));
 sky130_fd_sc_hd__nand2_1 _18779_ (.A(net35),
    .B(net21),
    .Y(_08683_));
 sky130_fd_sc_hd__a22oi_4 _18780_ (.A1(net34),
    .A2(net22),
    .B1(net24),
    .B2(net64),
    .Y(_08684_));
 sky130_fd_sc_hd__a22o_1 _18781_ (.A1(net34),
    .A2(net22),
    .B1(net24),
    .B2(net64),
    .X(_08685_));
 sky130_fd_sc_hd__and4_2 _18782_ (.A(net64),
    .B(net34),
    .C(net22),
    .D(net24),
    .X(_08686_));
 sky130_fd_sc_hd__nand4_4 _18783_ (.A(net64),
    .B(net34),
    .C(net22),
    .D(net24),
    .Y(_08687_));
 sky130_fd_sc_hd__o211ai_1 _18784_ (.A1(_01934_),
    .A2(_02185_),
    .B1(_08685_),
    .C1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__a21o_1 _18785_ (.A1(_08685_),
    .A2(_08687_),
    .B1(_08683_),
    .X(_08689_));
 sky130_fd_sc_hd__nand4_4 _18786_ (.A(_08685_),
    .B(_08687_),
    .C(net35),
    .D(net21),
    .Y(_08690_));
 sky130_fd_sc_hd__o22ai_4 _18787_ (.A1(_01934_),
    .A2(_02185_),
    .B1(_08684_),
    .B2(_08686_),
    .Y(_08691_));
 sky130_fd_sc_hd__o211a_2 _18788_ (.A1(_08368_),
    .A2(_08679_),
    .B1(_08690_),
    .C1(_08691_),
    .X(_08693_));
 sky130_fd_sc_hd__o211ai_4 _18789_ (.A1(_08368_),
    .A2(_08679_),
    .B1(_08690_),
    .C1(_08691_),
    .Y(_08694_));
 sky130_fd_sc_hd__a21oi_2 _18790_ (.A1(_08690_),
    .A2(_08691_),
    .B1(_08680_),
    .Y(_08695_));
 sky130_fd_sc_hd__nand3_2 _18791_ (.A(_08682_),
    .B(_08688_),
    .C(_08689_),
    .Y(_08696_));
 sky130_fd_sc_hd__o22ai_4 _18792_ (.A1(_08675_),
    .A2(_08676_),
    .B1(_08693_),
    .B2(_08695_),
    .Y(_08697_));
 sky130_fd_sc_hd__o211ai_4 _18793_ (.A1(_08677_),
    .A2(_08678_),
    .B1(_08694_),
    .C1(_08696_),
    .Y(_08698_));
 sky130_fd_sc_hd__o21ai_4 _18794_ (.A1(_08675_),
    .A2(_08676_),
    .B1(_08696_),
    .Y(_08699_));
 sky130_fd_sc_hd__o22ai_2 _18795_ (.A1(_08677_),
    .A2(_08678_),
    .B1(_08693_),
    .B2(_08695_),
    .Y(_08700_));
 sky130_fd_sc_hd__a21oi_2 _18796_ (.A1(_08329_),
    .A2(_08344_),
    .B1(_08342_),
    .Y(_08701_));
 sky130_fd_sc_hd__nand3_4 _18797_ (.A(_08697_),
    .B(_08698_),
    .C(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__o221a_2 _18798_ (.A1(_08342_),
    .A2(_08345_),
    .B1(_08693_),
    .B2(_08699_),
    .C1(_08700_),
    .X(_08703_));
 sky130_fd_sc_hd__o221ai_4 _18799_ (.A1(_08342_),
    .A2(_08345_),
    .B1(_08693_),
    .B2(_08699_),
    .C1(_08700_),
    .Y(_08704_));
 sky130_fd_sc_hd__a32oi_4 _18800_ (.A1(_08362_),
    .A2(_08372_),
    .A3(_08373_),
    .B1(_08376_),
    .B2(_08387_),
    .Y(_08705_));
 sky130_fd_sc_hd__a32o_2 _18801_ (.A1(_08362_),
    .A2(_08372_),
    .A3(_08373_),
    .B1(_08376_),
    .B2(_08387_),
    .X(_08706_));
 sky130_fd_sc_hd__a21oi_1 _18802_ (.A1(_08702_),
    .A2(_08704_),
    .B1(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__a21o_2 _18803_ (.A1(_08702_),
    .A2(_08704_),
    .B1(_08706_),
    .X(_08708_));
 sky130_fd_sc_hd__a31oi_2 _18804_ (.A1(_08697_),
    .A2(_08698_),
    .A3(_08701_),
    .B1(_08705_),
    .Y(_08709_));
 sky130_fd_sc_hd__a31o_1 _18805_ (.A1(_08697_),
    .A2(_08698_),
    .A3(_08701_),
    .B1(_08705_),
    .X(_08710_));
 sky130_fd_sc_hd__and3_1 _18806_ (.A(_08702_),
    .B(_08704_),
    .C(_08706_),
    .X(_08711_));
 sky130_fd_sc_hd__nand3_2 _18807_ (.A(_08702_),
    .B(_08704_),
    .C(_08706_),
    .Y(_08712_));
 sky130_fd_sc_hd__a22oi_4 _18808_ (.A1(_08667_),
    .A2(_08669_),
    .B1(_08708_),
    .B2(_08712_),
    .Y(_08714_));
 sky130_fd_sc_hd__o2bb2ai_1 _18809_ (.A1_N(_08667_),
    .A2_N(_08669_),
    .B1(_08707_),
    .B2(_08711_),
    .Y(_08715_));
 sky130_fd_sc_hd__o2111a_2 _18810_ (.A1(_08710_),
    .A2(_08703_),
    .B1(_08669_),
    .C1(_08667_),
    .D1(_08708_),
    .X(_08716_));
 sky130_fd_sc_hd__o2111ai_4 _18811_ (.A1(_08710_),
    .A2(_08703_),
    .B1(_08669_),
    .C1(_08667_),
    .D1(_08708_),
    .Y(_08717_));
 sky130_fd_sc_hd__nand4_4 _18812_ (.A(_08359_),
    .B(_08641_),
    .C(_08715_),
    .D(_08717_),
    .Y(_08718_));
 sky130_fd_sc_hd__o22ai_4 _18813_ (.A1(_08358_),
    .A2(_08640_),
    .B1(_08714_),
    .B2(_08716_),
    .Y(_08719_));
 sky130_fd_sc_hd__nor2_1 _18814_ (.A(_08393_),
    .B(_08399_),
    .Y(_08720_));
 sky130_fd_sc_hd__a31o_1 _18815_ (.A1(_08445_),
    .A2(net45),
    .A3(net10),
    .B1(_08443_),
    .X(_08721_));
 sky130_fd_sc_hd__nand2_1 _18816_ (.A(net11),
    .B(net45),
    .Y(_08722_));
 sky130_fd_sc_hd__nand2_1 _18817_ (.A(net43),
    .B(net14),
    .Y(_08723_));
 sky130_fd_sc_hd__nand4_2 _18818_ (.A(net42),
    .B(net43),
    .C(net13),
    .D(net14),
    .Y(_08725_));
 sky130_fd_sc_hd__a22oi_1 _18819_ (.A1(net43),
    .A2(net13),
    .B1(net14),
    .B2(net42),
    .Y(_08726_));
 sky130_fd_sc_hd__a22o_1 _18820_ (.A1(net43),
    .A2(net13),
    .B1(net14),
    .B2(net42),
    .X(_08727_));
 sky130_fd_sc_hd__o2bb2ai_2 _18821_ (.A1_N(_08725_),
    .A2_N(_08727_),
    .B1(_02032_),
    .B2(_02054_),
    .Y(_08728_));
 sky130_fd_sc_hd__and4_1 _18822_ (.A(_08727_),
    .B(net45),
    .C(net11),
    .D(_08725_),
    .X(_08729_));
 sky130_fd_sc_hd__nand4_2 _18823_ (.A(_08727_),
    .B(net45),
    .C(net11),
    .D(_08725_),
    .Y(_08730_));
 sky130_fd_sc_hd__a21oi_2 _18824_ (.A1(_08728_),
    .A2(_08730_),
    .B1(_08721_),
    .Y(_08731_));
 sky130_fd_sc_hd__a21o_1 _18825_ (.A1(_08728_),
    .A2(_08730_),
    .B1(_08721_),
    .X(_08732_));
 sky130_fd_sc_hd__nand2_1 _18826_ (.A(_08721_),
    .B(_08728_),
    .Y(_08733_));
 sky130_fd_sc_hd__nand3_1 _18827_ (.A(_08721_),
    .B(_08728_),
    .C(_08730_),
    .Y(_08734_));
 sky130_fd_sc_hd__nand2_1 _18828_ (.A(net8),
    .B(net48),
    .Y(_08736_));
 sky130_fd_sc_hd__nand2_1 _18829_ (.A(net10),
    .B(net46),
    .Y(_08737_));
 sky130_fd_sc_hd__and4_1 _18830_ (.A(net9),
    .B(net10),
    .C(net46),
    .D(net47),
    .X(_08738_));
 sky130_fd_sc_hd__nand4_1 _18831_ (.A(net9),
    .B(net10),
    .C(net46),
    .D(net47),
    .Y(_08739_));
 sky130_fd_sc_hd__a22o_1 _18832_ (.A1(net10),
    .A2(net46),
    .B1(net47),
    .B2(net9),
    .X(_08740_));
 sky130_fd_sc_hd__o211a_1 _18833_ (.A1(_01988_),
    .A2(_02109_),
    .B1(_08739_),
    .C1(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__a21oi_1 _18834_ (.A1(_08739_),
    .A2(_08740_),
    .B1(_08736_),
    .Y(_08742_));
 sky130_fd_sc_hd__nor2_2 _18835_ (.A(_08741_),
    .B(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__a21oi_2 _18836_ (.A1(_08732_),
    .A2(_08734_),
    .B1(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__and3_1 _18837_ (.A(_08732_),
    .B(_08734_),
    .C(_08743_),
    .X(_08745_));
 sky130_fd_sc_hd__a21boi_2 _18838_ (.A1(_08732_),
    .A2(_08734_),
    .B1_N(_08743_),
    .Y(_08747_));
 sky130_fd_sc_hd__o221a_2 _18839_ (.A1(_08741_),
    .A2(_08742_),
    .B1(_08729_),
    .B2(_08733_),
    .C1(_08732_),
    .X(_08748_));
 sky130_fd_sc_hd__o21ai_2 _18840_ (.A1(_08148_),
    .A2(_08426_),
    .B1(_08425_),
    .Y(_08749_));
 sky130_fd_sc_hd__o21a_1 _18841_ (.A1(_02010_),
    .A2(_02065_),
    .B1(_08417_),
    .X(_08750_));
 sky130_fd_sc_hd__o31a_1 _18842_ (.A1(_02010_),
    .A2(_02065_),
    .A3(_08414_),
    .B1(_08417_),
    .X(_08751_));
 sky130_fd_sc_hd__nor2_2 _18843_ (.A(_08377_),
    .B(_08380_),
    .Y(_08752_));
 sky130_fd_sc_hd__o21ai_2 _18844_ (.A1(_08377_),
    .A2(_08380_),
    .B1(_08379_),
    .Y(_08753_));
 sky130_fd_sc_hd__o21a_1 _18845_ (.A1(_08377_),
    .A2(_08380_),
    .B1(_08379_),
    .X(_08754_));
 sky130_fd_sc_hd__nor2_1 _18846_ (.A(_02010_),
    .B(_02076_),
    .Y(_08755_));
 sky130_fd_sc_hd__a22oi_4 _18847_ (.A1(net40),
    .A2(net16),
    .B1(net17),
    .B2(net39),
    .Y(_08756_));
 sky130_fd_sc_hd__a22o_1 _18848_ (.A1(net40),
    .A2(net16),
    .B1(net17),
    .B2(net39),
    .X(_08758_));
 sky130_fd_sc_hd__and4_1 _18849_ (.A(net39),
    .B(net40),
    .C(net16),
    .D(net17),
    .X(_08759_));
 sky130_fd_sc_hd__nand4_4 _18850_ (.A(net39),
    .B(net40),
    .C(net16),
    .D(net17),
    .Y(_08760_));
 sky130_fd_sc_hd__o211ai_2 _18851_ (.A1(_02010_),
    .A2(_02076_),
    .B1(_08758_),
    .C1(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__o21ai_1 _18852_ (.A1(_08756_),
    .A2(_08759_),
    .B1(_08755_),
    .Y(_08762_));
 sky130_fd_sc_hd__o22ai_4 _18853_ (.A1(_02010_),
    .A2(_02076_),
    .B1(_08756_),
    .B2(_08759_),
    .Y(_08763_));
 sky130_fd_sc_hd__nand4_4 _18854_ (.A(_08758_),
    .B(_08760_),
    .C(net41),
    .D(net15),
    .Y(_08764_));
 sky130_fd_sc_hd__a2bb2oi_2 _18855_ (.A1_N(_08378_),
    .A2_N(_08752_),
    .B1(_08761_),
    .B2(_08762_),
    .Y(_08765_));
 sky130_fd_sc_hd__o211ai_4 _18856_ (.A1(_08378_),
    .A2(_08752_),
    .B1(_08763_),
    .C1(_08764_),
    .Y(_08766_));
 sky130_fd_sc_hd__a21oi_2 _18857_ (.A1(_08763_),
    .A2(_08764_),
    .B1(_08753_),
    .Y(_08767_));
 sky130_fd_sc_hd__a21o_1 _18858_ (.A1(_08763_),
    .A2(_08764_),
    .B1(_08753_),
    .X(_08769_));
 sky130_fd_sc_hd__a31oi_1 _18859_ (.A1(_08754_),
    .A2(_08761_),
    .A3(_08762_),
    .B1(_08751_),
    .Y(_08770_));
 sky130_fd_sc_hd__nand3b_4 _18860_ (.A_N(_08751_),
    .B(_08766_),
    .C(_08769_),
    .Y(_08771_));
 sky130_fd_sc_hd__o22ai_4 _18861_ (.A1(_08414_),
    .A2(_08750_),
    .B1(_08765_),
    .B2(_08767_),
    .Y(_08772_));
 sky130_fd_sc_hd__o211a_1 _18862_ (.A1(_08424_),
    .A2(_08430_),
    .B1(_08771_),
    .C1(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__o211ai_4 _18863_ (.A1(_08424_),
    .A2(_08430_),
    .B1(_08771_),
    .C1(_08772_),
    .Y(_08774_));
 sky130_fd_sc_hd__a22oi_4 _18864_ (.A1(_08423_),
    .A2(_08749_),
    .B1(_08771_),
    .B2(_08772_),
    .Y(_08775_));
 sky130_fd_sc_hd__a22o_1 _18865_ (.A1(_08423_),
    .A2(_08749_),
    .B1(_08771_),
    .B2(_08772_),
    .X(_08776_));
 sky130_fd_sc_hd__o211a_1 _18866_ (.A1(_08744_),
    .A2(_08745_),
    .B1(_08774_),
    .C1(_08776_),
    .X(_08777_));
 sky130_fd_sc_hd__o211ai_2 _18867_ (.A1(_08744_),
    .A2(_08745_),
    .B1(_08774_),
    .C1(_08776_),
    .Y(_08778_));
 sky130_fd_sc_hd__o22ai_4 _18868_ (.A1(_08747_),
    .A2(_08748_),
    .B1(_08773_),
    .B2(_08775_),
    .Y(_08780_));
 sky130_fd_sc_hd__o211ai_2 _18869_ (.A1(_08747_),
    .A2(_08748_),
    .B1(_08774_),
    .C1(_08776_),
    .Y(_08781_));
 sky130_fd_sc_hd__o22ai_2 _18870_ (.A1(_08744_),
    .A2(_08745_),
    .B1(_08773_),
    .B2(_08775_),
    .Y(_08782_));
 sky130_fd_sc_hd__o21ai_2 _18871_ (.A1(_08393_),
    .A2(_08399_),
    .B1(_08780_),
    .Y(_08783_));
 sky130_fd_sc_hd__a2bb2oi_1 _18872_ (.A1_N(_08393_),
    .A2_N(_08399_),
    .B1(_08781_),
    .B2(_08782_),
    .Y(_08784_));
 sky130_fd_sc_hd__o211ai_4 _18873_ (.A1(_08393_),
    .A2(_08399_),
    .B1(_08778_),
    .C1(_08780_),
    .Y(_08785_));
 sky130_fd_sc_hd__nand3_4 _18874_ (.A(_08782_),
    .B(_08720_),
    .C(_08781_),
    .Y(_08786_));
 sky130_fd_sc_hd__o21a_1 _18875_ (.A1(_08470_),
    .A2(_08471_),
    .B1(_08438_),
    .X(_08787_));
 sky130_fd_sc_hd__o21ai_4 _18876_ (.A1(_08436_),
    .A2(_08472_),
    .B1(_08438_),
    .Y(_08788_));
 sky130_fd_sc_hd__a21boi_1 _18877_ (.A1(_08785_),
    .A2(_08786_),
    .B1_N(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__a21bo_1 _18878_ (.A1(_08785_),
    .A2(_08786_),
    .B1_N(_08788_),
    .X(_08791_));
 sky130_fd_sc_hd__o211a_1 _18879_ (.A1(_08436_),
    .A2(_08787_),
    .B1(_08786_),
    .C1(_08785_),
    .X(_08792_));
 sky130_fd_sc_hd__o2111ai_4 _18880_ (.A1(_08436_),
    .A2(_08472_),
    .B1(_08785_),
    .C1(_08786_),
    .D1(_08438_),
    .Y(_08793_));
 sky130_fd_sc_hd__a21oi_1 _18881_ (.A1(_08785_),
    .A2(_08786_),
    .B1(_08788_),
    .Y(_08794_));
 sky130_fd_sc_hd__o2bb2ai_2 _18882_ (.A1_N(_08785_),
    .A2_N(_08786_),
    .B1(_08787_),
    .B2(_08436_),
    .Y(_08795_));
 sky130_fd_sc_hd__and3_1 _18883_ (.A(_08785_),
    .B(_08786_),
    .C(_08788_),
    .X(_08796_));
 sky130_fd_sc_hd__o211ai_4 _18884_ (.A1(_08777_),
    .A2(_08783_),
    .B1(_08786_),
    .C1(_08788_),
    .Y(_08797_));
 sky130_fd_sc_hd__nand4_4 _18885_ (.A(_08718_),
    .B(_08719_),
    .C(_08791_),
    .D(_08793_),
    .Y(_08798_));
 sky130_fd_sc_hd__o2bb2ai_4 _18886_ (.A1_N(_08718_),
    .A2_N(_08719_),
    .B1(_08789_),
    .B2(_08792_),
    .Y(_08799_));
 sky130_fd_sc_hd__o2bb2ai_1 _18887_ (.A1_N(_08718_),
    .A2_N(_08719_),
    .B1(_08794_),
    .B2(_08796_),
    .Y(_08800_));
 sky130_fd_sc_hd__nand4_2 _18888_ (.A(_08718_),
    .B(_08719_),
    .C(_08795_),
    .D(_08797_),
    .Y(_08802_));
 sky130_fd_sc_hd__a22oi_4 _18889_ (.A1(_08409_),
    .A2(_08638_),
    .B1(_08798_),
    .B2(_08799_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand3_4 _18890_ (.A(_08639_),
    .B(_08800_),
    .C(_08802_),
    .Y(_08804_));
 sky130_fd_sc_hd__o211a_1 _18891_ (.A1(_08406_),
    .A2(_08636_),
    .B1(_08798_),
    .C1(_08799_),
    .X(_08805_));
 sky130_fd_sc_hd__o211ai_4 _18892_ (.A1(_08406_),
    .A2(_08636_),
    .B1(_08798_),
    .C1(_08799_),
    .Y(_08806_));
 sky130_fd_sc_hd__o21a_1 _18893_ (.A1(_08168_),
    .A2(_08483_),
    .B1(_08482_),
    .X(_08807_));
 sky130_fd_sc_hd__o21ai_1 _18894_ (.A1(_08168_),
    .A2(_08483_),
    .B1(_08482_),
    .Y(_08808_));
 sky130_fd_sc_hd__a41o_1 _18895_ (.A1(_08074_),
    .A2(_08083_),
    .A3(_08476_),
    .A4(_08477_),
    .B1(_08486_),
    .X(_08809_));
 sky130_fd_sc_hd__o21ai_2 _18896_ (.A1(_08486_),
    .A2(_08480_),
    .B1(_08482_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand2_1 _18897_ (.A(_08519_),
    .B(_08526_),
    .Y(_08811_));
 sky130_fd_sc_hd__o21ai_1 _18898_ (.A1(_01912_),
    .A2(_02207_),
    .B1(_08513_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_1 _18899_ (.A(net2),
    .B(net54),
    .Y(_08814_));
 sky130_fd_sc_hd__nand2_1 _18900_ (.A(net4),
    .B(net53),
    .Y(_08815_));
 sky130_fd_sc_hd__nand4_2 _18901_ (.A(net3),
    .B(net4),
    .C(net52),
    .D(net53),
    .Y(_08816_));
 sky130_fd_sc_hd__a22oi_1 _18902_ (.A1(net4),
    .A2(net52),
    .B1(net53),
    .B2(net3),
    .Y(_08817_));
 sky130_fd_sc_hd__a22o_1 _18903_ (.A1(net4),
    .A2(net52),
    .B1(net53),
    .B2(net3),
    .X(_08818_));
 sky130_fd_sc_hd__o2111a_1 _18904_ (.A1(_08509_),
    .A2(_08815_),
    .B1(net2),
    .C1(net54),
    .D1(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__o2111ai_4 _18905_ (.A1(_08509_),
    .A2(_08815_),
    .B1(net2),
    .C1(net54),
    .D1(_08818_),
    .Y(_08820_));
 sky130_fd_sc_hd__a22oi_1 _18906_ (.A1(net2),
    .A2(net54),
    .B1(_08816_),
    .B2(_08818_),
    .Y(_08821_));
 sky130_fd_sc_hd__o2bb2ai_1 _18907_ (.A1_N(_08816_),
    .A2_N(_08818_),
    .B1(_01901_),
    .B2(_02207_),
    .Y(_08822_));
 sky130_fd_sc_hd__nand4_1 _18908_ (.A(_08511_),
    .B(_08813_),
    .C(_08820_),
    .D(_08822_),
    .Y(_08824_));
 sky130_fd_sc_hd__a22oi_1 _18909_ (.A1(_08511_),
    .A2(_08813_),
    .B1(_08820_),
    .B2(_08822_),
    .Y(_08825_));
 sky130_fd_sc_hd__o2bb2ai_1 _18910_ (.A1_N(_08511_),
    .A2_N(_08813_),
    .B1(_08819_),
    .B2(_08821_),
    .Y(_08826_));
 sky130_fd_sc_hd__and4b_2 _18911_ (.A_N(net31),
    .B(net32),
    .C(net56),
    .D(net57),
    .X(_08827_));
 sky130_fd_sc_hd__a22oi_1 _18912_ (.A1(net32),
    .A2(net56),
    .B1(_01879_),
    .B2(net57),
    .Y(_08828_));
 sky130_fd_sc_hd__or2_1 _18913_ (.A(_08827_),
    .B(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__o2bb2ai_1 _18914_ (.A1_N(_08824_),
    .A2_N(_08826_),
    .B1(_08827_),
    .B2(_08828_),
    .Y(_08830_));
 sky130_fd_sc_hd__nand3b_1 _18915_ (.A_N(_08829_),
    .B(_08826_),
    .C(_08824_),
    .Y(_08831_));
 sky130_fd_sc_hd__a21o_1 _18916_ (.A1(_08830_),
    .A2(_08831_),
    .B1(_08811_),
    .X(_08832_));
 sky130_fd_sc_hd__nand3_2 _18917_ (.A(_08811_),
    .B(_08830_),
    .C(_08831_),
    .Y(_08833_));
 sky130_fd_sc_hd__inv_2 _18918_ (.A(_08833_),
    .Y(_08835_));
 sky130_fd_sc_hd__a21o_4 _18919_ (.A1(_08832_),
    .A2(_08833_),
    .B1(_08521_),
    .X(_08836_));
 sky130_fd_sc_hd__nand2_2 _18920_ (.A(_08832_),
    .B(_08521_),
    .Y(_08837_));
 sky130_fd_sc_hd__and3_1 _18921_ (.A(_08832_),
    .B(_08833_),
    .C(_08521_),
    .X(_08838_));
 sky130_fd_sc_hd__nand3_2 _18922_ (.A(_08832_),
    .B(_08833_),
    .C(_08521_),
    .Y(_08839_));
 sky130_fd_sc_hd__o21ai_4 _18923_ (.A1(_08835_),
    .A2(_08837_),
    .B1(_08836_),
    .Y(_08840_));
 sky130_fd_sc_hd__o21ai_1 _18924_ (.A1(_08460_),
    .A2(_08456_),
    .B1(_08459_),
    .Y(_08841_));
 sky130_fd_sc_hd__o22a_1 _18925_ (.A1(_08117_),
    .A2(_08458_),
    .B1(_08460_),
    .B2(_08456_),
    .X(_08842_));
 sky130_fd_sc_hd__nor2_1 _18926_ (.A(_01956_),
    .B(_02152_),
    .Y(_08843_));
 sky130_fd_sc_hd__a22oi_4 _18927_ (.A1(net7),
    .A2(net49),
    .B1(net50),
    .B2(net6),
    .Y(_08844_));
 sky130_fd_sc_hd__a22o_1 _18928_ (.A1(net7),
    .A2(net49),
    .B1(net50),
    .B2(net6),
    .X(_08846_));
 sky130_fd_sc_hd__and4_1 _18929_ (.A(net6),
    .B(net7),
    .C(net49),
    .D(net50),
    .X(_08847_));
 sky130_fd_sc_hd__nand4_2 _18930_ (.A(net6),
    .B(net7),
    .C(net49),
    .D(net50),
    .Y(_08848_));
 sky130_fd_sc_hd__o211ai_4 _18931_ (.A1(_01956_),
    .A2(_02152_),
    .B1(_08846_),
    .C1(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__o21ai_2 _18932_ (.A1(_08844_),
    .A2(_08847_),
    .B1(_08843_),
    .Y(_08850_));
 sky130_fd_sc_hd__o22ai_1 _18933_ (.A1(_01956_),
    .A2(_02152_),
    .B1(_08844_),
    .B2(_08847_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand4_1 _18934_ (.A(_08846_),
    .B(_08848_),
    .C(net5),
    .D(net51),
    .Y(_08852_));
 sky130_fd_sc_hd__nand3_4 _18935_ (.A(_08842_),
    .B(_08849_),
    .C(_08850_),
    .Y(_08853_));
 sky130_fd_sc_hd__and3_2 _18936_ (.A(_08851_),
    .B(_08852_),
    .C(_08841_),
    .X(_08854_));
 sky130_fd_sc_hd__nand3_2 _18937_ (.A(_08851_),
    .B(_08852_),
    .C(_08841_),
    .Y(_08855_));
 sky130_fd_sc_hd__o21a_1 _18938_ (.A1(_01945_),
    .A2(_02152_),
    .B1(_08549_),
    .X(_08857_));
 sky130_fd_sc_hd__a31o_1 _18939_ (.A1(_08547_),
    .A2(net51),
    .A3(net4),
    .B1(_08548_),
    .X(_08858_));
 sky130_fd_sc_hd__o31a_1 _18940_ (.A1(_01945_),
    .A2(_02152_),
    .A3(_08546_),
    .B1(_08549_),
    .X(_08859_));
 sky130_fd_sc_hd__o2bb2ai_2 _18941_ (.A1_N(_08853_),
    .A2_N(_08855_),
    .B1(_08857_),
    .B2(_08546_),
    .Y(_08860_));
 sky130_fd_sc_hd__a311oi_2 _18942_ (.A1(_08842_),
    .A2(_08849_),
    .A3(_08850_),
    .B1(_08857_),
    .C1(_08546_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand3_1 _18943_ (.A(_08853_),
    .B(_08855_),
    .C(_08858_),
    .Y(_08862_));
 sky130_fd_sc_hd__a21o_1 _18944_ (.A1(_08853_),
    .A2(_08855_),
    .B1(_08859_),
    .X(_08863_));
 sky130_fd_sc_hd__o2111ai_4 _18945_ (.A1(_08545_),
    .A2(_08546_),
    .B1(_08549_),
    .C1(_08853_),
    .D1(_08855_),
    .Y(_08864_));
 sky130_fd_sc_hd__a2bb2oi_2 _18946_ (.A1_N(_08448_),
    .A2_N(_08453_),
    .B1(_08466_),
    .B2(_08452_),
    .Y(_08865_));
 sky130_fd_sc_hd__o22ai_4 _18947_ (.A1(_08448_),
    .A2(_08453_),
    .B1(_08467_),
    .B2(_08450_),
    .Y(_08866_));
 sky130_fd_sc_hd__and3_1 _18948_ (.A(_08863_),
    .B(_08865_),
    .C(_08864_),
    .X(_08868_));
 sky130_fd_sc_hd__nand3_4 _18949_ (.A(_08863_),
    .B(_08865_),
    .C(_08864_),
    .Y(_08869_));
 sky130_fd_sc_hd__nand3_4 _18950_ (.A(_08860_),
    .B(_08862_),
    .C(_08866_),
    .Y(_08870_));
 sky130_fd_sc_hd__o311a_1 _18951_ (.A1(_01923_),
    .A2(_02152_),
    .A3(_08245_),
    .B1(_08248_),
    .C1(_08557_),
    .X(_08871_));
 sky130_fd_sc_hd__o21ai_2 _18952_ (.A1(_08560_),
    .A2(_08555_),
    .B1(_08557_),
    .Y(_08872_));
 sky130_fd_sc_hd__o21a_1 _18953_ (.A1(_08560_),
    .A2(_08555_),
    .B1(_08557_),
    .X(_08873_));
 sky130_fd_sc_hd__o2bb2ai_2 _18954_ (.A1_N(_08869_),
    .A2_N(_08870_),
    .B1(_08871_),
    .B2(_08555_),
    .Y(_08874_));
 sky130_fd_sc_hd__nand2_1 _18955_ (.A(_08869_),
    .B(_08872_),
    .Y(_08875_));
 sky130_fd_sc_hd__nand3_2 _18956_ (.A(_08869_),
    .B(_08870_),
    .C(_08872_),
    .Y(_08876_));
 sky130_fd_sc_hd__a21o_1 _18957_ (.A1(_08869_),
    .A2(_08870_),
    .B1(_08873_),
    .X(_08877_));
 sky130_fd_sc_hd__o2111ai_2 _18958_ (.A1(_08560_),
    .A2(_08555_),
    .B1(_08557_),
    .C1(_08869_),
    .D1(_08870_),
    .Y(_08879_));
 sky130_fd_sc_hd__o2bb2ai_4 _18959_ (.A1_N(_08542_),
    .A2_N(_08568_),
    .B1(_08569_),
    .B2(_08563_),
    .Y(_08880_));
 sky130_fd_sc_hd__a2bb2oi_1 _18960_ (.A1_N(_08563_),
    .A2_N(_08569_),
    .B1(_08568_),
    .B2(_08542_),
    .Y(_08881_));
 sky130_fd_sc_hd__and3_2 _18961_ (.A(_08877_),
    .B(_08879_),
    .C(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__nand3_2 _18962_ (.A(_08877_),
    .B(_08879_),
    .C(_08881_),
    .Y(_08883_));
 sky130_fd_sc_hd__nand3_4 _18963_ (.A(_08874_),
    .B(_08880_),
    .C(_08876_),
    .Y(_08884_));
 sky130_fd_sc_hd__nand2_1 _18964_ (.A(_08883_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__nand3_2 _18965_ (.A(_08840_),
    .B(_08883_),
    .C(_08884_),
    .Y(_08886_));
 sky130_fd_sc_hd__o211ai_4 _18966_ (.A1(_08837_),
    .A2(_08835_),
    .B1(_08836_),
    .C1(_08885_),
    .Y(_08887_));
 sky130_fd_sc_hd__a22o_2 _18967_ (.A1(_08836_),
    .A2(_08839_),
    .B1(_08883_),
    .B2(_08884_),
    .X(_08888_));
 sky130_fd_sc_hd__o2111ai_4 _18968_ (.A1(_08837_),
    .A2(_08835_),
    .B1(_08836_),
    .C1(_08883_),
    .D1(_08884_),
    .Y(_08890_));
 sky130_fd_sc_hd__a22oi_4 _18969_ (.A1(_08481_),
    .A2(_08808_),
    .B1(_08888_),
    .B2(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__o211ai_4 _18970_ (.A1(_08480_),
    .A2(_08807_),
    .B1(_08886_),
    .C1(_08887_),
    .Y(_08892_));
 sky130_fd_sc_hd__a22oi_4 _18971_ (.A1(_08482_),
    .A2(_08809_),
    .B1(_08886_),
    .B2(_08887_),
    .Y(_08893_));
 sky130_fd_sc_hd__nand3_4 _18972_ (.A(_08888_),
    .B(_08890_),
    .C(_08810_),
    .Y(_08894_));
 sky130_fd_sc_hd__and3_1 _18973_ (.A(_08536_),
    .B(_08538_),
    .C(_08577_),
    .X(_08895_));
 sky130_fd_sc_hd__a31o_1 _18974_ (.A1(_08536_),
    .A2(_08538_),
    .A3(_08577_),
    .B1(_08578_),
    .X(_08896_));
 sky130_fd_sc_hd__a21boi_1 _18975_ (.A1(_08892_),
    .A2(_08894_),
    .B1_N(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__o2bb2ai_2 _18976_ (.A1_N(_08892_),
    .A2_N(_08894_),
    .B1(_08895_),
    .B2(_08578_),
    .Y(_08898_));
 sky130_fd_sc_hd__o311a_1 _18977_ (.A1(_08535_),
    .A2(_08537_),
    .A3(_08576_),
    .B1(_08579_),
    .C1(_08892_),
    .X(_08899_));
 sky130_fd_sc_hd__o211a_1 _18978_ (.A1(_08576_),
    .A2(_08582_),
    .B1(_08892_),
    .C1(_08894_),
    .X(_08901_));
 sky130_fd_sc_hd__o211ai_4 _18979_ (.A1(_08576_),
    .A2(_08582_),
    .B1(_08892_),
    .C1(_08894_),
    .Y(_08902_));
 sky130_fd_sc_hd__a21oi_1 _18980_ (.A1(_08892_),
    .A2(_08894_),
    .B1(_08896_),
    .Y(_08903_));
 sky130_fd_sc_hd__o22ai_4 _18981_ (.A1(_08576_),
    .A2(_08582_),
    .B1(_08891_),
    .B2(_08893_),
    .Y(_08904_));
 sky130_fd_sc_hd__and3_1 _18982_ (.A(_08892_),
    .B(_08894_),
    .C(_08896_),
    .X(_08905_));
 sky130_fd_sc_hd__o2111ai_4 _18983_ (.A1(_08578_),
    .A2(_08540_),
    .B1(_08577_),
    .C1(_08892_),
    .D1(_08894_),
    .Y(_08906_));
 sky130_fd_sc_hd__o22a_1 _18984_ (.A1(_08803_),
    .A2(_08805_),
    .B1(_08897_),
    .B2(_08901_),
    .X(_08907_));
 sky130_fd_sc_hd__o2bb2ai_1 _18985_ (.A1_N(_08804_),
    .A2_N(_08806_),
    .B1(_08897_),
    .B2(_08901_),
    .Y(_08908_));
 sky130_fd_sc_hd__nand4_2 _18986_ (.A(_08804_),
    .B(_08806_),
    .C(_08898_),
    .D(_08902_),
    .Y(_08909_));
 sky130_fd_sc_hd__nand4_2 _18987_ (.A(_08804_),
    .B(_08806_),
    .C(_08904_),
    .D(_08906_),
    .Y(_08910_));
 sky130_fd_sc_hd__o2bb2ai_2 _18988_ (.A1_N(_08804_),
    .A2_N(_08806_),
    .B1(_08903_),
    .B2(_08905_),
    .Y(_08912_));
 sky130_fd_sc_hd__nand3_1 _18989_ (.A(_08500_),
    .B(_08634_),
    .C(_08909_),
    .Y(_08913_));
 sky130_fd_sc_hd__a22oi_1 _18990_ (.A1(_08499_),
    .A2(_08635_),
    .B1(_08910_),
    .B2(_08912_),
    .Y(_08914_));
 sky130_fd_sc_hd__nand4_2 _18991_ (.A(_08500_),
    .B(_08634_),
    .C(_08908_),
    .D(_08909_),
    .Y(_08915_));
 sky130_fd_sc_hd__a22oi_1 _18992_ (.A1(_08500_),
    .A2(_08634_),
    .B1(_08908_),
    .B2(_08909_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand4_4 _18993_ (.A(_08499_),
    .B(_08635_),
    .C(_08910_),
    .D(_08912_),
    .Y(_08917_));
 sky130_fd_sc_hd__and3_1 _18994_ (.A(_08278_),
    .B(_08280_),
    .C(_08587_),
    .X(_08918_));
 sky130_fd_sc_hd__a31o_1 _18995_ (.A1(_08275_),
    .A2(_08501_),
    .A3(_08589_),
    .B1(_08586_),
    .X(_08919_));
 sky130_fd_sc_hd__o2111ai_1 _18996_ (.A1(_08588_),
    .A2(_08502_),
    .B1(_08587_),
    .C1(_08915_),
    .D1(_08917_),
    .Y(_08920_));
 sky130_fd_sc_hd__o22ai_1 _18997_ (.A1(_08586_),
    .A2(_08593_),
    .B1(_08914_),
    .B2(_08916_),
    .Y(_08921_));
 sky130_fd_sc_hd__o2bb2ai_2 _18998_ (.A1_N(_08915_),
    .A2_N(_08917_),
    .B1(_08918_),
    .B2(_08588_),
    .Y(_08923_));
 sky130_fd_sc_hd__o211ai_2 _18999_ (.A1(_08586_),
    .A2(_08593_),
    .B1(_08915_),
    .C1(_08917_),
    .Y(_08924_));
 sky130_fd_sc_hd__o2bb2ai_2 _19000_ (.A1_N(_08611_),
    .A2_N(_08607_),
    .B1(_08601_),
    .B2(_08608_),
    .Y(_08925_));
 sky130_fd_sc_hd__a2bb2oi_1 _19001_ (.A1_N(_08601_),
    .A2_N(_08608_),
    .B1(_08611_),
    .B2(_08607_),
    .Y(_08926_));
 sky130_fd_sc_hd__nand3_2 _19002_ (.A(_08920_),
    .B(_08921_),
    .C(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__nand3_4 _19003_ (.A(_08925_),
    .B(_08924_),
    .C(_08923_),
    .Y(_08928_));
 sky130_fd_sc_hd__o21ai_2 _19004_ (.A1(_08527_),
    .A2(_08529_),
    .B1(_08534_),
    .Y(_08929_));
 sky130_fd_sc_hd__a21oi_4 _19005_ (.A1(_08927_),
    .A2(_08928_),
    .B1(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__and3_1 _19006_ (.A(_08927_),
    .B(_08928_),
    .C(_08929_),
    .X(_08931_));
 sky130_fd_sc_hd__nand3_2 _19007_ (.A(_08927_),
    .B(_08928_),
    .C(_08929_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand2_1 _19008_ (.A(_08618_),
    .B(_08619_),
    .Y(_08934_));
 sky130_fd_sc_hd__o211ai_4 _19009_ (.A1(_08930_),
    .A2(_08931_),
    .B1(_08618_),
    .C1(_08623_),
    .Y(_08935_));
 sky130_fd_sc_hd__nand3_1 _19010_ (.A(_08617_),
    .B(_08932_),
    .C(_08934_),
    .Y(_08936_));
 sky130_fd_sc_hd__nor2_1 _19011_ (.A(_08930_),
    .B(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__o21ai_1 _19012_ (.A1(_08930_),
    .A2(_08936_),
    .B1(_08935_),
    .Y(_08938_));
 sky130_fd_sc_hd__xnor2_1 _19013_ (.A(_08633_),
    .B(_08938_),
    .Y(net97));
 sky130_fd_sc_hd__a31o_2 _19014_ (.A1(_08923_),
    .A2(_08924_),
    .A3(_08925_),
    .B1(_08931_),
    .X(_08939_));
 sky130_fd_sc_hd__a21oi_1 _19015_ (.A1(_08521_),
    .A2(_08832_),
    .B1(_08835_),
    .Y(_08940_));
 sky130_fd_sc_hd__a31oi_4 _19016_ (.A1(_08806_),
    .A2(_08898_),
    .A3(_08902_),
    .B1(_08803_),
    .Y(_08941_));
 sky130_fd_sc_hd__a31oi_4 _19017_ (.A1(_08804_),
    .A2(_08904_),
    .A3(_08906_),
    .B1(_08805_),
    .Y(_08942_));
 sky130_fd_sc_hd__nand3_4 _19018_ (.A(_08719_),
    .B(_08795_),
    .C(_08797_),
    .Y(_08944_));
 sky130_fd_sc_hd__o41ai_4 _19019_ (.A1(_08358_),
    .A2(_08640_),
    .A3(_08714_),
    .A4(_08716_),
    .B1(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__nand2_1 _19020_ (.A(_08667_),
    .B(_08712_),
    .Y(_08946_));
 sky130_fd_sc_hd__o21ai_1 _19021_ (.A1(_08707_),
    .A2(_08946_),
    .B1(_08669_),
    .Y(_08947_));
 sky130_fd_sc_hd__a31oi_2 _19022_ (.A1(_08667_),
    .A2(_08708_),
    .A3(_08712_),
    .B1(_08668_),
    .Y(_08948_));
 sky130_fd_sc_hd__nand3_1 _19023_ (.A(_08007_),
    .B(_08658_),
    .C(_08660_),
    .Y(_08949_));
 sky130_fd_sc_hd__a31o_2 _19024_ (.A1(_08661_),
    .A2(_08662_),
    .A3(_08008_),
    .B1(_08006_),
    .X(_08950_));
 sky130_fd_sc_hd__a31oi_1 _19025_ (.A1(_08661_),
    .A2(_08662_),
    .A3(_08008_),
    .B1(_08006_),
    .Y(_08951_));
 sky130_fd_sc_hd__o31a_2 _19026_ (.A1(_01890_),
    .A2(_02251_),
    .A3(_08332_),
    .B1(_08335_),
    .X(_08952_));
 sky130_fd_sc_hd__nand2_2 _19027_ (.A(_08335_),
    .B(_08646_),
    .Y(_08953_));
 sky130_fd_sc_hd__o21ai_4 _19028_ (.A1(_08651_),
    .A2(_08654_),
    .B1(_08952_),
    .Y(_08955_));
 sky130_fd_sc_hd__o211ai_4 _19029_ (.A1(_08647_),
    .A2(_08653_),
    .B1(_08953_),
    .C1(_08652_),
    .Y(_08956_));
 sky130_fd_sc_hd__o22ai_4 _19030_ (.A1(_08334_),
    .A2(_08645_),
    .B1(_08651_),
    .B2(_08654_),
    .Y(_08957_));
 sky130_fd_sc_hd__o211ai_4 _19031_ (.A1(_08647_),
    .A2(_08653_),
    .B1(_08952_),
    .C1(_08652_),
    .Y(_08958_));
 sky130_fd_sc_hd__nand2_4 _19032_ (.A(_08957_),
    .B(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__nand3_1 _19033_ (.A(_08009_),
    .B(_08955_),
    .C(_08956_),
    .Y(_08960_));
 sky130_fd_sc_hd__nand4_2 _19034_ (.A(_08004_),
    .B(_08007_),
    .C(_08957_),
    .D(_08958_),
    .Y(_08961_));
 sky130_fd_sc_hd__and3_2 _19035_ (.A(_08009_),
    .B(_08957_),
    .C(_08958_),
    .X(_08962_));
 sky130_fd_sc_hd__nand3_4 _19036_ (.A(_08009_),
    .B(_08957_),
    .C(_08958_),
    .Y(_08963_));
 sky130_fd_sc_hd__nand3_1 _19037_ (.A(_08955_),
    .B(_08956_),
    .C(_08008_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand2_2 _19038_ (.A(_08960_),
    .B(_08961_),
    .Y(_08966_));
 sky130_fd_sc_hd__and3_1 _19039_ (.A(_08951_),
    .B(_08960_),
    .C(_08961_),
    .X(_08967_));
 sky130_fd_sc_hd__nand3_2 _19040_ (.A(_08951_),
    .B(_08960_),
    .C(_08961_),
    .Y(_08968_));
 sky130_fd_sc_hd__nand4_4 _19041_ (.A(_08004_),
    .B(_08949_),
    .C(_08963_),
    .D(_08964_),
    .Y(_08969_));
 sky130_fd_sc_hd__nor2_1 _19042_ (.A(_08683_),
    .B(_08684_),
    .Y(_08970_));
 sky130_fd_sc_hd__o21a_1 _19043_ (.A1(_08683_),
    .A2(_08684_),
    .B1(_08687_),
    .X(_08971_));
 sky130_fd_sc_hd__nand2_2 _19044_ (.A(net35),
    .B(net22),
    .Y(_08972_));
 sky130_fd_sc_hd__nand2_1 _19045_ (.A(net64),
    .B(net25),
    .Y(_08973_));
 sky130_fd_sc_hd__a22oi_4 _19046_ (.A1(net34),
    .A2(net24),
    .B1(net25),
    .B2(net64),
    .Y(_08974_));
 sky130_fd_sc_hd__a22o_1 _19047_ (.A1(net34),
    .A2(net24),
    .B1(net25),
    .B2(net64),
    .X(_08975_));
 sky130_fd_sc_hd__nand2_1 _19048_ (.A(net34),
    .B(net25),
    .Y(_08977_));
 sky130_fd_sc_hd__nand2_2 _19049_ (.A(net64),
    .B(net34),
    .Y(_08978_));
 sky130_fd_sc_hd__nand3_4 _19050_ (.A(net64),
    .B(net34),
    .C(net25),
    .Y(_08979_));
 sky130_fd_sc_hd__and4_1 _19051_ (.A(net64),
    .B(net34),
    .C(net24),
    .D(net25),
    .X(_08980_));
 sky130_fd_sc_hd__o221ai_4 _19052_ (.A1(_01934_),
    .A2(_02196_),
    .B1(_02218_),
    .B2(_08979_),
    .C1(_08975_),
    .Y(_08981_));
 sky130_fd_sc_hd__o21bai_1 _19053_ (.A1(_08974_),
    .A2(_08980_),
    .B1_N(_08972_),
    .Y(_08982_));
 sky130_fd_sc_hd__o2111ai_4 _19054_ (.A1(_02218_),
    .A2(_08979_),
    .B1(net35),
    .C1(net22),
    .D1(_08975_),
    .Y(_08983_));
 sky130_fd_sc_hd__o21ai_1 _19055_ (.A1(_08974_),
    .A2(_08980_),
    .B1(_08972_),
    .Y(_08984_));
 sky130_fd_sc_hd__o211ai_4 _19056_ (.A1(_08686_),
    .A2(_08970_),
    .B1(_08983_),
    .C1(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__nand3_4 _19057_ (.A(_08971_),
    .B(_08981_),
    .C(_08982_),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_1 _19058_ (.A(net38),
    .B(net19),
    .Y(_08988_));
 sky130_fd_sc_hd__and4_1 _19059_ (.A(net36),
    .B(net37),
    .C(net20),
    .D(net21),
    .X(_08989_));
 sky130_fd_sc_hd__nand4_2 _19060_ (.A(net36),
    .B(net37),
    .C(net20),
    .D(net21),
    .Y(_08990_));
 sky130_fd_sc_hd__a22oi_4 _19061_ (.A1(net37),
    .A2(net20),
    .B1(net21),
    .B2(net36),
    .Y(_08991_));
 sky130_fd_sc_hd__a22o_1 _19062_ (.A1(net37),
    .A2(net20),
    .B1(net21),
    .B2(net36),
    .X(_08992_));
 sky130_fd_sc_hd__and3_1 _19063_ (.A(_08988_),
    .B(_08990_),
    .C(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__o211a_1 _19064_ (.A1(_08989_),
    .A2(_08991_),
    .B1(net38),
    .C1(net19),
    .X(_08994_));
 sky130_fd_sc_hd__o21a_1 _19065_ (.A1(_08989_),
    .A2(_08991_),
    .B1(_08988_),
    .X(_08995_));
 sky130_fd_sc_hd__and4_1 _19066_ (.A(_08992_),
    .B(net19),
    .C(net38),
    .D(_08990_),
    .X(_08996_));
 sky130_fd_sc_hd__o2bb2ai_4 _19067_ (.A1_N(_08985_),
    .A2_N(_08986_),
    .B1(_08993_),
    .B2(_08994_),
    .Y(_08997_));
 sky130_fd_sc_hd__o211ai_4 _19068_ (.A1(_08995_),
    .A2(_08996_),
    .B1(_08985_),
    .C1(_08986_),
    .Y(_08999_));
 sky130_fd_sc_hd__o2bb2ai_1 _19069_ (.A1_N(_08985_),
    .A2_N(_08986_),
    .B1(_08995_),
    .B2(_08996_),
    .Y(_09000_));
 sky130_fd_sc_hd__o21ai_1 _19070_ (.A1(_08993_),
    .A2(_08994_),
    .B1(_08986_),
    .Y(_09001_));
 sky130_fd_sc_hd__o211ai_1 _19071_ (.A1(_08993_),
    .A2(_08994_),
    .B1(_08985_),
    .C1(_08986_),
    .Y(_09002_));
 sky130_fd_sc_hd__o21ai_1 _19072_ (.A1(_08657_),
    .A2(_08651_),
    .B1(_08655_),
    .Y(_09003_));
 sky130_fd_sc_hd__a21oi_4 _19073_ (.A1(_08652_),
    .A2(_08656_),
    .B1(_08654_),
    .Y(_09004_));
 sky130_fd_sc_hd__nand3_2 _19074_ (.A(_08997_),
    .B(_08999_),
    .C(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__a21oi_4 _19075_ (.A1(_08997_),
    .A2(_08999_),
    .B1(_09004_),
    .Y(_09006_));
 sky130_fd_sc_hd__nand3_2 _19076_ (.A(_09000_),
    .B(_09002_),
    .C(_09003_),
    .Y(_09007_));
 sky130_fd_sc_hd__nand2_1 _19077_ (.A(_08694_),
    .B(_08699_),
    .Y(_09008_));
 sky130_fd_sc_hd__a21o_2 _19078_ (.A1(_09005_),
    .A2(_09007_),
    .B1(_09008_),
    .X(_09010_));
 sky130_fd_sc_hd__a32oi_4 _19079_ (.A1(_08997_),
    .A2(_08999_),
    .A3(_09004_),
    .B1(_08699_),
    .B2(_08694_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_1 _19080_ (.A(_09005_),
    .B(_09008_),
    .Y(_09012_));
 sky130_fd_sc_hd__nand3_2 _19081_ (.A(_09005_),
    .B(_09007_),
    .C(_09008_),
    .Y(_09013_));
 sky130_fd_sc_hd__a22o_1 _19082_ (.A1(_08694_),
    .A2(_08699_),
    .B1(_09005_),
    .B2(_09007_),
    .X(_09014_));
 sky130_fd_sc_hd__nand4_1 _19083_ (.A(_08694_),
    .B(_08699_),
    .C(_09005_),
    .D(_09007_),
    .Y(_09015_));
 sky130_fd_sc_hd__o2111a_1 _19084_ (.A1(_09012_),
    .A2(_09006_),
    .B1(_08969_),
    .C1(_08968_),
    .D1(_09010_),
    .X(_09016_));
 sky130_fd_sc_hd__o2111ai_4 _19085_ (.A1(_09012_),
    .A2(_09006_),
    .B1(_08969_),
    .C1(_08968_),
    .D1(_09010_),
    .Y(_09017_));
 sky130_fd_sc_hd__a22oi_2 _19086_ (.A1(_08968_),
    .A2(_08969_),
    .B1(_09010_),
    .B2(_09013_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand3b_4 _19087_ (.A_N(_09018_),
    .B(_08947_),
    .C(_09017_),
    .Y(_09019_));
 sky130_fd_sc_hd__o21a_1 _19088_ (.A1(_09016_),
    .A2(_09018_),
    .B1(_08948_),
    .X(_09021_));
 sky130_fd_sc_hd__o21ai_2 _19089_ (.A1(_09016_),
    .A2(_09018_),
    .B1(_08948_),
    .Y(_09022_));
 sky130_fd_sc_hd__nand2_1 _19090_ (.A(_08704_),
    .B(_08705_),
    .Y(_09023_));
 sky130_fd_sc_hd__o21ai_1 _19091_ (.A1(_08706_),
    .A2(_08703_),
    .B1(_08702_),
    .Y(_09024_));
 sky130_fd_sc_hd__o31a_1 _19092_ (.A1(_08414_),
    .A2(_08750_),
    .A3(_08767_),
    .B1(_08766_),
    .X(_09025_));
 sky130_fd_sc_hd__o21ai_1 _19093_ (.A1(_08751_),
    .A2(_08767_),
    .B1(_08766_),
    .Y(_09026_));
 sky130_fd_sc_hd__a21o_1 _19094_ (.A1(_08673_),
    .A2(_08671_),
    .B1(_08674_),
    .X(_09027_));
 sky130_fd_sc_hd__a21oi_1 _19095_ (.A1(_08673_),
    .A2(_08671_),
    .B1(_08674_),
    .Y(_09028_));
 sky130_fd_sc_hd__nand2_1 _19096_ (.A(net41),
    .B(net16),
    .Y(_09029_));
 sky130_fd_sc_hd__a22oi_4 _19097_ (.A1(net40),
    .A2(net17),
    .B1(net18),
    .B2(net39),
    .Y(_09030_));
 sky130_fd_sc_hd__a22o_1 _19098_ (.A1(net40),
    .A2(net17),
    .B1(net18),
    .B2(net39),
    .X(_09032_));
 sky130_fd_sc_hd__and4_1 _19099_ (.A(net39),
    .B(net40),
    .C(net17),
    .D(net18),
    .X(_09033_));
 sky130_fd_sc_hd__nand4_4 _19100_ (.A(net39),
    .B(net40),
    .C(net17),
    .D(net18),
    .Y(_09034_));
 sky130_fd_sc_hd__o211ai_2 _19101_ (.A1(_02010_),
    .A2(_02098_),
    .B1(_09032_),
    .C1(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__o21bai_1 _19102_ (.A1(_09030_),
    .A2(_09033_),
    .B1_N(_09029_),
    .Y(_09036_));
 sky130_fd_sc_hd__o21ai_2 _19103_ (.A1(_09030_),
    .A2(_09033_),
    .B1(_09029_),
    .Y(_09037_));
 sky130_fd_sc_hd__and4_1 _19104_ (.A(_09032_),
    .B(_09034_),
    .C(net41),
    .D(net16),
    .X(_09038_));
 sky130_fd_sc_hd__nand4_2 _19105_ (.A(_09032_),
    .B(_09034_),
    .C(net41),
    .D(net16),
    .Y(_09039_));
 sky130_fd_sc_hd__nand3_4 _19106_ (.A(_09028_),
    .B(_09035_),
    .C(_09036_),
    .Y(_09040_));
 sky130_fd_sc_hd__nand2_1 _19107_ (.A(_09027_),
    .B(_09037_),
    .Y(_09041_));
 sky130_fd_sc_hd__nand3_4 _19108_ (.A(_09027_),
    .B(_09037_),
    .C(_09039_),
    .Y(_09043_));
 sky130_fd_sc_hd__o21a_1 _19109_ (.A1(_02010_),
    .A2(_02076_),
    .B1(_08760_),
    .X(_09044_));
 sky130_fd_sc_hd__a31o_1 _19110_ (.A1(_08758_),
    .A2(net15),
    .A3(net41),
    .B1(_08759_),
    .X(_09045_));
 sky130_fd_sc_hd__o2bb2ai_2 _19111_ (.A1_N(_09040_),
    .A2_N(_09043_),
    .B1(_09044_),
    .B2(_08756_),
    .Y(_09046_));
 sky130_fd_sc_hd__nand2_1 _19112_ (.A(_09040_),
    .B(_09045_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand3_4 _19113_ (.A(_09040_),
    .B(_09043_),
    .C(_09045_),
    .Y(_09048_));
 sky130_fd_sc_hd__nand2_1 _19114_ (.A(_09046_),
    .B(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__a21oi_2 _19115_ (.A1(_09046_),
    .A2(_09048_),
    .B1(_09026_),
    .Y(_09050_));
 sky130_fd_sc_hd__a21o_1 _19116_ (.A1(_09046_),
    .A2(_09048_),
    .B1(_09026_),
    .X(_09051_));
 sky130_fd_sc_hd__o211a_1 _19117_ (.A1(_08765_),
    .A2(_08770_),
    .B1(_09046_),
    .C1(_09048_),
    .X(_09052_));
 sky130_fd_sc_hd__o211ai_1 _19118_ (.A1(_08765_),
    .A2(_08770_),
    .B1(_09046_),
    .C1(_09048_),
    .Y(_09054_));
 sky130_fd_sc_hd__o21ai_1 _19119_ (.A1(_08722_),
    .A2(_08726_),
    .B1(_08725_),
    .Y(_09055_));
 sky130_fd_sc_hd__nand2_2 _19120_ (.A(net13),
    .B(net45),
    .Y(_09056_));
 sky130_fd_sc_hd__nand2_2 _19121_ (.A(net42),
    .B(net15),
    .Y(_09057_));
 sky130_fd_sc_hd__and4_2 _19122_ (.A(net42),
    .B(net43),
    .C(net14),
    .D(net15),
    .X(_09058_));
 sky130_fd_sc_hd__nand4_1 _19123_ (.A(net42),
    .B(net43),
    .C(net14),
    .D(net15),
    .Y(_09059_));
 sky130_fd_sc_hd__a22oi_4 _19124_ (.A1(net43),
    .A2(net14),
    .B1(net15),
    .B2(net42),
    .Y(_09060_));
 sky130_fd_sc_hd__a22o_1 _19125_ (.A1(net43),
    .A2(net14),
    .B1(net15),
    .B2(net42),
    .X(_09061_));
 sky130_fd_sc_hd__a2bb2oi_1 _19126_ (.A1_N(_02043_),
    .A2_N(_02054_),
    .B1(_09059_),
    .B2(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__o21ai_2 _19127_ (.A1(_09058_),
    .A2(_09060_),
    .B1(_09056_),
    .Y(_09063_));
 sky130_fd_sc_hd__nor3_4 _19128_ (.A(_09060_),
    .B(_09056_),
    .C(_09058_),
    .Y(_09065_));
 sky130_fd_sc_hd__nand4_1 _19129_ (.A(_09061_),
    .B(net45),
    .C(net13),
    .D(_09059_),
    .Y(_09066_));
 sky130_fd_sc_hd__a21oi_1 _19130_ (.A1(_09063_),
    .A2(_09066_),
    .B1(_09055_),
    .Y(_09067_));
 sky130_fd_sc_hd__o21bai_2 _19131_ (.A1(_09062_),
    .A2(_09065_),
    .B1_N(_09055_),
    .Y(_09068_));
 sky130_fd_sc_hd__nand2_1 _19132_ (.A(_09063_),
    .B(_09055_),
    .Y(_09069_));
 sky130_fd_sc_hd__nand3_1 _19133_ (.A(_09063_),
    .B(_09066_),
    .C(_09055_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand2_1 _19134_ (.A(net9),
    .B(net48),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_2 _19135_ (.A(net11),
    .B(net47),
    .Y(_09072_));
 sky130_fd_sc_hd__nand2_1 _19136_ (.A(net11),
    .B(net46),
    .Y(_09073_));
 sky130_fd_sc_hd__and4_1 _19137_ (.A(net10),
    .B(net11),
    .C(net46),
    .D(net47),
    .X(_09074_));
 sky130_fd_sc_hd__nand4_1 _19138_ (.A(net10),
    .B(net11),
    .C(net46),
    .D(net47),
    .Y(_09076_));
 sky130_fd_sc_hd__a22o_1 _19139_ (.A1(net11),
    .A2(net46),
    .B1(net47),
    .B2(net10),
    .X(_09077_));
 sky130_fd_sc_hd__o221a_1 _19140_ (.A1(_01999_),
    .A2(_02109_),
    .B1(_08737_),
    .B2(_09072_),
    .C1(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__a21oi_1 _19141_ (.A1(_09076_),
    .A2(_09077_),
    .B1(_09071_),
    .Y(_09079_));
 sky130_fd_sc_hd__nor2_2 _19142_ (.A(_09078_),
    .B(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__o2bb2a_1 _19143_ (.A1_N(_09068_),
    .A2_N(_09070_),
    .B1(_09078_),
    .B2(_09079_),
    .X(_09081_));
 sky130_fd_sc_hd__a21o_1 _19144_ (.A1(_09068_),
    .A2(_09070_),
    .B1(_09080_),
    .X(_09082_));
 sky130_fd_sc_hd__and3_1 _19145_ (.A(_09068_),
    .B(_09080_),
    .C(_09070_),
    .X(_09083_));
 sky130_fd_sc_hd__o211ai_2 _19146_ (.A1(_09065_),
    .A2(_09069_),
    .B1(_09080_),
    .C1(_09068_),
    .Y(_09084_));
 sky130_fd_sc_hd__nand2_1 _19147_ (.A(_09082_),
    .B(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__o21bai_1 _19148_ (.A1(_09050_),
    .A2(_09052_),
    .B1_N(_09085_),
    .Y(_09087_));
 sky130_fd_sc_hd__o2bb2ai_2 _19149_ (.A1_N(_09049_),
    .A2_N(_09025_),
    .B1(_09083_),
    .B2(_09081_),
    .Y(_09088_));
 sky130_fd_sc_hd__o21ai_2 _19150_ (.A1(_09050_),
    .A2(_09052_),
    .B1(_09085_),
    .Y(_09089_));
 sky130_fd_sc_hd__nand4_2 _19151_ (.A(_09051_),
    .B(_09054_),
    .C(_09082_),
    .D(_09084_),
    .Y(_09090_));
 sky130_fd_sc_hd__nand2_1 _19152_ (.A(_09089_),
    .B(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__nand3_4 _19153_ (.A(_09089_),
    .B(_09090_),
    .C(_09024_),
    .Y(_09092_));
 sky130_fd_sc_hd__o221ai_4 _19154_ (.A1(_08703_),
    .A2(_08709_),
    .B1(_09052_),
    .B2(_09088_),
    .C1(_09087_),
    .Y(_09093_));
 sky130_fd_sc_hd__o31a_2 _19155_ (.A1(_08744_),
    .A2(_08745_),
    .A3(_08773_),
    .B1(_08776_),
    .X(_09094_));
 sky130_fd_sc_hd__o31a_2 _19156_ (.A1(_08747_),
    .A2(_08748_),
    .A3(_08775_),
    .B1(_08774_),
    .X(_09095_));
 sky130_fd_sc_hd__a21oi_1 _19157_ (.A1(_09092_),
    .A2(_09093_),
    .B1(_09094_),
    .Y(_09096_));
 sky130_fd_sc_hd__a21o_1 _19158_ (.A1(_09092_),
    .A2(_09093_),
    .B1(_09094_),
    .X(_09098_));
 sky130_fd_sc_hd__and3_1 _19159_ (.A(_09092_),
    .B(_09093_),
    .C(_09094_),
    .X(_09099_));
 sky130_fd_sc_hd__nand3_1 _19160_ (.A(_09092_),
    .B(_09093_),
    .C(_09094_),
    .Y(_09100_));
 sky130_fd_sc_hd__a21oi_1 _19161_ (.A1(_09092_),
    .A2(_09093_),
    .B1(_09095_),
    .Y(_09101_));
 sky130_fd_sc_hd__a21o_1 _19162_ (.A1(_09092_),
    .A2(_09093_),
    .B1(_09095_),
    .X(_09102_));
 sky130_fd_sc_hd__and3_1 _19163_ (.A(_09092_),
    .B(_09093_),
    .C(_09095_),
    .X(_09103_));
 sky130_fd_sc_hd__nand3_2 _19164_ (.A(_09092_),
    .B(_09093_),
    .C(_09095_),
    .Y(_09104_));
 sky130_fd_sc_hd__nand4_2 _19165_ (.A(_09019_),
    .B(_09022_),
    .C(_09102_),
    .D(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__o2bb2ai_1 _19166_ (.A1_N(_09019_),
    .A2_N(_09022_),
    .B1(_09101_),
    .B2(_09103_),
    .Y(_09106_));
 sky130_fd_sc_hd__o2bb2ai_2 _19167_ (.A1_N(_09019_),
    .A2_N(_09022_),
    .B1(_09096_),
    .B2(_09099_),
    .Y(_09107_));
 sky130_fd_sc_hd__nand4_2 _19168_ (.A(_09019_),
    .B(_09022_),
    .C(_09098_),
    .D(_09100_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand3_4 _19169_ (.A(_08945_),
    .B(_09107_),
    .C(_09109_),
    .Y(_09110_));
 sky130_fd_sc_hd__a21oi_2 _19170_ (.A1(_09107_),
    .A2(_09109_),
    .B1(_08945_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand4_4 _19171_ (.A(_08718_),
    .B(_08944_),
    .C(_09105_),
    .D(_09106_),
    .Y(_09112_));
 sky130_fd_sc_hd__o21ai_1 _19172_ (.A1(_08829_),
    .A2(_08825_),
    .B1(_08824_),
    .Y(_09113_));
 sky130_fd_sc_hd__o22ai_1 _19173_ (.A1(_08509_),
    .A2(_08815_),
    .B1(_08814_),
    .B2(_08817_),
    .Y(_09114_));
 sky130_fd_sc_hd__nand2_1 _19174_ (.A(net3),
    .B(net54),
    .Y(_09115_));
 sky130_fd_sc_hd__a22oi_4 _19175_ (.A1(net5),
    .A2(net52),
    .B1(net53),
    .B2(net4),
    .Y(_09116_));
 sky130_fd_sc_hd__a22o_1 _19176_ (.A1(net5),
    .A2(net52),
    .B1(net53),
    .B2(net4),
    .X(_09117_));
 sky130_fd_sc_hd__and4_1 _19177_ (.A(net4),
    .B(net5),
    .C(net52),
    .D(net53),
    .X(_09118_));
 sky130_fd_sc_hd__nand4_2 _19178_ (.A(net4),
    .B(net5),
    .C(net52),
    .D(net53),
    .Y(_09120_));
 sky130_fd_sc_hd__o211ai_1 _19179_ (.A1(_01923_),
    .A2(_02207_),
    .B1(_09117_),
    .C1(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__o21bai_1 _19180_ (.A1(_09116_),
    .A2(_09118_),
    .B1_N(_09115_),
    .Y(_09122_));
 sky130_fd_sc_hd__o21ai_1 _19181_ (.A1(_09116_),
    .A2(_09118_),
    .B1(_09115_),
    .Y(_09123_));
 sky130_fd_sc_hd__nand4_1 _19182_ (.A(_09117_),
    .B(_09120_),
    .C(net3),
    .D(net54),
    .Y(_09124_));
 sky130_fd_sc_hd__nand3b_1 _19183_ (.A_N(_09114_),
    .B(_09121_),
    .C(_09122_),
    .Y(_09125_));
 sky130_fd_sc_hd__a22oi_1 _19184_ (.A1(_08816_),
    .A2(_08820_),
    .B1(_09121_),
    .B2(_09122_),
    .Y(_09126_));
 sky130_fd_sc_hd__nand3_1 _19185_ (.A(_09114_),
    .B(_09123_),
    .C(_09124_),
    .Y(_09127_));
 sky130_fd_sc_hd__nand2_1 _19186_ (.A(_01912_),
    .B(net57),
    .Y(_09128_));
 sky130_fd_sc_hd__and4_2 _19187_ (.A(_01912_),
    .B(net56),
    .C(net57),
    .D(net2),
    .X(_09129_));
 sky130_fd_sc_hd__o22a_1 _19188_ (.A1(net32),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01901_),
    .X(_09131_));
 sky130_fd_sc_hd__nor2_1 _19189_ (.A(_09129_),
    .B(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__o2bb2ai_1 _19190_ (.A1_N(_09125_),
    .A2_N(_09127_),
    .B1(_09129_),
    .B2(_09131_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand3_1 _19191_ (.A(_09125_),
    .B(_09127_),
    .C(_09132_),
    .Y(_09134_));
 sky130_fd_sc_hd__a21oi_2 _19192_ (.A1(_09133_),
    .A2(_09134_),
    .B1(_09113_),
    .Y(_09135_));
 sky130_fd_sc_hd__and3_1 _19193_ (.A(_09113_),
    .B(_09133_),
    .C(_09134_),
    .X(_09136_));
 sky130_fd_sc_hd__nor3_2 _19194_ (.A(_08827_),
    .B(_09135_),
    .C(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__o21a_1 _19195_ (.A1(_09135_),
    .A2(_09136_),
    .B1(_08827_),
    .X(_09138_));
 sky130_fd_sc_hd__nor2_2 _19196_ (.A(_09137_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__a21oi_2 _19197_ (.A1(_08458_),
    .A2(_08737_),
    .B1(_08736_),
    .Y(_09140_));
 sky130_fd_sc_hd__nor2_1 _19198_ (.A(_08738_),
    .B(_09140_),
    .Y(_09142_));
 sky130_fd_sc_hd__nor2_1 _19199_ (.A(_01966_),
    .B(_02152_),
    .Y(_09143_));
 sky130_fd_sc_hd__a22oi_4 _19200_ (.A1(net8),
    .A2(net49),
    .B1(net50),
    .B2(net7),
    .Y(_09144_));
 sky130_fd_sc_hd__a22o_1 _19201_ (.A1(net8),
    .A2(net49),
    .B1(net50),
    .B2(net7),
    .X(_09145_));
 sky130_fd_sc_hd__nand2_2 _19202_ (.A(net8),
    .B(net50),
    .Y(_09146_));
 sky130_fd_sc_hd__and4_1 _19203_ (.A(net7),
    .B(net8),
    .C(net49),
    .D(net50),
    .X(_09147_));
 sky130_fd_sc_hd__nand4_1 _19204_ (.A(net7),
    .B(net8),
    .C(net49),
    .D(net50),
    .Y(_09148_));
 sky130_fd_sc_hd__o211ai_2 _19205_ (.A1(_01966_),
    .A2(_02152_),
    .B1(_09145_),
    .C1(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__o21ai_1 _19206_ (.A1(_09144_),
    .A2(_09147_),
    .B1(_09143_),
    .Y(_09150_));
 sky130_fd_sc_hd__o22ai_2 _19207_ (.A1(_01966_),
    .A2(_02152_),
    .B1(_09144_),
    .B2(_09147_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand4_1 _19208_ (.A(_09145_),
    .B(_09148_),
    .C(net6),
    .D(net51),
    .Y(_09153_));
 sky130_fd_sc_hd__nand3_4 _19209_ (.A(_09142_),
    .B(_09149_),
    .C(_09150_),
    .Y(_09154_));
 sky130_fd_sc_hd__o211ai_4 _19210_ (.A1(_08738_),
    .A2(_09140_),
    .B1(_09151_),
    .C1(_09153_),
    .Y(_09155_));
 sky130_fd_sc_hd__inv_2 _19211_ (.A(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__o21a_1 _19212_ (.A1(_01956_),
    .A2(_02152_),
    .B1(_08848_),
    .X(_09157_));
 sky130_fd_sc_hd__a31o_2 _19213_ (.A1(_08846_),
    .A2(net51),
    .A3(net5),
    .B1(_08847_),
    .X(_09158_));
 sky130_fd_sc_hd__o2bb2ai_4 _19214_ (.A1_N(_09154_),
    .A2_N(_09155_),
    .B1(_09157_),
    .B2(_08844_),
    .Y(_09159_));
 sky130_fd_sc_hd__nand2_1 _19215_ (.A(_09154_),
    .B(_09158_),
    .Y(_09160_));
 sky130_fd_sc_hd__and3_1 _19216_ (.A(_09154_),
    .B(_09155_),
    .C(_09158_),
    .X(_09161_));
 sky130_fd_sc_hd__nand3_2 _19217_ (.A(_09154_),
    .B(_09155_),
    .C(_09158_),
    .Y(_09162_));
 sky130_fd_sc_hd__nand2_1 _19218_ (.A(_09159_),
    .B(_09162_),
    .Y(_09164_));
 sky130_fd_sc_hd__o22a_1 _19219_ (.A1(_08729_),
    .A2(_08733_),
    .B1(_08743_),
    .B2(_08731_),
    .X(_09165_));
 sky130_fd_sc_hd__o22ai_4 _19220_ (.A1(_08729_),
    .A2(_08733_),
    .B1(_08743_),
    .B2(_08731_),
    .Y(_09166_));
 sky130_fd_sc_hd__a21oi_4 _19221_ (.A1(_09159_),
    .A2(_09162_),
    .B1(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__a21o_1 _19222_ (.A1(_09159_),
    .A2(_09162_),
    .B1(_09166_),
    .X(_09168_));
 sky130_fd_sc_hd__o211a_2 _19223_ (.A1(_09160_),
    .A2(_09156_),
    .B1(_09159_),
    .C1(_09166_),
    .X(_09169_));
 sky130_fd_sc_hd__o211ai_4 _19224_ (.A1(_09160_),
    .A2(_09156_),
    .B1(_09159_),
    .C1(_09166_),
    .Y(_09170_));
 sky130_fd_sc_hd__a21oi_4 _19225_ (.A1(_08853_),
    .A2(_08858_),
    .B1(_08854_),
    .Y(_09171_));
 sky130_fd_sc_hd__a21oi_2 _19226_ (.A1(_09164_),
    .A2(_09165_),
    .B1(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__o21ai_2 _19227_ (.A1(_09164_),
    .A2(_09165_),
    .B1(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__o21ai_1 _19228_ (.A1(_09167_),
    .A2(_09169_),
    .B1(_09171_),
    .Y(_09175_));
 sky130_fd_sc_hd__o22ai_4 _19229_ (.A1(_08854_),
    .A2(_08861_),
    .B1(_09167_),
    .B2(_09169_),
    .Y(_09176_));
 sky130_fd_sc_hd__nand3_4 _19230_ (.A(_09168_),
    .B(_09170_),
    .C(_09171_),
    .Y(_09177_));
 sky130_fd_sc_hd__o21a_1 _19231_ (.A1(_08555_),
    .A2(_08871_),
    .B1(_08870_),
    .X(_09178_));
 sky130_fd_sc_hd__a31o_1 _19232_ (.A1(_08860_),
    .A2(_08862_),
    .A3(_08866_),
    .B1(_08872_),
    .X(_09179_));
 sky130_fd_sc_hd__a22oi_4 _19233_ (.A1(_08870_),
    .A2(_08875_),
    .B1(_09176_),
    .B2(_09177_),
    .Y(_09180_));
 sky130_fd_sc_hd__nand4_4 _19234_ (.A(_08869_),
    .B(_09173_),
    .C(_09175_),
    .D(_09179_),
    .Y(_09181_));
 sky130_fd_sc_hd__o211a_2 _19235_ (.A1(_08868_),
    .A2(_09178_),
    .B1(_09177_),
    .C1(_09176_),
    .X(_09182_));
 sky130_fd_sc_hd__o2111ai_4 _19236_ (.A1(_08873_),
    .A2(_08868_),
    .B1(_08870_),
    .C1(_09176_),
    .D1(_09177_),
    .Y(_09183_));
 sky130_fd_sc_hd__o31a_1 _19237_ (.A1(_09137_),
    .A2(_09138_),
    .A3(_09180_),
    .B1(_09183_),
    .X(_09184_));
 sky130_fd_sc_hd__nand3_1 _19238_ (.A(_09139_),
    .B(_09181_),
    .C(_09183_),
    .Y(_09186_));
 sky130_fd_sc_hd__o22ai_2 _19239_ (.A1(_09137_),
    .A2(_09138_),
    .B1(_09180_),
    .B2(_09182_),
    .Y(_09187_));
 sky130_fd_sc_hd__o21ai_2 _19240_ (.A1(_09180_),
    .A2(_09182_),
    .B1(_09139_),
    .Y(_09188_));
 sky130_fd_sc_hd__o211ai_2 _19241_ (.A1(_09137_),
    .A2(_09138_),
    .B1(_09181_),
    .C1(_09183_),
    .Y(_09189_));
 sky130_fd_sc_hd__o2bb2ai_2 _19242_ (.A1_N(_08788_),
    .A2_N(_08786_),
    .B1(_08783_),
    .B2(_08777_),
    .Y(_09190_));
 sky130_fd_sc_hd__a21oi_2 _19243_ (.A1(_08786_),
    .A2(_08788_),
    .B1(_08784_),
    .Y(_09191_));
 sky130_fd_sc_hd__nand3_4 _19244_ (.A(_09186_),
    .B(_09187_),
    .C(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__inv_2 _19245_ (.A(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__and3_2 _19246_ (.A(_09188_),
    .B(_09189_),
    .C(_09190_),
    .X(_09194_));
 sky130_fd_sc_hd__nand3_4 _19247_ (.A(_09188_),
    .B(_09189_),
    .C(_09190_),
    .Y(_09195_));
 sky130_fd_sc_hd__a32oi_4 _19248_ (.A1(_08874_),
    .A2(_08880_),
    .A3(_08876_),
    .B1(_08836_),
    .B2(_08839_),
    .Y(_09197_));
 sky130_fd_sc_hd__o21ai_2 _19249_ (.A1(_08840_),
    .A2(_08882_),
    .B1(_08884_),
    .Y(_09198_));
 sky130_fd_sc_hd__a21oi_1 _19250_ (.A1(_09192_),
    .A2(_09195_),
    .B1(_09198_),
    .Y(_09199_));
 sky130_fd_sc_hd__o2bb2ai_2 _19251_ (.A1_N(_09192_),
    .A2_N(_09195_),
    .B1(_09197_),
    .B2(_08882_),
    .Y(_09200_));
 sky130_fd_sc_hd__nand2_2 _19252_ (.A(_09192_),
    .B(_09198_),
    .Y(_09201_));
 sky130_fd_sc_hd__and3_1 _19253_ (.A(_09192_),
    .B(_09195_),
    .C(_09198_),
    .X(_09202_));
 sky130_fd_sc_hd__a21boi_1 _19254_ (.A1(_09192_),
    .A2(_09195_),
    .B1_N(_09198_),
    .Y(_09203_));
 sky130_fd_sc_hd__a21bo_1 _19255_ (.A1(_09192_),
    .A2(_09195_),
    .B1_N(_09198_),
    .X(_09204_));
 sky130_fd_sc_hd__o211a_1 _19256_ (.A1(_08882_),
    .A2(_09197_),
    .B1(_09195_),
    .C1(_09192_),
    .X(_09205_));
 sky130_fd_sc_hd__o2111ai_2 _19257_ (.A1(_08840_),
    .A2(_08882_),
    .B1(_08884_),
    .C1(_09192_),
    .D1(_09195_),
    .Y(_09206_));
 sky130_fd_sc_hd__o21ai_2 _19258_ (.A1(_09194_),
    .A2(_09201_),
    .B1(_09200_),
    .Y(_09208_));
 sky130_fd_sc_hd__nand4_2 _19259_ (.A(_09110_),
    .B(_09112_),
    .C(_09204_),
    .D(_09206_),
    .Y(_09209_));
 sky130_fd_sc_hd__o2bb2ai_2 _19260_ (.A1_N(_09110_),
    .A2_N(_09112_),
    .B1(_09203_),
    .B2(_09205_),
    .Y(_09210_));
 sky130_fd_sc_hd__o2bb2ai_2 _19261_ (.A1_N(_09110_),
    .A2_N(_09112_),
    .B1(_09199_),
    .B2(_09202_),
    .Y(_09211_));
 sky130_fd_sc_hd__o2111ai_4 _19262_ (.A1(_09194_),
    .A2(_09201_),
    .B1(_09200_),
    .C1(_09110_),
    .D1(_09112_),
    .Y(_09212_));
 sky130_fd_sc_hd__nand3_2 _19263_ (.A(_09210_),
    .B(_08941_),
    .C(_09209_),
    .Y(_09213_));
 sky130_fd_sc_hd__and3_2 _19264_ (.A(_08942_),
    .B(_09211_),
    .C(_09212_),
    .X(_09214_));
 sky130_fd_sc_hd__nand3_1 _19265_ (.A(_08942_),
    .B(_09211_),
    .C(_09212_),
    .Y(_09215_));
 sky130_fd_sc_hd__and3_1 _19266_ (.A(_08577_),
    .B(_08584_),
    .C(_08894_),
    .X(_09216_));
 sky130_fd_sc_hd__a31o_1 _19267_ (.A1(_08810_),
    .A2(_08888_),
    .A3(_08890_),
    .B1(_08899_),
    .X(_09217_));
 sky130_fd_sc_hd__a31o_1 _19268_ (.A1(_08577_),
    .A2(_08584_),
    .A3(_08894_),
    .B1(_08891_),
    .X(_09219_));
 sky130_fd_sc_hd__o2bb2ai_2 _19269_ (.A1_N(_09213_),
    .A2_N(_09215_),
    .B1(_09216_),
    .B2(_08891_),
    .Y(_09220_));
 sky130_fd_sc_hd__a31oi_2 _19270_ (.A1(_09210_),
    .A2(_08941_),
    .A3(_09209_),
    .B1(_09219_),
    .Y(_09221_));
 sky130_fd_sc_hd__a31o_1 _19271_ (.A1(_09210_),
    .A2(_08941_),
    .A3(_09209_),
    .B1(_09219_),
    .X(_09222_));
 sky130_fd_sc_hd__o211ai_1 _19272_ (.A1(_08893_),
    .A2(_08899_),
    .B1(_09213_),
    .C1(_09215_),
    .Y(_09223_));
 sky130_fd_sc_hd__o2bb2ai_2 _19273_ (.A1_N(_08919_),
    .A2_N(_08917_),
    .B1(_08913_),
    .B2(_08907_),
    .Y(_09224_));
 sky130_fd_sc_hd__a21oi_1 _19274_ (.A1(_09220_),
    .A2(_09223_),
    .B1(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__a21o_1 _19275_ (.A1(_09220_),
    .A2(_09223_),
    .B1(_09224_),
    .X(_09226_));
 sky130_fd_sc_hd__o211a_1 _19276_ (.A1(_09214_),
    .A2(_09222_),
    .B1(_09224_),
    .C1(_09220_),
    .X(_09227_));
 sky130_fd_sc_hd__o211ai_2 _19277_ (.A1(_09214_),
    .A2(_09222_),
    .B1(_09224_),
    .C1(_09220_),
    .Y(_09228_));
 sky130_fd_sc_hd__o22ai_2 _19278_ (.A1(_08835_),
    .A2(_08838_),
    .B1(_09225_),
    .B2(_09227_),
    .Y(_09230_));
 sky130_fd_sc_hd__nand3_1 _19279_ (.A(_09226_),
    .B(_09228_),
    .C(_08940_),
    .Y(_09231_));
 sky130_fd_sc_hd__nand2_2 _19280_ (.A(_09230_),
    .B(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__a22oi_2 _19281_ (.A1(_08928_),
    .A2(_08932_),
    .B1(_09230_),
    .B2(_09231_),
    .Y(_09233_));
 sky130_fd_sc_hd__xor2_4 _19282_ (.A(_08939_),
    .B(_09232_),
    .X(_09234_));
 sky130_fd_sc_hd__o2111a_2 _19283_ (.A1(_08930_),
    .A2(_08936_),
    .B1(_08935_),
    .C1(_08625_),
    .D1(_08626_),
    .X(_09235_));
 sky130_fd_sc_hd__o2111ai_1 _19284_ (.A1(_08930_),
    .A2(_08936_),
    .B1(_08935_),
    .C1(_08625_),
    .D1(_08626_),
    .Y(_09236_));
 sky130_fd_sc_hd__nor2_1 _19285_ (.A(_08631_),
    .B(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand4_4 _19286_ (.A(_09235_),
    .B(_07984_),
    .C(_08324_),
    .D(_07985_),
    .Y(_09238_));
 sky130_fd_sc_hd__a221oi_4 _19287_ (.A1(_08628_),
    .A2(_08935_),
    .B1(_09235_),
    .B2(_08630_),
    .C1(_08937_),
    .Y(_09239_));
 sky130_fd_sc_hd__o21ai_4 _19288_ (.A1(_09238_),
    .A2(_07989_),
    .B1(_09239_),
    .Y(_09241_));
 sky130_fd_sc_hd__nand2_1 _19289_ (.A(_07990_),
    .B(_09237_),
    .Y(_09242_));
 sky130_fd_sc_hd__a31oi_4 _19290_ (.A1(_06596_),
    .A2(_06598_),
    .A3(_06600_),
    .B1(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__o21a_1 _19291_ (.A1(_09241_),
    .A2(_09243_),
    .B1(_09234_),
    .X(_09244_));
 sky130_fd_sc_hd__a311oi_2 _19292_ (.A1(_06601_),
    .A2(_07990_),
    .A3(_09237_),
    .B1(_09234_),
    .C1(_09241_),
    .Y(_09245_));
 sky130_fd_sc_hd__nor2_1 _19293_ (.A(_09244_),
    .B(_09245_),
    .Y(net99));
 sky130_fd_sc_hd__a32oi_4 _19294_ (.A1(_08942_),
    .A2(_09211_),
    .A3(_09212_),
    .B1(_09213_),
    .B2(_09217_),
    .Y(_09246_));
 sky130_fd_sc_hd__nand3_1 _19295_ (.A(_09110_),
    .B(_09204_),
    .C(_09206_),
    .Y(_09247_));
 sky130_fd_sc_hd__o211ai_2 _19296_ (.A1(_09194_),
    .A2(_09201_),
    .B1(_09200_),
    .C1(_09112_),
    .Y(_09248_));
 sky130_fd_sc_hd__o21ai_1 _19297_ (.A1(_09111_),
    .A2(_09208_),
    .B1(_09110_),
    .Y(_09249_));
 sky130_fd_sc_hd__o21ai_2 _19298_ (.A1(_09008_),
    .A2(_09006_),
    .B1(_09005_),
    .Y(_09251_));
 sky130_fd_sc_hd__o22a_1 _19299_ (.A1(_02043_),
    .A2(_02054_),
    .B1(_08723_),
    .B2(_09057_),
    .X(_09252_));
 sky130_fd_sc_hd__a21oi_2 _19300_ (.A1(_08723_),
    .A2(_09057_),
    .B1(_09056_),
    .Y(_09253_));
 sky130_fd_sc_hd__nand2_1 _19301_ (.A(net43),
    .B(net16),
    .Y(_09254_));
 sky130_fd_sc_hd__nand4_2 _19302_ (.A(net42),
    .B(net43),
    .C(net15),
    .D(net16),
    .Y(_09255_));
 sky130_fd_sc_hd__a22oi_4 _19303_ (.A1(net43),
    .A2(net15),
    .B1(net16),
    .B2(net42),
    .Y(_09256_));
 sky130_fd_sc_hd__a22o_2 _19304_ (.A1(net43),
    .A2(net15),
    .B1(net16),
    .B2(net42),
    .X(_09257_));
 sky130_fd_sc_hd__a2bb2oi_1 _19305_ (.A1_N(_02054_),
    .A2_N(_02065_),
    .B1(_09255_),
    .B2(_09257_),
    .Y(_09258_));
 sky130_fd_sc_hd__o2bb2ai_2 _19306_ (.A1_N(_09255_),
    .A2_N(_09257_),
    .B1(_02054_),
    .B2(_02065_),
    .Y(_09259_));
 sky130_fd_sc_hd__o2111a_2 _19307_ (.A1(_09057_),
    .A2(_09254_),
    .B1(net45),
    .C1(net14),
    .D1(_09257_),
    .X(_09260_));
 sky130_fd_sc_hd__o2111ai_2 _19308_ (.A1(_09057_),
    .A2(_09254_),
    .B1(net45),
    .C1(net14),
    .D1(_09257_),
    .Y(_09262_));
 sky130_fd_sc_hd__o22ai_4 _19309_ (.A1(_09060_),
    .A2(_09252_),
    .B1(_09258_),
    .B2(_09260_),
    .Y(_09263_));
 sky130_fd_sc_hd__o21ai_2 _19310_ (.A1(_09058_),
    .A2(_09253_),
    .B1(_09259_),
    .Y(_09264_));
 sky130_fd_sc_hd__o211a_1 _19311_ (.A1(_09058_),
    .A2(_09253_),
    .B1(_09259_),
    .C1(_09262_),
    .X(_09265_));
 sky130_fd_sc_hd__o211ai_2 _19312_ (.A1(_09058_),
    .A2(_09253_),
    .B1(_09259_),
    .C1(_09262_),
    .Y(_09266_));
 sky130_fd_sc_hd__nand2_1 _19313_ (.A(net13),
    .B(net46),
    .Y(_09267_));
 sky130_fd_sc_hd__a22o_2 _19314_ (.A1(net13),
    .A2(net46),
    .B1(net47),
    .B2(net11),
    .X(_09268_));
 sky130_fd_sc_hd__nand2_1 _19315_ (.A(net13),
    .B(net47),
    .Y(_09269_));
 sky130_fd_sc_hd__and4_2 _19316_ (.A(net11),
    .B(net13),
    .C(net46),
    .D(net47),
    .X(_09270_));
 sky130_fd_sc_hd__nand4_2 _19317_ (.A(net11),
    .B(net13),
    .C(net46),
    .D(net47),
    .Y(_09271_));
 sky130_fd_sc_hd__nand2_1 _19318_ (.A(net10),
    .B(net48),
    .Y(_09273_));
 sky130_fd_sc_hd__a22oi_4 _19319_ (.A1(net10),
    .A2(net48),
    .B1(_09268_),
    .B2(_09271_),
    .Y(_09274_));
 sky130_fd_sc_hd__a22o_1 _19320_ (.A1(net10),
    .A2(net48),
    .B1(_09268_),
    .B2(_09271_),
    .X(_09275_));
 sky130_fd_sc_hd__o2111a_1 _19321_ (.A1(_09073_),
    .A2(_09269_),
    .B1(net10),
    .C1(net48),
    .D1(_09268_),
    .X(_09276_));
 sky130_fd_sc_hd__or4b_1 _19322_ (.A(_02021_),
    .B(_09270_),
    .C(_02109_),
    .D_N(_09268_),
    .X(_09277_));
 sky130_fd_sc_hd__nor2_1 _19323_ (.A(_09274_),
    .B(_09276_),
    .Y(_09278_));
 sky130_fd_sc_hd__a211oi_1 _19324_ (.A1(_09263_),
    .A2(_09266_),
    .B1(_09274_),
    .C1(_09276_),
    .Y(_09279_));
 sky130_fd_sc_hd__a211o_1 _19325_ (.A1(_09263_),
    .A2(_09266_),
    .B1(_09274_),
    .C1(_09276_),
    .X(_09280_));
 sky130_fd_sc_hd__o221a_1 _19326_ (.A1(_09274_),
    .A2(_09276_),
    .B1(_09260_),
    .B2(_09264_),
    .C1(_09263_),
    .X(_09281_));
 sky130_fd_sc_hd__o221ai_2 _19327_ (.A1(_09274_),
    .A2(_09276_),
    .B1(_09260_),
    .B2(_09264_),
    .C1(_09263_),
    .Y(_09282_));
 sky130_fd_sc_hd__o2bb2a_1 _19328_ (.A1_N(_09263_),
    .A2_N(_09266_),
    .B1(_09274_),
    .B2(_09276_),
    .X(_09284_));
 sky130_fd_sc_hd__a22o_1 _19329_ (.A1(_09263_),
    .A2(_09266_),
    .B1(_09275_),
    .B2(_09277_),
    .X(_09285_));
 sky130_fd_sc_hd__nand2_1 _19330_ (.A(_09263_),
    .B(_09278_),
    .Y(_09286_));
 sky130_fd_sc_hd__and3_1 _19331_ (.A(_09263_),
    .B(_09278_),
    .C(_09266_),
    .X(_09287_));
 sky130_fd_sc_hd__o21ai_2 _19332_ (.A1(_09038_),
    .A2(_09041_),
    .B1(_09047_),
    .Y(_09288_));
 sky130_fd_sc_hd__o21a_1 _19333_ (.A1(_02010_),
    .A2(_02098_),
    .B1(_09034_),
    .X(_09289_));
 sky130_fd_sc_hd__and3_1 _19334_ (.A(_09032_),
    .B(net16),
    .C(net41),
    .X(_09290_));
 sky130_fd_sc_hd__a31o_1 _19335_ (.A1(_09032_),
    .A2(net16),
    .A3(net41),
    .B1(_09033_),
    .X(_09291_));
 sky130_fd_sc_hd__o31a_1 _19336_ (.A1(_02010_),
    .A2(_02098_),
    .A3(_09030_),
    .B1(_09034_),
    .X(_09292_));
 sky130_fd_sc_hd__nor2_1 _19337_ (.A(_08988_),
    .B(_08991_),
    .Y(_09293_));
 sky130_fd_sc_hd__o21ai_2 _19338_ (.A1(_08988_),
    .A2(_08991_),
    .B1(_08990_),
    .Y(_09295_));
 sky130_fd_sc_hd__o21a_1 _19339_ (.A1(_08988_),
    .A2(_08991_),
    .B1(_08990_),
    .X(_09296_));
 sky130_fd_sc_hd__nand2_2 _19340_ (.A(net41),
    .B(net17),
    .Y(_09297_));
 sky130_fd_sc_hd__nand2_2 _19341_ (.A(net39),
    .B(net19),
    .Y(_09298_));
 sky130_fd_sc_hd__a22oi_4 _19342_ (.A1(net40),
    .A2(net18),
    .B1(net19),
    .B2(net39),
    .Y(_09299_));
 sky130_fd_sc_hd__a22o_1 _19343_ (.A1(net40),
    .A2(net18),
    .B1(net19),
    .B2(net39),
    .X(_09300_));
 sky130_fd_sc_hd__nand2_1 _19344_ (.A(net40),
    .B(net19),
    .Y(_09301_));
 sky130_fd_sc_hd__and4_1 _19345_ (.A(net39),
    .B(net40),
    .C(net18),
    .D(net19),
    .X(_09302_));
 sky130_fd_sc_hd__nand4_4 _19346_ (.A(net39),
    .B(net40),
    .C(net18),
    .D(net19),
    .Y(_09303_));
 sky130_fd_sc_hd__nand3_4 _19347_ (.A(_09297_),
    .B(_09300_),
    .C(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__o21bai_4 _19348_ (.A1(_09299_),
    .A2(_09302_),
    .B1_N(_09297_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand4_2 _19349_ (.A(_09300_),
    .B(_09303_),
    .C(net41),
    .D(net17),
    .Y(_09307_));
 sky130_fd_sc_hd__o2bb2ai_2 _19350_ (.A1_N(net41),
    .A2_N(net17),
    .B1(_09299_),
    .B2(_09302_),
    .Y(_09308_));
 sky130_fd_sc_hd__a2bb2oi_4 _19351_ (.A1_N(_08989_),
    .A2_N(_09293_),
    .B1(_09304_),
    .B2(_09306_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand3_4 _19352_ (.A(_09308_),
    .B(_09295_),
    .C(_09307_),
    .Y(_09310_));
 sky130_fd_sc_hd__a21oi_2 _19353_ (.A1(_09307_),
    .A2(_09308_),
    .B1(_09295_),
    .Y(_09311_));
 sky130_fd_sc_hd__nand3_2 _19354_ (.A(_09296_),
    .B(_09304_),
    .C(_09306_),
    .Y(_09312_));
 sky130_fd_sc_hd__a31oi_4 _19355_ (.A1(_09296_),
    .A2(_09304_),
    .A3(_09306_),
    .B1(_09292_),
    .Y(_09313_));
 sky130_fd_sc_hd__o211a_1 _19356_ (.A1(_09033_),
    .A2(_09290_),
    .B1(_09310_),
    .C1(_09312_),
    .X(_09314_));
 sky130_fd_sc_hd__nand2_1 _19357_ (.A(_09313_),
    .B(_09310_),
    .Y(_09315_));
 sky130_fd_sc_hd__a2bb2oi_2 _19358_ (.A1_N(_09030_),
    .A2_N(_09289_),
    .B1(_09310_),
    .B2(_09312_),
    .Y(_09317_));
 sky130_fd_sc_hd__o22ai_4 _19359_ (.A1(_09030_),
    .A2(_09289_),
    .B1(_09309_),
    .B2(_09311_),
    .Y(_09318_));
 sky130_fd_sc_hd__a221oi_4 _19360_ (.A1(_09313_),
    .A2(_09310_),
    .B1(_09047_),
    .B2(_09043_),
    .C1(_09317_),
    .Y(_09319_));
 sky130_fd_sc_hd__nand3_2 _19361_ (.A(_09288_),
    .B(_09315_),
    .C(_09318_),
    .Y(_09320_));
 sky130_fd_sc_hd__a21oi_4 _19362_ (.A1(_09315_),
    .A2(_09318_),
    .B1(_09288_),
    .Y(_09321_));
 sky130_fd_sc_hd__o221ai_4 _19363_ (.A1(_09041_),
    .A2(_09038_),
    .B1(_09317_),
    .B2(_09314_),
    .C1(_09048_),
    .Y(_09322_));
 sky130_fd_sc_hd__o211a_2 _19364_ (.A1(_09286_),
    .A2(_09265_),
    .B1(_09285_),
    .C1(_09322_),
    .X(_09323_));
 sky130_fd_sc_hd__o2111ai_4 _19365_ (.A1(_09286_),
    .A2(_09265_),
    .B1(_09285_),
    .C1(_09320_),
    .D1(_09322_),
    .Y(_09324_));
 sky130_fd_sc_hd__o22ai_2 _19366_ (.A1(_09284_),
    .A2(_09287_),
    .B1(_09319_),
    .B2(_09321_),
    .Y(_09325_));
 sky130_fd_sc_hd__o22ai_2 _19367_ (.A1(_09279_),
    .A2(_09281_),
    .B1(_09319_),
    .B2(_09321_),
    .Y(_09326_));
 sky130_fd_sc_hd__o211ai_2 _19368_ (.A1(_09284_),
    .A2(_09287_),
    .B1(_09320_),
    .C1(_09322_),
    .Y(_09328_));
 sky130_fd_sc_hd__o211ai_4 _19369_ (.A1(_09006_),
    .A2(_09011_),
    .B1(_09324_),
    .C1(_09325_),
    .Y(_09329_));
 sky130_fd_sc_hd__nand3_4 _19370_ (.A(_09326_),
    .B(_09328_),
    .C(_09251_),
    .Y(_09330_));
 sky130_fd_sc_hd__and3_1 _19371_ (.A(_09054_),
    .B(_09082_),
    .C(_09084_),
    .X(_09331_));
 sky130_fd_sc_hd__o21ai_2 _19372_ (.A1(_09025_),
    .A2(_09049_),
    .B1(_09088_),
    .Y(_09332_));
 sky130_fd_sc_hd__o2bb2ai_4 _19373_ (.A1_N(_09329_),
    .A2_N(_09330_),
    .B1(_09331_),
    .B2(_09050_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_1 _19374_ (.A(_09330_),
    .B(_09332_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand3_4 _19375_ (.A(_09329_),
    .B(_09330_),
    .C(_09332_),
    .Y(_09335_));
 sky130_fd_sc_hd__a22oi_4 _19376_ (.A1(_08950_),
    .A2(_08966_),
    .B1(_09010_),
    .B2(_09013_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand3_2 _19377_ (.A(_08969_),
    .B(_09014_),
    .C(_09015_),
    .Y(_09337_));
 sky130_fd_sc_hd__a31oi_4 _19378_ (.A1(_08644_),
    .A2(_08649_),
    .A3(_07698_),
    .B1(_08953_),
    .Y(_09339_));
 sky130_fd_sc_hd__o211ai_4 _19379_ (.A1(_07699_),
    .A2(_08643_),
    .B1(_08646_),
    .C1(_08335_),
    .Y(_09340_));
 sky130_fd_sc_hd__o22ai_4 _19380_ (.A1(_08647_),
    .A2(_08653_),
    .B1(_08952_),
    .B2(_08651_),
    .Y(_09341_));
 sky130_fd_sc_hd__a31o_2 _19381_ (.A1(_08335_),
    .A2(_08646_),
    .A3(_08653_),
    .B1(_08651_),
    .X(_09342_));
 sky130_fd_sc_hd__o22ai_4 _19382_ (.A1(_02218_),
    .A2(_08979_),
    .B1(_08972_),
    .B2(_08974_),
    .Y(_09343_));
 sky130_fd_sc_hd__o22a_1 _19383_ (.A1(_02218_),
    .A2(_08979_),
    .B1(_08972_),
    .B2(_08974_),
    .X(_09344_));
 sky130_fd_sc_hd__and2_1 _19384_ (.A(net35),
    .B(net24),
    .X(_09345_));
 sky130_fd_sc_hd__o21a_4 _19385_ (.A1(net64),
    .A2(net34),
    .B1(net25),
    .X(_09346_));
 sky130_fd_sc_hd__o2bb2ai_1 _19386_ (.A1_N(_08973_),
    .A2_N(_08977_),
    .B1(_08978_),
    .B2(_02251_),
    .Y(_09347_));
 sky130_fd_sc_hd__o221ai_2 _19387_ (.A1(_01934_),
    .A2(_02218_),
    .B1(_02251_),
    .B2(_08978_),
    .C1(_09346_),
    .Y(_09348_));
 sky130_fd_sc_hd__nand2_1 _19388_ (.A(_09347_),
    .B(_09345_),
    .Y(_09350_));
 sky130_fd_sc_hd__o2bb2ai_2 _19389_ (.A1_N(_08979_),
    .A2_N(_09346_),
    .B1(_01934_),
    .B2(_02218_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand4_2 _19390_ (.A(_09346_),
    .B(net24),
    .C(net35),
    .D(_08979_),
    .Y(_09352_));
 sky130_fd_sc_hd__a21oi_1 _19391_ (.A1(_09351_),
    .A2(_09352_),
    .B1(_09343_),
    .Y(_09353_));
 sky130_fd_sc_hd__nand3_2 _19392_ (.A(_09344_),
    .B(_09348_),
    .C(_09350_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand3_4 _19393_ (.A(_09351_),
    .B(_09352_),
    .C(_09343_),
    .Y(_09355_));
 sky130_fd_sc_hd__nand2_1 _19394_ (.A(net38),
    .B(net20),
    .Y(_09356_));
 sky130_fd_sc_hd__nand2_1 _19395_ (.A(net37),
    .B(net22),
    .Y(_09357_));
 sky130_fd_sc_hd__and4_1 _19396_ (.A(net36),
    .B(net37),
    .C(net21),
    .D(net22),
    .X(_09358_));
 sky130_fd_sc_hd__nand4_4 _19397_ (.A(net36),
    .B(net37),
    .C(net21),
    .D(net22),
    .Y(_09359_));
 sky130_fd_sc_hd__a22oi_2 _19398_ (.A1(net37),
    .A2(net21),
    .B1(net22),
    .B2(net36),
    .Y(_09361_));
 sky130_fd_sc_hd__a22o_1 _19399_ (.A1(net37),
    .A2(net21),
    .B1(net22),
    .B2(net36),
    .X(_09362_));
 sky130_fd_sc_hd__and3_1 _19400_ (.A(_09356_),
    .B(_09359_),
    .C(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__o211a_1 _19401_ (.A1(_09358_),
    .A2(_09361_),
    .B1(net38),
    .C1(net20),
    .X(_09364_));
 sky130_fd_sc_hd__o2bb2a_1 _19402_ (.A1_N(net38),
    .A2_N(net20),
    .B1(_09358_),
    .B2(_09361_),
    .X(_09365_));
 sky130_fd_sc_hd__a22o_1 _19403_ (.A1(net38),
    .A2(net20),
    .B1(_09359_),
    .B2(_09362_),
    .X(_09366_));
 sky130_fd_sc_hd__and4_1 _19404_ (.A(_09362_),
    .B(net20),
    .C(net38),
    .D(_09359_),
    .X(_09367_));
 sky130_fd_sc_hd__nand4_1 _19405_ (.A(_09362_),
    .B(net20),
    .C(net38),
    .D(_09359_),
    .Y(_09368_));
 sky130_fd_sc_hd__nand2_1 _19406_ (.A(_09366_),
    .B(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__o2bb2ai_1 _19407_ (.A1_N(_09354_),
    .A2_N(_09355_),
    .B1(_09363_),
    .B2(_09364_),
    .Y(_09370_));
 sky130_fd_sc_hd__o211ai_2 _19408_ (.A1(_09365_),
    .A2(_09367_),
    .B1(_09354_),
    .C1(_09355_),
    .Y(_09372_));
 sky130_fd_sc_hd__o2bb2ai_2 _19409_ (.A1_N(_09354_),
    .A2_N(_09355_),
    .B1(_09365_),
    .B2(_09367_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand4_2 _19410_ (.A(_09354_),
    .B(_09355_),
    .C(_09366_),
    .D(_09368_),
    .Y(_09374_));
 sky130_fd_sc_hd__nand2_1 _19411_ (.A(_09373_),
    .B(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__nand3_4 _19412_ (.A(_09342_),
    .B(_09370_),
    .C(_09372_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand3_4 _19413_ (.A(_09373_),
    .B(_09374_),
    .C(_09341_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand2_4 _19414_ (.A(_08985_),
    .B(_09001_),
    .Y(_09378_));
 sky130_fd_sc_hd__a21oi_2 _19415_ (.A1(_09376_),
    .A2(_09377_),
    .B1(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__a21o_1 _19416_ (.A1(_09376_),
    .A2(_09377_),
    .B1(_09378_),
    .X(_09380_));
 sky130_fd_sc_hd__nand3_4 _19417_ (.A(_09376_),
    .B(_09377_),
    .C(_09378_),
    .Y(_09381_));
 sky130_fd_sc_hd__a21oi_4 _19418_ (.A1(_08955_),
    .A2(_08956_),
    .B1(_08004_),
    .Y(_09383_));
 sky130_fd_sc_hd__a21o_4 _19419_ (.A1(_08955_),
    .A2(_08956_),
    .B1(_08004_),
    .X(_09384_));
 sky130_fd_sc_hd__and3_4 _19420_ (.A(_08955_),
    .B(_08956_),
    .C(_08006_),
    .X(_09385_));
 sky130_fd_sc_hd__nand3_4 _19421_ (.A(_08955_),
    .B(_08956_),
    .C(_08006_),
    .Y(_09386_));
 sky130_fd_sc_hd__o21a_2 _19422_ (.A1(_08004_),
    .A2(_08959_),
    .B1(_09386_),
    .X(_09387_));
 sky130_fd_sc_hd__o21ai_2 _19423_ (.A1(_08004_),
    .A2(_08959_),
    .B1(_09386_),
    .Y(_09388_));
 sky130_fd_sc_hd__a21oi_4 _19424_ (.A1(_09380_),
    .A2(_09381_),
    .B1(_09387_),
    .Y(_09389_));
 sky130_fd_sc_hd__a21o_1 _19425_ (.A1(_09380_),
    .A2(_09381_),
    .B1(_09387_),
    .X(_09390_));
 sky130_fd_sc_hd__a31o_1 _19426_ (.A1(_09376_),
    .A2(_09377_),
    .A3(_09378_),
    .B1(_09383_),
    .X(_09391_));
 sky130_fd_sc_hd__nor3_2 _19427_ (.A(_09379_),
    .B(_09385_),
    .C(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__nand3_2 _19428_ (.A(_09380_),
    .B(_09381_),
    .C(_09387_),
    .Y(_09394_));
 sky130_fd_sc_hd__o211ai_4 _19429_ (.A1(_08966_),
    .A2(_08950_),
    .B1(_09394_),
    .C1(_09337_),
    .Y(_09395_));
 sky130_fd_sc_hd__nor2_1 _19430_ (.A(_09389_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__nand4_2 _19431_ (.A(_08968_),
    .B(_09337_),
    .C(_09390_),
    .D(_09394_),
    .Y(_09397_));
 sky130_fd_sc_hd__o22a_2 _19432_ (.A1(_08967_),
    .A2(_09336_),
    .B1(_09389_),
    .B2(_09392_),
    .X(_09398_));
 sky130_fd_sc_hd__o22ai_4 _19433_ (.A1(_08967_),
    .A2(_09336_),
    .B1(_09389_),
    .B2(_09392_),
    .Y(_09399_));
 sky130_fd_sc_hd__a22oi_4 _19434_ (.A1(_09333_),
    .A2(_09335_),
    .B1(_09397_),
    .B2(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__o2111a_1 _19435_ (.A1(_09395_),
    .A2(_09389_),
    .B1(_09335_),
    .C1(_09333_),
    .D1(_09399_),
    .X(_09401_));
 sky130_fd_sc_hd__o2111ai_4 _19436_ (.A1(_09395_),
    .A2(_09389_),
    .B1(_09335_),
    .C1(_09333_),
    .D1(_09399_),
    .Y(_09402_));
 sky130_fd_sc_hd__a2bb2oi_2 _19437_ (.A1_N(_09395_),
    .A2_N(_09389_),
    .B1(_09335_),
    .B2(_09333_),
    .Y(_09403_));
 sky130_fd_sc_hd__a2bb2o_1 _19438_ (.A1_N(_09395_),
    .A2_N(_09389_),
    .B1(_09335_),
    .B2(_09333_),
    .X(_09405_));
 sky130_fd_sc_hd__a31oi_4 _19439_ (.A1(_09333_),
    .A2(_09335_),
    .A3(_09399_),
    .B1(_09396_),
    .Y(_09406_));
 sky130_fd_sc_hd__a31oi_2 _19440_ (.A1(_09019_),
    .A2(_09102_),
    .A3(_09104_),
    .B1(_09021_),
    .Y(_09407_));
 sky130_fd_sc_hd__a31o_1 _19441_ (.A1(_09019_),
    .A2(_09102_),
    .A3(_09104_),
    .B1(_09021_),
    .X(_09408_));
 sky130_fd_sc_hd__o21ai_4 _19442_ (.A1(_09400_),
    .A2(_09401_),
    .B1(_09408_),
    .Y(_09409_));
 sky130_fd_sc_hd__nand3b_4 _19443_ (.A_N(_09400_),
    .B(_09407_),
    .C(_09402_),
    .Y(_09410_));
 sky130_fd_sc_hd__a32oi_4 _19444_ (.A1(_09091_),
    .A2(_09023_),
    .A3(_08702_),
    .B1(_09094_),
    .B2(_09092_),
    .Y(_09411_));
 sky130_fd_sc_hd__a21boi_2 _19445_ (.A1(_09093_),
    .A2(_09095_),
    .B1_N(_09092_),
    .Y(_09412_));
 sky130_fd_sc_hd__a21o_1 _19446_ (.A1(_09125_),
    .A2(_09132_),
    .B1(_09126_),
    .X(_09413_));
 sky130_fd_sc_hd__o21a_1 _19447_ (.A1(_01923_),
    .A2(_02207_),
    .B1(_09120_),
    .X(_09414_));
 sky130_fd_sc_hd__o21ai_1 _19448_ (.A1(_09115_),
    .A2(_09116_),
    .B1(_09120_),
    .Y(_09416_));
 sky130_fd_sc_hd__nand2_1 _19449_ (.A(net6),
    .B(net52),
    .Y(_09417_));
 sky130_fd_sc_hd__a22o_2 _19450_ (.A1(net6),
    .A2(net52),
    .B1(net53),
    .B2(net5),
    .X(_09418_));
 sky130_fd_sc_hd__and4_1 _19451_ (.A(net5),
    .B(net6),
    .C(net52),
    .D(net53),
    .X(_09419_));
 sky130_fd_sc_hd__nand4_4 _19452_ (.A(net5),
    .B(net6),
    .C(net52),
    .D(net53),
    .Y(_09420_));
 sky130_fd_sc_hd__a22oi_2 _19453_ (.A1(net4),
    .A2(net54),
    .B1(_09418_),
    .B2(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__a22o_1 _19454_ (.A1(net4),
    .A2(net54),
    .B1(_09418_),
    .B2(_09420_),
    .X(_09422_));
 sky130_fd_sc_hd__and4_2 _19455_ (.A(_09418_),
    .B(_09420_),
    .C(net4),
    .D(net54),
    .X(_09423_));
 sky130_fd_sc_hd__nand4_1 _19456_ (.A(_09418_),
    .B(_09420_),
    .C(net4),
    .D(net54),
    .Y(_09424_));
 sky130_fd_sc_hd__o22ai_4 _19457_ (.A1(_09116_),
    .A2(_09414_),
    .B1(_09421_),
    .B2(_09423_),
    .Y(_09425_));
 sky130_fd_sc_hd__nand2_1 _19458_ (.A(_09422_),
    .B(_09416_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand3_1 _19459_ (.A(_09422_),
    .B(_09424_),
    .C(_09416_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand2_1 _19460_ (.A(net3),
    .B(net56),
    .Y(_09429_));
 sky130_fd_sc_hd__and4_2 _19461_ (.A(_01901_),
    .B(net3),
    .C(net56),
    .D(net57),
    .X(_09430_));
 sky130_fd_sc_hd__o22a_1 _19462_ (.A1(net2),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01923_),
    .X(_09431_));
 sky130_fd_sc_hd__nor2_1 _19463_ (.A(_09430_),
    .B(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__o2bb2ai_2 _19464_ (.A1_N(_09425_),
    .A2_N(_09428_),
    .B1(_09430_),
    .B2(_09431_),
    .Y(_09433_));
 sky130_fd_sc_hd__o211ai_2 _19465_ (.A1(_09423_),
    .A2(_09427_),
    .B1(_09432_),
    .C1(_09425_),
    .Y(_09434_));
 sky130_fd_sc_hd__nand3_2 _19466_ (.A(_09413_),
    .B(_09433_),
    .C(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__a21oi_1 _19467_ (.A1(_09433_),
    .A2(_09434_),
    .B1(_09413_),
    .Y(_09436_));
 sky130_fd_sc_hd__a21o_1 _19468_ (.A1(_09433_),
    .A2(_09434_),
    .B1(_09413_),
    .X(_09438_));
 sky130_fd_sc_hd__and3_2 _19469_ (.A(_09438_),
    .B(_09129_),
    .C(_09435_),
    .X(_09439_));
 sky130_fd_sc_hd__a21oi_2 _19470_ (.A1(_09435_),
    .A2(_09438_),
    .B1(_09129_),
    .Y(_09440_));
 sky130_fd_sc_hd__o311a_1 _19471_ (.A1(_01901_),
    .A2(_02229_),
    .A3(_09128_),
    .B1(_09435_),
    .C1(_09438_),
    .X(_09441_));
 sky130_fd_sc_hd__a21boi_2 _19472_ (.A1(_09435_),
    .A2(_09438_),
    .B1_N(_09129_),
    .Y(_09442_));
 sky130_fd_sc_hd__a21oi_2 _19473_ (.A1(_09154_),
    .A2(_09158_),
    .B1(_09156_),
    .Y(_09443_));
 sky130_fd_sc_hd__nand2_1 _19474_ (.A(_09155_),
    .B(_09160_),
    .Y(_09444_));
 sky130_fd_sc_hd__a31o_1 _19475_ (.A1(_09077_),
    .A2(net48),
    .A3(net9),
    .B1(_09074_),
    .X(_09445_));
 sky130_fd_sc_hd__a31oi_2 _19476_ (.A1(_09077_),
    .A2(net48),
    .A3(net9),
    .B1(_09074_),
    .Y(_09446_));
 sky130_fd_sc_hd__nand2_1 _19477_ (.A(net7),
    .B(net51),
    .Y(_09447_));
 sky130_fd_sc_hd__nand2_1 _19478_ (.A(net9),
    .B(net49),
    .Y(_09449_));
 sky130_fd_sc_hd__a22oi_4 _19479_ (.A1(net9),
    .A2(net49),
    .B1(net50),
    .B2(net8),
    .Y(_09450_));
 sky130_fd_sc_hd__nand2_2 _19480_ (.A(_09146_),
    .B(_09449_),
    .Y(_09451_));
 sky130_fd_sc_hd__and4_2 _19481_ (.A(net8),
    .B(net9),
    .C(net49),
    .D(net50),
    .X(_09452_));
 sky130_fd_sc_hd__nand4_4 _19482_ (.A(net8),
    .B(net9),
    .C(net49),
    .D(net50),
    .Y(_09453_));
 sky130_fd_sc_hd__o211ai_2 _19483_ (.A1(_01977_),
    .A2(_02152_),
    .B1(_09451_),
    .C1(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__o21bai_4 _19484_ (.A1(_09450_),
    .A2(_09452_),
    .B1_N(_09447_),
    .Y(_09455_));
 sky130_fd_sc_hd__a22o_1 _19485_ (.A1(net7),
    .A2(net51),
    .B1(_09451_),
    .B2(_09453_),
    .X(_09456_));
 sky130_fd_sc_hd__nand4_2 _19486_ (.A(_09451_),
    .B(_09453_),
    .C(net7),
    .D(net51),
    .Y(_09457_));
 sky130_fd_sc_hd__nand3_4 _19487_ (.A(_09446_),
    .B(_09454_),
    .C(_09455_),
    .Y(_09458_));
 sky130_fd_sc_hd__and3_1 _19488_ (.A(_09445_),
    .B(_09456_),
    .C(_09457_),
    .X(_09460_));
 sky130_fd_sc_hd__nand3_4 _19489_ (.A(_09445_),
    .B(_09456_),
    .C(_09457_),
    .Y(_09461_));
 sky130_fd_sc_hd__o32a_1 _19490_ (.A1(_01977_),
    .A2(_02120_),
    .A3(_09146_),
    .B1(_02152_),
    .B2(_01966_),
    .X(_09462_));
 sky130_fd_sc_hd__a31o_1 _19491_ (.A1(_09145_),
    .A2(net51),
    .A3(net6),
    .B1(_09147_),
    .X(_09463_));
 sky130_fd_sc_hd__o2bb2ai_4 _19492_ (.A1_N(_09458_),
    .A2_N(_09461_),
    .B1(_09462_),
    .B2(_09144_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand2_1 _19493_ (.A(_09458_),
    .B(_09463_),
    .Y(_09465_));
 sky130_fd_sc_hd__nand3_4 _19494_ (.A(_09458_),
    .B(_09461_),
    .C(_09463_),
    .Y(_09466_));
 sky130_fd_sc_hd__o22ai_4 _19495_ (.A1(_09065_),
    .A2(_09069_),
    .B1(_09080_),
    .B2(_09067_),
    .Y(_09467_));
 sky130_fd_sc_hd__a21oi_4 _19496_ (.A1(_09464_),
    .A2(_09466_),
    .B1(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__a21o_1 _19497_ (.A1(_09464_),
    .A2(_09466_),
    .B1(_09467_),
    .X(_09469_));
 sky130_fd_sc_hd__o211a_1 _19498_ (.A1(_09465_),
    .A2(_09460_),
    .B1(_09464_),
    .C1(_09467_),
    .X(_09471_));
 sky130_fd_sc_hd__o211ai_4 _19499_ (.A1(_09465_),
    .A2(_09460_),
    .B1(_09464_),
    .C1(_09467_),
    .Y(_09472_));
 sky130_fd_sc_hd__o211ai_2 _19500_ (.A1(_09156_),
    .A2(_09161_),
    .B1(_09469_),
    .C1(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__o21ai_2 _19501_ (.A1(_09468_),
    .A2(_09471_),
    .B1(_09443_),
    .Y(_09474_));
 sky130_fd_sc_hd__nand3_2 _19502_ (.A(_09469_),
    .B(_09472_),
    .C(_09443_),
    .Y(_09475_));
 sky130_fd_sc_hd__o22ai_2 _19503_ (.A1(_09156_),
    .A2(_09161_),
    .B1(_09468_),
    .B2(_09471_),
    .Y(_09476_));
 sky130_fd_sc_hd__o2111a_2 _19504_ (.A1(_09171_),
    .A2(_09167_),
    .B1(_09170_),
    .C1(_09475_),
    .D1(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__o2111ai_4 _19505_ (.A1(_09171_),
    .A2(_09167_),
    .B1(_09170_),
    .C1(_09475_),
    .D1(_09476_),
    .Y(_09478_));
 sky130_fd_sc_hd__o211a_2 _19506_ (.A1(_09169_),
    .A2(_09172_),
    .B1(_09473_),
    .C1(_09474_),
    .X(_09479_));
 sky130_fd_sc_hd__o211ai_4 _19507_ (.A1(_09169_),
    .A2(_09172_),
    .B1(_09473_),
    .C1(_09474_),
    .Y(_09480_));
 sky130_fd_sc_hd__o21ai_1 _19508_ (.A1(_09441_),
    .A2(_09442_),
    .B1(_09480_),
    .Y(_09482_));
 sky130_fd_sc_hd__o211a_2 _19509_ (.A1(_09441_),
    .A2(_09442_),
    .B1(_09478_),
    .C1(_09480_),
    .X(_09483_));
 sky130_fd_sc_hd__o22ai_2 _19510_ (.A1(_09439_),
    .A2(_09440_),
    .B1(_09477_),
    .B2(_09479_),
    .Y(_09484_));
 sky130_fd_sc_hd__o22ai_2 _19511_ (.A1(_09441_),
    .A2(_09442_),
    .B1(_09477_),
    .B2(_09479_),
    .Y(_09485_));
 sky130_fd_sc_hd__o211ai_2 _19512_ (.A1(_09439_),
    .A2(_09440_),
    .B1(_09478_),
    .C1(_09480_),
    .Y(_09486_));
 sky130_fd_sc_hd__o211ai_4 _19513_ (.A1(_09482_),
    .A2(_09477_),
    .B1(_09412_),
    .C1(_09484_),
    .Y(_09487_));
 sky130_fd_sc_hd__nand3_4 _19514_ (.A(_09485_),
    .B(_09486_),
    .C(_09411_),
    .Y(_09488_));
 sky130_fd_sc_hd__inv_2 _19515_ (.A(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__a21oi_1 _19516_ (.A1(_09487_),
    .A2(_09488_),
    .B1(_09184_),
    .Y(_09490_));
 sky130_fd_sc_hd__a21o_1 _19517_ (.A1(_09487_),
    .A2(_09488_),
    .B1(_09184_),
    .X(_09491_));
 sky130_fd_sc_hd__and3_1 _19518_ (.A(_09487_),
    .B(_09488_),
    .C(_09184_),
    .X(_09493_));
 sky130_fd_sc_hd__nand3_1 _19519_ (.A(_09487_),
    .B(_09488_),
    .C(_09184_),
    .Y(_09494_));
 sky130_fd_sc_hd__a21boi_1 _19520_ (.A1(_09487_),
    .A2(_09488_),
    .B1_N(_09184_),
    .Y(_09495_));
 sky130_fd_sc_hd__a21bo_1 _19521_ (.A1(_09487_),
    .A2(_09488_),
    .B1_N(_09184_),
    .X(_09496_));
 sky130_fd_sc_hd__o2111a_1 _19522_ (.A1(_09182_),
    .A2(_09139_),
    .B1(_09181_),
    .C1(_09487_),
    .D1(_09488_),
    .X(_09497_));
 sky130_fd_sc_hd__o2111ai_4 _19523_ (.A1(_09182_),
    .A2(_09139_),
    .B1(_09181_),
    .C1(_09487_),
    .D1(_09488_),
    .Y(_09498_));
 sky130_fd_sc_hd__o2bb2ai_2 _19524_ (.A1_N(_09409_),
    .A2_N(_09410_),
    .B1(_09495_),
    .B2(_09497_),
    .Y(_09499_));
 sky130_fd_sc_hd__nand4_4 _19525_ (.A(_09409_),
    .B(_09410_),
    .C(_09496_),
    .D(_09498_),
    .Y(_09500_));
 sky130_fd_sc_hd__o2bb2ai_1 _19526_ (.A1_N(_09409_),
    .A2_N(_09410_),
    .B1(_09490_),
    .B2(_09493_),
    .Y(_09501_));
 sky130_fd_sc_hd__nand4_1 _19527_ (.A(_09409_),
    .B(_09410_),
    .C(_09491_),
    .D(_09494_),
    .Y(_09502_));
 sky130_fd_sc_hd__a22oi_4 _19528_ (.A1(_09110_),
    .A2(_09248_),
    .B1(_09499_),
    .B2(_09500_),
    .Y(_09504_));
 sky130_fd_sc_hd__nand3_1 _19529_ (.A(_09249_),
    .B(_09501_),
    .C(_09502_),
    .Y(_09505_));
 sky130_fd_sc_hd__a22oi_2 _19530_ (.A1(_09112_),
    .A2(_09247_),
    .B1(_09501_),
    .B2(_09502_),
    .Y(_09506_));
 sky130_fd_sc_hd__o2111ai_4 _19531_ (.A1(_09208_),
    .A2(_09111_),
    .B1(_09110_),
    .C1(_09500_),
    .D1(_09499_),
    .Y(_09507_));
 sky130_fd_sc_hd__o211a_1 _19532_ (.A1(_08840_),
    .A2(_08882_),
    .B1(_08884_),
    .C1(_09195_),
    .X(_09508_));
 sky130_fd_sc_hd__a21o_1 _19533_ (.A1(_09192_),
    .A2(_09198_),
    .B1(_09194_),
    .X(_09509_));
 sky130_fd_sc_hd__o31a_1 _19534_ (.A1(_08882_),
    .A2(_09193_),
    .A3(_09197_),
    .B1(_09195_),
    .X(_09510_));
 sky130_fd_sc_hd__o22ai_2 _19535_ (.A1(_09194_),
    .A2(_09202_),
    .B1(_09504_),
    .B2(_09506_),
    .Y(_09511_));
 sky130_fd_sc_hd__o211ai_2 _19536_ (.A1(_09193_),
    .A2(_09508_),
    .B1(_09507_),
    .C1(_09505_),
    .Y(_09512_));
 sky130_fd_sc_hd__o2bb2ai_1 _19537_ (.A1_N(_09505_),
    .A2_N(_09507_),
    .B1(_09508_),
    .B2(_09193_),
    .Y(_09513_));
 sky130_fd_sc_hd__o21ai_1 _19538_ (.A1(_09194_),
    .A2(_09202_),
    .B1(_09507_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand3_1 _19539_ (.A(_09511_),
    .B(_09512_),
    .C(_09246_),
    .Y(_09516_));
 sky130_fd_sc_hd__o221a_2 _19540_ (.A1(_09214_),
    .A2(_09221_),
    .B1(_09504_),
    .B2(_09515_),
    .C1(_09513_),
    .X(_09517_));
 sky130_fd_sc_hd__o221ai_2 _19541_ (.A1(_09214_),
    .A2(_09221_),
    .B1(_09504_),
    .B2(_09515_),
    .C1(_09513_),
    .Y(_09518_));
 sky130_fd_sc_hd__nor2_1 _19542_ (.A(_08827_),
    .B(_09136_),
    .Y(_09519_));
 sky130_fd_sc_hd__nor2_1 _19543_ (.A(_09135_),
    .B(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__inv_2 _19544_ (.A(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__o2bb2ai_1 _19545_ (.A1_N(_09516_),
    .A2_N(_09518_),
    .B1(_09519_),
    .B2(_09135_),
    .Y(_09522_));
 sky130_fd_sc_hd__a31oi_2 _19546_ (.A1(_09511_),
    .A2(_09512_),
    .A3(_09246_),
    .B1(_09521_),
    .Y(_09523_));
 sky130_fd_sc_hd__a31o_1 _19547_ (.A1(_09511_),
    .A2(_09512_),
    .A3(_09246_),
    .B1(_09521_),
    .X(_09524_));
 sky130_fd_sc_hd__nand3_1 _19548_ (.A(_09516_),
    .B(_09518_),
    .C(_09520_),
    .Y(_09526_));
 sky130_fd_sc_hd__o21ai_2 _19549_ (.A1(_08940_),
    .A2(_09225_),
    .B1(_09228_),
    .Y(_09527_));
 sky130_fd_sc_hd__a21oi_2 _19550_ (.A1(_09522_),
    .A2(_09526_),
    .B1(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__o211a_1 _19551_ (.A1(_09517_),
    .A2(_09524_),
    .B1(_09522_),
    .C1(_09527_),
    .X(_09529_));
 sky130_fd_sc_hd__nor2_2 _19552_ (.A(_09528_),
    .B(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__a21oi_1 _19553_ (.A1(_08939_),
    .A2(_09232_),
    .B1(_09244_),
    .Y(_09531_));
 sky130_fd_sc_hd__xnor2_1 _19554_ (.A(_09530_),
    .B(_09531_),
    .Y(net100));
 sky130_fd_sc_hd__nand3_4 _19555_ (.A(_09410_),
    .B(_09496_),
    .C(_09498_),
    .Y(_09532_));
 sky130_fd_sc_hd__o21ai_4 _19556_ (.A1(_09439_),
    .A2(_09440_),
    .B1(_09480_),
    .Y(_09533_));
 sky130_fd_sc_hd__a21boi_1 _19557_ (.A1(_09330_),
    .A2(_09332_),
    .B1_N(_09329_),
    .Y(_09534_));
 sky130_fd_sc_hd__nand2_1 _19558_ (.A(_09329_),
    .B(_09334_),
    .Y(_09536_));
 sky130_fd_sc_hd__a21o_2 _19559_ (.A1(_09458_),
    .A2(_09463_),
    .B1(_09460_),
    .X(_09537_));
 sky130_fd_sc_hd__a2bb2oi_1 _19560_ (.A1_N(_09260_),
    .A2_N(_09264_),
    .B1(_09278_),
    .B2(_09263_),
    .Y(_09538_));
 sky130_fd_sc_hd__o2bb2ai_2 _19561_ (.A1_N(_09278_),
    .A2_N(_09263_),
    .B1(_09260_),
    .B2(_09264_),
    .Y(_09539_));
 sky130_fd_sc_hd__o32a_1 _19562_ (.A1(_01999_),
    .A2(_02120_),
    .A3(_09146_),
    .B1(_02152_),
    .B2(_01977_),
    .X(_09540_));
 sky130_fd_sc_hd__and3_1 _19563_ (.A(_09451_),
    .B(net51),
    .C(net7),
    .X(_09541_));
 sky130_fd_sc_hd__a21oi_2 _19564_ (.A1(_09072_),
    .A2(_09267_),
    .B1(_09273_),
    .Y(_09542_));
 sky130_fd_sc_hd__a31o_1 _19565_ (.A1(_09268_),
    .A2(net48),
    .A3(net10),
    .B1(_09270_),
    .X(_09543_));
 sky130_fd_sc_hd__nor2_1 _19566_ (.A(_09270_),
    .B(_09542_),
    .Y(_09544_));
 sky130_fd_sc_hd__a22oi_4 _19567_ (.A1(net10),
    .A2(net49),
    .B1(net50),
    .B2(net9),
    .Y(_09545_));
 sky130_fd_sc_hd__a22o_2 _19568_ (.A1(net10),
    .A2(net49),
    .B1(net50),
    .B2(net9),
    .X(_09547_));
 sky130_fd_sc_hd__and4_1 _19569_ (.A(net9),
    .B(net10),
    .C(net49),
    .D(net50),
    .X(_09548_));
 sky130_fd_sc_hd__nand4_4 _19570_ (.A(net9),
    .B(net10),
    .C(net49),
    .D(net50),
    .Y(_09549_));
 sky130_fd_sc_hd__o211ai_1 _19571_ (.A1(_01988_),
    .A2(_02152_),
    .B1(_09547_),
    .C1(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__o211ai_1 _19572_ (.A1(_09545_),
    .A2(_09548_),
    .B1(net8),
    .C1(net51),
    .Y(_09551_));
 sky130_fd_sc_hd__nand4_4 _19573_ (.A(_09547_),
    .B(_09549_),
    .C(net8),
    .D(net51),
    .Y(_09552_));
 sky130_fd_sc_hd__o22ai_4 _19574_ (.A1(_01988_),
    .A2(_02152_),
    .B1(_09545_),
    .B2(_09548_),
    .Y(_09553_));
 sky130_fd_sc_hd__o211a_4 _19575_ (.A1(_09270_),
    .A2(_09542_),
    .B1(_09552_),
    .C1(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__o211ai_4 _19576_ (.A1(_09270_),
    .A2(_09542_),
    .B1(_09552_),
    .C1(_09553_),
    .Y(_09555_));
 sky130_fd_sc_hd__a21oi_2 _19577_ (.A1(_09552_),
    .A2(_09553_),
    .B1(_09543_),
    .Y(_09556_));
 sky130_fd_sc_hd__nand3_2 _19578_ (.A(_09544_),
    .B(_09550_),
    .C(_09551_),
    .Y(_09558_));
 sky130_fd_sc_hd__o21a_1 _19579_ (.A1(_09452_),
    .A2(_09541_),
    .B1(_09558_),
    .X(_09559_));
 sky130_fd_sc_hd__o21ai_4 _19580_ (.A1(_09452_),
    .A2(_09541_),
    .B1(_09558_),
    .Y(_09560_));
 sky130_fd_sc_hd__o22ai_2 _19581_ (.A1(_09450_),
    .A2(_09540_),
    .B1(_09554_),
    .B2(_09556_),
    .Y(_09561_));
 sky130_fd_sc_hd__o2111ai_4 _19582_ (.A1(_09447_),
    .A2(_09450_),
    .B1(_09453_),
    .C1(_09555_),
    .D1(_09558_),
    .Y(_09562_));
 sky130_fd_sc_hd__o22ai_2 _19583_ (.A1(_09452_),
    .A2(_09541_),
    .B1(_09554_),
    .B2(_09556_),
    .Y(_09563_));
 sky130_fd_sc_hd__o211a_1 _19584_ (.A1(_09554_),
    .A2(_09560_),
    .B1(_09561_),
    .C1(_09539_),
    .X(_09564_));
 sky130_fd_sc_hd__o211ai_4 _19585_ (.A1(_09554_),
    .A2(_09560_),
    .B1(_09561_),
    .C1(_09539_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand3_4 _19586_ (.A(_09563_),
    .B(_09538_),
    .C(_09562_),
    .Y(_09566_));
 sky130_fd_sc_hd__nand3_1 _19587_ (.A(_09537_),
    .B(_09565_),
    .C(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__a21o_1 _19588_ (.A1(_09565_),
    .A2(_09566_),
    .B1(_09537_),
    .X(_09569_));
 sky130_fd_sc_hd__a22o_1 _19589_ (.A1(_09461_),
    .A2(_09466_),
    .B1(_09565_),
    .B2(_09566_),
    .X(_09570_));
 sky130_fd_sc_hd__nand4_2 _19590_ (.A(_09461_),
    .B(_09466_),
    .C(_09565_),
    .D(_09566_),
    .Y(_09571_));
 sky130_fd_sc_hd__a31oi_2 _19591_ (.A1(_09464_),
    .A2(_09466_),
    .A3(_09467_),
    .B1(_09444_),
    .Y(_09572_));
 sky130_fd_sc_hd__o21ai_2 _19592_ (.A1(_09443_),
    .A2(_09468_),
    .B1(_09472_),
    .Y(_09573_));
 sky130_fd_sc_hd__o211a_1 _19593_ (.A1(_09468_),
    .A2(_09572_),
    .B1(_09571_),
    .C1(_09570_),
    .X(_09574_));
 sky130_fd_sc_hd__o211ai_4 _19594_ (.A1(_09468_),
    .A2(_09572_),
    .B1(_09571_),
    .C1(_09570_),
    .Y(_09575_));
 sky130_fd_sc_hd__nand3_4 _19595_ (.A(_09567_),
    .B(_09569_),
    .C(_09573_),
    .Y(_09576_));
 sky130_fd_sc_hd__inv_2 _19596_ (.A(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__o2bb2ai_2 _19597_ (.A1_N(_09432_),
    .A2_N(_09425_),
    .B1(_09423_),
    .B2(_09427_),
    .Y(_09578_));
 sky130_fd_sc_hd__o21ai_2 _19598_ (.A1(_01945_),
    .A2(_02207_),
    .B1(_09420_),
    .Y(_09580_));
 sky130_fd_sc_hd__a31o_1 _19599_ (.A1(_09418_),
    .A2(net54),
    .A3(net4),
    .B1(_09419_),
    .X(_09581_));
 sky130_fd_sc_hd__and2_1 _19600_ (.A(net5),
    .B(net54),
    .X(_09582_));
 sky130_fd_sc_hd__nand2_1 _19601_ (.A(net7),
    .B(net53),
    .Y(_09583_));
 sky130_fd_sc_hd__nand4_1 _19602_ (.A(net6),
    .B(net7),
    .C(net52),
    .D(net53),
    .Y(_09584_));
 sky130_fd_sc_hd__a22o_1 _19603_ (.A1(net7),
    .A2(net52),
    .B1(net53),
    .B2(net6),
    .X(_09585_));
 sky130_fd_sc_hd__o211a_2 _19604_ (.A1(_09417_),
    .A2(_09583_),
    .B1(_09582_),
    .C1(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__o2111ai_2 _19605_ (.A1(_09417_),
    .A2(_09583_),
    .B1(net5),
    .C1(net54),
    .D1(_09585_),
    .Y(_09587_));
 sky130_fd_sc_hd__a21oi_1 _19606_ (.A1(_09584_),
    .A2(_09585_),
    .B1(_09582_),
    .Y(_09588_));
 sky130_fd_sc_hd__a22o_1 _19607_ (.A1(net5),
    .A2(net54),
    .B1(_09584_),
    .B2(_09585_),
    .X(_09589_));
 sky130_fd_sc_hd__nand2_2 _19608_ (.A(_09581_),
    .B(_09589_),
    .Y(_09591_));
 sky130_fd_sc_hd__nand3_1 _19609_ (.A(_09589_),
    .B(_09581_),
    .C(_09587_),
    .Y(_09592_));
 sky130_fd_sc_hd__o2bb2ai_4 _19610_ (.A1_N(_09418_),
    .A2_N(_09580_),
    .B1(_09586_),
    .B2(_09588_),
    .Y(_09593_));
 sky130_fd_sc_hd__nand2_1 _19611_ (.A(net4),
    .B(net56),
    .Y(_09594_));
 sky130_fd_sc_hd__nand2_1 _19612_ (.A(_01923_),
    .B(net57),
    .Y(_09595_));
 sky130_fd_sc_hd__and4_1 _19613_ (.A(_01923_),
    .B(net4),
    .C(net56),
    .D(net57),
    .X(_09596_));
 sky130_fd_sc_hd__o22a_1 _19614_ (.A1(net3),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01945_),
    .X(_09597_));
 sky130_fd_sc_hd__and3_1 _19615_ (.A(_01923_),
    .B(_09594_),
    .C(net57),
    .X(_09598_));
 sky130_fd_sc_hd__and3_1 _19616_ (.A(_09595_),
    .B(net56),
    .C(net4),
    .X(_09599_));
 sky130_fd_sc_hd__nor2_1 _19617_ (.A(_09596_),
    .B(_09597_),
    .Y(_09600_));
 sky130_fd_sc_hd__o211a_1 _19618_ (.A1(_09598_),
    .A2(_09599_),
    .B1(_09592_),
    .C1(_09593_),
    .X(_09602_));
 sky130_fd_sc_hd__o221ai_4 _19619_ (.A1(_09598_),
    .A2(_09599_),
    .B1(_09586_),
    .B2(_09591_),
    .C1(_09593_),
    .Y(_09603_));
 sky130_fd_sc_hd__a21oi_1 _19620_ (.A1(_09592_),
    .A2(_09593_),
    .B1(_09600_),
    .Y(_09604_));
 sky130_fd_sc_hd__o2bb2ai_2 _19621_ (.A1_N(_09592_),
    .A2_N(_09593_),
    .B1(_09596_),
    .B2(_09597_),
    .Y(_09605_));
 sky130_fd_sc_hd__nand2_1 _19622_ (.A(_09578_),
    .B(_09605_),
    .Y(_09606_));
 sky130_fd_sc_hd__nand3_4 _19623_ (.A(_09578_),
    .B(_09603_),
    .C(_09605_),
    .Y(_09607_));
 sky130_fd_sc_hd__inv_2 _19624_ (.A(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__o21bai_2 _19625_ (.A1(_09602_),
    .A2(_09604_),
    .B1_N(_09578_),
    .Y(_09609_));
 sky130_fd_sc_hd__or4b_1 _19626_ (.A(net2),
    .B(_02240_),
    .C(_09429_),
    .D_N(_09609_),
    .X(_09610_));
 sky130_fd_sc_hd__inv_2 _19627_ (.A(_09610_),
    .Y(_09611_));
 sky130_fd_sc_hd__o211a_1 _19628_ (.A1(_09602_),
    .A2(_09606_),
    .B1(_09430_),
    .C1(_09609_),
    .X(_09613_));
 sky130_fd_sc_hd__a21oi_2 _19629_ (.A1(_09607_),
    .A2(_09609_),
    .B1(_09430_),
    .Y(_09614_));
 sky130_fd_sc_hd__o311a_2 _19630_ (.A1(net2),
    .A2(_02240_),
    .A3(_09429_),
    .B1(_09607_),
    .C1(_09609_),
    .X(_09615_));
 sky130_fd_sc_hd__a21boi_2 _19631_ (.A1(_09607_),
    .A2(_09609_),
    .B1_N(_09430_),
    .Y(_09616_));
 sky130_fd_sc_hd__nor2_1 _19632_ (.A(_09615_),
    .B(_09616_),
    .Y(_09617_));
 sky130_fd_sc_hd__o2bb2ai_1 _19633_ (.A1_N(_09575_),
    .A2_N(_09576_),
    .B1(_09613_),
    .B2(_09614_),
    .Y(_09618_));
 sky130_fd_sc_hd__o211ai_2 _19634_ (.A1(_09615_),
    .A2(_09616_),
    .B1(_09575_),
    .C1(_09576_),
    .Y(_09619_));
 sky130_fd_sc_hd__o2bb2ai_2 _19635_ (.A1_N(_09575_),
    .A2_N(_09576_),
    .B1(_09615_),
    .B2(_09616_),
    .Y(_09620_));
 sky130_fd_sc_hd__o211ai_4 _19636_ (.A1(_09613_),
    .A2(_09614_),
    .B1(_09575_),
    .C1(_09576_),
    .Y(_09621_));
 sky130_fd_sc_hd__a22oi_4 _19637_ (.A1(_09329_),
    .A2(_09334_),
    .B1(_09620_),
    .B2(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__nand3_2 _19638_ (.A(_09536_),
    .B(_09618_),
    .C(_09619_),
    .Y(_09624_));
 sky130_fd_sc_hd__a21oi_1 _19639_ (.A1(_09618_),
    .A2(_09619_),
    .B1(_09536_),
    .Y(_09625_));
 sky130_fd_sc_hd__nand3_4 _19640_ (.A(_09534_),
    .B(_09620_),
    .C(_09621_),
    .Y(_09626_));
 sky130_fd_sc_hd__o21ai_4 _19641_ (.A1(_09479_),
    .A2(_09483_),
    .B1(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__o211a_2 _19642_ (.A1(_09479_),
    .A2(_09483_),
    .B1(_09624_),
    .C1(_09626_),
    .X(_09628_));
 sky130_fd_sc_hd__o211ai_4 _19643_ (.A1(_09479_),
    .A2(_09483_),
    .B1(_09624_),
    .C1(_09626_),
    .Y(_09629_));
 sky130_fd_sc_hd__a22oi_4 _19644_ (.A1(_09478_),
    .A2(_09533_),
    .B1(_09624_),
    .B2(_09626_),
    .Y(_09630_));
 sky130_fd_sc_hd__o2bb2ai_4 _19645_ (.A1_N(_09478_),
    .A2_N(_09533_),
    .B1(_09622_),
    .B2(_09625_),
    .Y(_09631_));
 sky130_fd_sc_hd__o21ai_4 _19646_ (.A1(_09379_),
    .A2(_09391_),
    .B1(_09386_),
    .Y(_09632_));
 sky130_fd_sc_hd__nand2_1 _19647_ (.A(net38),
    .B(net21),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2_2 _19648_ (.A(net36),
    .B(net24),
    .Y(_09635_));
 sky130_fd_sc_hd__a22oi_2 _19649_ (.A1(net37),
    .A2(net22),
    .B1(net24),
    .B2(net36),
    .Y(_09636_));
 sky130_fd_sc_hd__a22o_1 _19650_ (.A1(net37),
    .A2(net22),
    .B1(net24),
    .B2(net36),
    .X(_09637_));
 sky130_fd_sc_hd__nand3_1 _19651_ (.A(net36),
    .B(net37),
    .C(net22),
    .Y(_09638_));
 sky130_fd_sc_hd__and4_2 _19652_ (.A(net36),
    .B(net37),
    .C(net22),
    .D(net24),
    .X(_09639_));
 sky130_fd_sc_hd__o211a_2 _19653_ (.A1(_02218_),
    .A2(_09638_),
    .B1(_09637_),
    .C1(_09633_),
    .X(_09640_));
 sky130_fd_sc_hd__o21ba_2 _19654_ (.A1(_09636_),
    .A2(_09639_),
    .B1_N(_09633_),
    .X(_09641_));
 sky130_fd_sc_hd__o21ai_1 _19655_ (.A1(_09636_),
    .A2(_09639_),
    .B1(_09633_),
    .Y(_09642_));
 sky130_fd_sc_hd__o2111ai_2 _19656_ (.A1(_02218_),
    .A2(_09638_),
    .B1(net38),
    .C1(net21),
    .D1(_09637_),
    .Y(_09643_));
 sky130_fd_sc_hd__nand2_1 _19657_ (.A(_09642_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__o2111ai_4 _19658_ (.A1(net64),
    .A2(net34),
    .B1(net35),
    .C1(net24),
    .D1(net25),
    .Y(_09646_));
 sky130_fd_sc_hd__o21ai_2 _19659_ (.A1(_02251_),
    .A2(_08978_),
    .B1(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__o21a_1 _19660_ (.A1(_02251_),
    .A2(_08978_),
    .B1(_09646_),
    .X(_09648_));
 sky130_fd_sc_hd__and2_4 _19661_ (.A(net35),
    .B(net25),
    .X(_09649_));
 sky130_fd_sc_hd__o211ai_4 _19662_ (.A1(_01934_),
    .A2(_02251_),
    .B1(_08979_),
    .C1(_09346_),
    .Y(_09650_));
 sky130_fd_sc_hd__nand2_1 _19663_ (.A(_09347_),
    .B(_09649_),
    .Y(_09651_));
 sky130_fd_sc_hd__o21ai_1 _19664_ (.A1(_01934_),
    .A2(_02251_),
    .B1(_09347_),
    .Y(_09652_));
 sky130_fd_sc_hd__and3_1 _19665_ (.A(_08979_),
    .B(_09346_),
    .C(_09649_),
    .X(_09653_));
 sky130_fd_sc_hd__o2111ai_1 _19666_ (.A1(net64),
    .A2(net34),
    .B1(net35),
    .C1(net25),
    .D1(_08979_),
    .Y(_09654_));
 sky130_fd_sc_hd__nand3_1 _19667_ (.A(_09648_),
    .B(_09650_),
    .C(_09651_),
    .Y(_09655_));
 sky130_fd_sc_hd__and4_4 _19668_ (.A(net64),
    .B(net34),
    .C(net35),
    .D(net25),
    .X(_09657_));
 sky130_fd_sc_hd__nand4_4 _19669_ (.A(net64),
    .B(net34),
    .C(net35),
    .D(net25),
    .Y(_09658_));
 sky130_fd_sc_hd__nand3_4 _19670_ (.A(_09651_),
    .B(_09647_),
    .C(_09650_),
    .Y(_09659_));
 sky130_fd_sc_hd__o211ai_2 _19671_ (.A1(_09649_),
    .A2(_09346_),
    .B1(_08979_),
    .C1(_09646_),
    .Y(_09660_));
 sky130_fd_sc_hd__nand3_1 _19672_ (.A(_09648_),
    .B(_09652_),
    .C(_09654_),
    .Y(_09661_));
 sky130_fd_sc_hd__a2bb2oi_4 _19673_ (.A1_N(_09640_),
    .A2_N(_09641_),
    .B1(_09659_),
    .B2(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__o221ai_4 _19674_ (.A1(_01934_),
    .A2(_08979_),
    .B1(_09640_),
    .B2(_09641_),
    .C1(_09655_),
    .Y(_09663_));
 sky130_fd_sc_hd__a32oi_1 _19675_ (.A1(_09651_),
    .A2(_09647_),
    .A3(_09650_),
    .B1(_09643_),
    .B2(_09642_),
    .Y(_09664_));
 sky130_fd_sc_hd__o211a_1 _19676_ (.A1(_09653_),
    .A2(_09660_),
    .B1(_09659_),
    .C1(_09644_),
    .X(_09665_));
 sky130_fd_sc_hd__o211ai_4 _19677_ (.A1(_09660_),
    .A2(_09653_),
    .B1(_09659_),
    .C1(_09644_),
    .Y(_09666_));
 sky130_fd_sc_hd__a21oi_1 _19678_ (.A1(_09661_),
    .A2(_09664_),
    .B1(_09662_),
    .Y(_09668_));
 sky130_fd_sc_hd__a21oi_2 _19679_ (.A1(_09663_),
    .A2(_09666_),
    .B1(_09341_),
    .Y(_09669_));
 sky130_fd_sc_hd__o22ai_4 _19680_ (.A1(_08651_),
    .A2(_09339_),
    .B1(_09662_),
    .B2(_09665_),
    .Y(_09670_));
 sky130_fd_sc_hd__o2111a_1 _19681_ (.A1(_07698_),
    .A2(_08650_),
    .B1(_09340_),
    .C1(_09663_),
    .D1(_09666_),
    .X(_09671_));
 sky130_fd_sc_hd__nand3_4 _19682_ (.A(_09341_),
    .B(_09663_),
    .C(_09666_),
    .Y(_09672_));
 sky130_fd_sc_hd__nand2_1 _19683_ (.A(_09670_),
    .B(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__o21a_1 _19684_ (.A1(_09353_),
    .A2(_09369_),
    .B1(_09355_),
    .X(_09674_));
 sky130_fd_sc_hd__o21ai_2 _19685_ (.A1(_09353_),
    .A2(_09369_),
    .B1(_09355_),
    .Y(_09675_));
 sky130_fd_sc_hd__a21oi_2 _19686_ (.A1(_09670_),
    .A2(_09672_),
    .B1(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__o21ai_2 _19687_ (.A1(_09669_),
    .A2(_09671_),
    .B1(_09674_),
    .Y(_09677_));
 sky130_fd_sc_hd__and3_1 _19688_ (.A(_09670_),
    .B(_09672_),
    .C(_09675_),
    .X(_09679_));
 sky130_fd_sc_hd__nand3_2 _19689_ (.A(_09670_),
    .B(_09672_),
    .C(_09675_),
    .Y(_09680_));
 sky130_fd_sc_hd__a22oi_1 _19690_ (.A1(_09384_),
    .A2(_09386_),
    .B1(_09677_),
    .B2(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__o22ai_4 _19691_ (.A1(_09383_),
    .A2(_09385_),
    .B1(_09676_),
    .B2(_09679_),
    .Y(_09682_));
 sky130_fd_sc_hd__o41ai_2 _19692_ (.A1(_06880_),
    .A2(_07129_),
    .A3(_07680_),
    .A4(_08959_),
    .B1(_09680_),
    .Y(_09683_));
 sky130_fd_sc_hd__a21oi_1 _19693_ (.A1(_09673_),
    .A2(_09674_),
    .B1(_09388_),
    .Y(_09684_));
 sky130_fd_sc_hd__nand4_4 _19694_ (.A(_09384_),
    .B(_09386_),
    .C(_09677_),
    .D(_09680_),
    .Y(_09685_));
 sky130_fd_sc_hd__a21oi_1 _19695_ (.A1(_09680_),
    .A2(_09684_),
    .B1(_09681_),
    .Y(_09686_));
 sky130_fd_sc_hd__a21oi_4 _19696_ (.A1(_09682_),
    .A2(_09685_),
    .B1(_09632_),
    .Y(_09687_));
 sky130_fd_sc_hd__a21o_2 _19697_ (.A1(_09682_),
    .A2(_09685_),
    .B1(_09632_),
    .X(_09688_));
 sky130_fd_sc_hd__o311a_4 _19698_ (.A1(_09385_),
    .A2(_09676_),
    .A3(_09683_),
    .B1(_09682_),
    .C1(_09632_),
    .X(_09690_));
 sky130_fd_sc_hd__nand3_2 _19699_ (.A(_09632_),
    .B(_09682_),
    .C(_09685_),
    .Y(_09691_));
 sky130_fd_sc_hd__a21boi_4 _19700_ (.A1(_09376_),
    .A2(_09378_),
    .B1_N(_09377_),
    .Y(_09692_));
 sky130_fd_sc_hd__o21ai_2 _19701_ (.A1(_09342_),
    .A2(_09375_),
    .B1(_09381_),
    .Y(_09693_));
 sky130_fd_sc_hd__a21oi_2 _19702_ (.A1(_09312_),
    .A2(_09291_),
    .B1(_09309_),
    .Y(_09694_));
 sky130_fd_sc_hd__o21ai_2 _19703_ (.A1(_09356_),
    .A2(_09361_),
    .B1(_09359_),
    .Y(_09695_));
 sky130_fd_sc_hd__o21a_1 _19704_ (.A1(_09356_),
    .A2(_09361_),
    .B1(_09359_),
    .X(_09696_));
 sky130_fd_sc_hd__nand2_4 _19705_ (.A(net39),
    .B(net20),
    .Y(_09697_));
 sky130_fd_sc_hd__a22oi_2 _19706_ (.A1(net40),
    .A2(net19),
    .B1(net20),
    .B2(net39),
    .Y(_09698_));
 sky130_fd_sc_hd__a22o_2 _19707_ (.A1(net40),
    .A2(net19),
    .B1(net20),
    .B2(net39),
    .X(_09699_));
 sky130_fd_sc_hd__nand2_4 _19708_ (.A(net40),
    .B(net20),
    .Y(_09701_));
 sky130_fd_sc_hd__and4_2 _19709_ (.A(net39),
    .B(net40),
    .C(net19),
    .D(net20),
    .X(_09702_));
 sky130_fd_sc_hd__o2bb2ai_2 _19710_ (.A1_N(_09301_),
    .A2_N(_09697_),
    .B1(_09701_),
    .B2(_09298_),
    .Y(_09703_));
 sky130_fd_sc_hd__o221ai_4 _19711_ (.A1(_02010_),
    .A2(_02131_),
    .B1(_09298_),
    .B2(_09701_),
    .C1(_09699_),
    .Y(_09704_));
 sky130_fd_sc_hd__nand3_2 _19712_ (.A(_09703_),
    .B(net18),
    .C(net41),
    .Y(_09705_));
 sky130_fd_sc_hd__o21ai_2 _19713_ (.A1(_02010_),
    .A2(_02131_),
    .B1(_09703_),
    .Y(_09706_));
 sky130_fd_sc_hd__o2111ai_4 _19714_ (.A1(_09298_),
    .A2(_09701_),
    .B1(net41),
    .C1(net18),
    .D1(_09699_),
    .Y(_09707_));
 sky130_fd_sc_hd__and3_1 _19715_ (.A(_09696_),
    .B(_09704_),
    .C(_09705_),
    .X(_09708_));
 sky130_fd_sc_hd__nand3_2 _19716_ (.A(_09696_),
    .B(_09704_),
    .C(_09705_),
    .Y(_09709_));
 sky130_fd_sc_hd__and3_1 _19717_ (.A(_09706_),
    .B(_09707_),
    .C(_09695_),
    .X(_09710_));
 sky130_fd_sc_hd__nand3_4 _19718_ (.A(_09706_),
    .B(_09707_),
    .C(_09695_),
    .Y(_09712_));
 sky130_fd_sc_hd__a31o_1 _19719_ (.A1(_09300_),
    .A2(net17),
    .A3(net41),
    .B1(_09302_),
    .X(_09713_));
 sky130_fd_sc_hd__o21a_1 _19720_ (.A1(_09297_),
    .A2(_09299_),
    .B1(_09303_),
    .X(_09714_));
 sky130_fd_sc_hd__a21oi_1 _19721_ (.A1(_09709_),
    .A2(_09712_),
    .B1(_09713_),
    .Y(_09715_));
 sky130_fd_sc_hd__a21o_1 _19722_ (.A1(_09709_),
    .A2(_09712_),
    .B1(_09713_),
    .X(_09716_));
 sky130_fd_sc_hd__a31oi_4 _19723_ (.A1(_09696_),
    .A2(_09704_),
    .A3(_09705_),
    .B1(_09714_),
    .Y(_09717_));
 sky130_fd_sc_hd__and3_1 _19724_ (.A(_09709_),
    .B(_09712_),
    .C(_09713_),
    .X(_09718_));
 sky130_fd_sc_hd__nand2_1 _19725_ (.A(_09717_),
    .B(_09712_),
    .Y(_09719_));
 sky130_fd_sc_hd__a21o_1 _19726_ (.A1(_09709_),
    .A2(_09712_),
    .B1(_09714_),
    .X(_09720_));
 sky130_fd_sc_hd__o2111ai_4 _19727_ (.A1(_09297_),
    .A2(_09299_),
    .B1(_09303_),
    .C1(_09709_),
    .D1(_09712_),
    .Y(_09721_));
 sky130_fd_sc_hd__o221a_2 _19728_ (.A1(_09292_),
    .A2(_09311_),
    .B1(_09715_),
    .B2(_09718_),
    .C1(_09310_),
    .X(_09723_));
 sky130_fd_sc_hd__nand3_4 _19729_ (.A(_09720_),
    .B(_09721_),
    .C(_09694_),
    .Y(_09724_));
 sky130_fd_sc_hd__o211a_1 _19730_ (.A1(_09309_),
    .A2(_09313_),
    .B1(_09716_),
    .C1(_09719_),
    .X(_09725_));
 sky130_fd_sc_hd__o211ai_4 _19731_ (.A1(_09309_),
    .A2(_09313_),
    .B1(_09716_),
    .C1(_09719_),
    .Y(_09726_));
 sky130_fd_sc_hd__o22a_2 _19732_ (.A1(_02054_),
    .A2(_02065_),
    .B1(_09057_),
    .B2(_09254_),
    .X(_09727_));
 sky130_fd_sc_hd__o21ai_2 _19733_ (.A1(_02054_),
    .A2(_02065_),
    .B1(_09255_),
    .Y(_09728_));
 sky130_fd_sc_hd__nand2_1 _19734_ (.A(net42),
    .B(net17),
    .Y(_09729_));
 sky130_fd_sc_hd__a22oi_1 _19735_ (.A1(net43),
    .A2(net16),
    .B1(net17),
    .B2(net42),
    .Y(_09730_));
 sky130_fd_sc_hd__a22o_1 _19736_ (.A1(net43),
    .A2(net16),
    .B1(net17),
    .B2(net42),
    .X(_09731_));
 sky130_fd_sc_hd__nand4_4 _19737_ (.A(net42),
    .B(net43),
    .C(net16),
    .D(net17),
    .Y(_09732_));
 sky130_fd_sc_hd__nand2_1 _19738_ (.A(net45),
    .B(net15),
    .Y(_09734_));
 sky130_fd_sc_hd__a22oi_2 _19739_ (.A1(net45),
    .A2(net15),
    .B1(_09731_),
    .B2(_09732_),
    .Y(_09735_));
 sky130_fd_sc_hd__a22o_1 _19740_ (.A1(net45),
    .A2(net15),
    .B1(_09731_),
    .B2(_09732_),
    .X(_09736_));
 sky130_fd_sc_hd__and4_1 _19741_ (.A(_09731_),
    .B(_09732_),
    .C(net45),
    .D(net15),
    .X(_09737_));
 sky130_fd_sc_hd__nand4_4 _19742_ (.A(_09731_),
    .B(_09732_),
    .C(net45),
    .D(net15),
    .Y(_09738_));
 sky130_fd_sc_hd__nand2_1 _19743_ (.A(_09736_),
    .B(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__a22oi_2 _19744_ (.A1(_09257_),
    .A2(_09728_),
    .B1(_09736_),
    .B2(_09738_),
    .Y(_09740_));
 sky130_fd_sc_hd__o22ai_4 _19745_ (.A1(_09256_),
    .A2(_09727_),
    .B1(_09735_),
    .B2(_09737_),
    .Y(_09741_));
 sky130_fd_sc_hd__and4_2 _19746_ (.A(_09257_),
    .B(_09728_),
    .C(_09736_),
    .D(_09738_),
    .X(_09742_));
 sky130_fd_sc_hd__nand4_4 _19747_ (.A(_09257_),
    .B(_09728_),
    .C(_09736_),
    .D(_09738_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand2_2 _19748_ (.A(net11),
    .B(net48),
    .Y(_09745_));
 sky130_fd_sc_hd__and4_1 _19749_ (.A(net13),
    .B(net14),
    .C(net46),
    .D(net47),
    .X(_09746_));
 sky130_fd_sc_hd__nand4_2 _19750_ (.A(net13),
    .B(net14),
    .C(net46),
    .D(net47),
    .Y(_09747_));
 sky130_fd_sc_hd__a22oi_4 _19751_ (.A1(net14),
    .A2(net46),
    .B1(net47),
    .B2(net13),
    .Y(_09748_));
 sky130_fd_sc_hd__a22o_1 _19752_ (.A1(net14),
    .A2(net46),
    .B1(net47),
    .B2(net13),
    .X(_09749_));
 sky130_fd_sc_hd__o311a_1 _19753_ (.A1(_02065_),
    .A2(_02087_),
    .A3(_09267_),
    .B1(_09745_),
    .C1(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__a211o_1 _19754_ (.A1(net11),
    .A2(net48),
    .B1(_09746_),
    .C1(_09748_),
    .X(_09751_));
 sky130_fd_sc_hd__a21oi_2 _19755_ (.A1(_09747_),
    .A2(_09749_),
    .B1(_09745_),
    .Y(_09752_));
 sky130_fd_sc_hd__a211o_1 _19756_ (.A1(_09747_),
    .A2(_09749_),
    .B1(_02032_),
    .C1(_02109_),
    .X(_09753_));
 sky130_fd_sc_hd__nor2_1 _19757_ (.A(_09750_),
    .B(_09752_),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_1 _19758_ (.A(_09751_),
    .B(_09753_),
    .Y(_09756_));
 sky130_fd_sc_hd__and3_1 _19759_ (.A(_09754_),
    .B(_09743_),
    .C(_09741_),
    .X(_09757_));
 sky130_fd_sc_hd__o2bb2a_1 _19760_ (.A1_N(_09741_),
    .A2_N(_09743_),
    .B1(_09750_),
    .B2(_09752_),
    .X(_09758_));
 sky130_fd_sc_hd__a21oi_2 _19761_ (.A1(_09741_),
    .A2(_09743_),
    .B1(_09756_),
    .Y(_09759_));
 sky130_fd_sc_hd__a21o_1 _19762_ (.A1(_09741_),
    .A2(_09743_),
    .B1(_09756_),
    .X(_09760_));
 sky130_fd_sc_hd__o21ai_4 _19763_ (.A1(_09750_),
    .A2(_09752_),
    .B1(_09741_),
    .Y(_09761_));
 sky130_fd_sc_hd__o311a_1 _19764_ (.A1(_09256_),
    .A2(_09727_),
    .A3(_09739_),
    .B1(_09741_),
    .C1(_09756_),
    .X(_09762_));
 sky130_fd_sc_hd__o21ai_2 _19765_ (.A1(_09742_),
    .A2(_09761_),
    .B1(_09760_),
    .Y(_09763_));
 sky130_fd_sc_hd__o2bb2ai_4 _19766_ (.A1_N(_09724_),
    .A2_N(_09726_),
    .B1(_09757_),
    .B2(_09758_),
    .Y(_09764_));
 sky130_fd_sc_hd__o32a_2 _19767_ (.A1(_09694_),
    .A2(_09715_),
    .A3(_09718_),
    .B1(_09759_),
    .B2(_09762_),
    .X(_09765_));
 sky130_fd_sc_hd__o211ai_4 _19768_ (.A1(_09759_),
    .A2(_09762_),
    .B1(_09724_),
    .C1(_09726_),
    .Y(_09767_));
 sky130_fd_sc_hd__o2bb2ai_1 _19769_ (.A1_N(_09724_),
    .A2_N(_09726_),
    .B1(_09759_),
    .B2(_09762_),
    .Y(_09768_));
 sky130_fd_sc_hd__o2111ai_4 _19770_ (.A1(_09742_),
    .A2(_09761_),
    .B1(_09760_),
    .C1(_09724_),
    .D1(_09726_),
    .Y(_09769_));
 sky130_fd_sc_hd__nand3_4 _19771_ (.A(_09764_),
    .B(_09767_),
    .C(_09692_),
    .Y(_09770_));
 sky130_fd_sc_hd__a21oi_4 _19772_ (.A1(_09764_),
    .A2(_09767_),
    .B1(_09692_),
    .Y(_09771_));
 sky130_fd_sc_hd__nand3_4 _19773_ (.A(_09693_),
    .B(_09768_),
    .C(_09769_),
    .Y(_09772_));
 sky130_fd_sc_hd__and3_1 _19774_ (.A(_09280_),
    .B(_09282_),
    .C(_09320_),
    .X(_09773_));
 sky130_fd_sc_hd__a31o_1 _19775_ (.A1(_09280_),
    .A2(_09282_),
    .A3(_09320_),
    .B1(_09321_),
    .X(_09774_));
 sky130_fd_sc_hd__o21a_1 _19776_ (.A1(_09319_),
    .A2(_09323_),
    .B1(_09770_),
    .X(_09775_));
 sky130_fd_sc_hd__o21ai_4 _19777_ (.A1(_09319_),
    .A2(_09323_),
    .B1(_09770_),
    .Y(_09776_));
 sky130_fd_sc_hd__o211ai_2 _19778_ (.A1(_09319_),
    .A2(_09323_),
    .B1(_09770_),
    .C1(_09772_),
    .Y(_09778_));
 sky130_fd_sc_hd__o2bb2ai_4 _19779_ (.A1_N(_09770_),
    .A2_N(_09772_),
    .B1(_09773_),
    .B2(_09321_),
    .Y(_09779_));
 sky130_fd_sc_hd__and3_1 _19780_ (.A(_09770_),
    .B(_09772_),
    .C(_09774_),
    .X(_09780_));
 sky130_fd_sc_hd__a21oi_2 _19781_ (.A1(_09770_),
    .A2(_09772_),
    .B1(_09774_),
    .Y(_09781_));
 sky130_fd_sc_hd__o21a_1 _19782_ (.A1(_09771_),
    .A2(_09776_),
    .B1(_09779_),
    .X(_09782_));
 sky130_fd_sc_hd__o21ai_2 _19783_ (.A1(_09771_),
    .A2(_09776_),
    .B1(_09779_),
    .Y(_09783_));
 sky130_fd_sc_hd__nand3_2 _19784_ (.A(_09688_),
    .B(_09691_),
    .C(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__o22ai_4 _19785_ (.A1(_09687_),
    .A2(_09690_),
    .B1(_09780_),
    .B2(_09781_),
    .Y(_09785_));
 sky130_fd_sc_hd__o21ai_4 _19786_ (.A1(_09687_),
    .A2(_09690_),
    .B1(_09783_),
    .Y(_09786_));
 sky130_fd_sc_hd__o2111ai_4 _19787_ (.A1(_09771_),
    .A2(_09776_),
    .B1(_09779_),
    .C1(_09691_),
    .D1(_09688_),
    .Y(_09787_));
 sky130_fd_sc_hd__nand2_2 _19788_ (.A(_09786_),
    .B(_09787_),
    .Y(_09789_));
 sky130_fd_sc_hd__a2bb2oi_4 _19789_ (.A1_N(_09398_),
    .A2_N(_09403_),
    .B1(_09786_),
    .B2(_09787_),
    .Y(_09790_));
 sky130_fd_sc_hd__o211ai_4 _19790_ (.A1(_09398_),
    .A2(_09403_),
    .B1(_09784_),
    .C1(_09785_),
    .Y(_09791_));
 sky130_fd_sc_hd__a21oi_4 _19791_ (.A1(_09784_),
    .A2(_09785_),
    .B1(_09406_),
    .Y(_09792_));
 sky130_fd_sc_hd__nand4_4 _19792_ (.A(_09399_),
    .B(_09405_),
    .C(_09786_),
    .D(_09787_),
    .Y(_09793_));
 sky130_fd_sc_hd__o221ai_4 _19793_ (.A1(_09622_),
    .A2(_09627_),
    .B1(_09406_),
    .B2(_09789_),
    .C1(_09631_),
    .Y(_09794_));
 sky130_fd_sc_hd__o2111a_1 _19794_ (.A1(_09622_),
    .A2(_09627_),
    .B1(_09631_),
    .C1(_09791_),
    .D1(_09793_),
    .X(_09795_));
 sky130_fd_sc_hd__o2111ai_4 _19795_ (.A1(_09622_),
    .A2(_09627_),
    .B1(_09631_),
    .C1(_09791_),
    .D1(_09793_),
    .Y(_09796_));
 sky130_fd_sc_hd__a22oi_4 _19796_ (.A1(_09629_),
    .A2(_09631_),
    .B1(_09791_),
    .B2(_09793_),
    .Y(_09797_));
 sky130_fd_sc_hd__o22ai_4 _19797_ (.A1(_09628_),
    .A2(_09630_),
    .B1(_09790_),
    .B2(_09792_),
    .Y(_09798_));
 sky130_fd_sc_hd__a22oi_4 _19798_ (.A1(_09409_),
    .A2(_09532_),
    .B1(_09796_),
    .B2(_09798_),
    .Y(_09800_));
 sky130_fd_sc_hd__o2bb2ai_4 _19799_ (.A1_N(_09409_),
    .A2_N(_09532_),
    .B1(_09795_),
    .B2(_09797_),
    .Y(_09801_));
 sky130_fd_sc_hd__o211ai_4 _19800_ (.A1(_09790_),
    .A2(_09794_),
    .B1(_09409_),
    .C1(_09532_),
    .Y(_09802_));
 sky130_fd_sc_hd__o2111a_1 _19801_ (.A1(_09790_),
    .A2(_09794_),
    .B1(_09798_),
    .C1(_09532_),
    .D1(_09409_),
    .X(_09803_));
 sky130_fd_sc_hd__o2111ai_4 _19802_ (.A1(_09790_),
    .A2(_09794_),
    .B1(_09798_),
    .C1(_09532_),
    .D1(_09409_),
    .Y(_09804_));
 sky130_fd_sc_hd__o21ai_1 _19803_ (.A1(_09797_),
    .A2(_09802_),
    .B1(_09801_),
    .Y(_09805_));
 sky130_fd_sc_hd__o211a_1 _19804_ (.A1(_09182_),
    .A2(_09139_),
    .B1(_09181_),
    .C1(_09487_),
    .X(_09806_));
 sky130_fd_sc_hd__or2_2 _19805_ (.A(_09489_),
    .B(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__inv_2 _19806_ (.A(_09807_),
    .Y(_09808_));
 sky130_fd_sc_hd__o2bb2ai_1 _19807_ (.A1_N(_09801_),
    .A2_N(_09804_),
    .B1(_09806_),
    .B2(_09489_),
    .Y(_09809_));
 sky130_fd_sc_hd__o211ai_2 _19808_ (.A1(_09797_),
    .A2(_09802_),
    .B1(_09808_),
    .C1(_09801_),
    .Y(_09811_));
 sky130_fd_sc_hd__o21ai_2 _19809_ (.A1(_09800_),
    .A2(_09803_),
    .B1(_09808_),
    .Y(_09812_));
 sky130_fd_sc_hd__o211ai_4 _19810_ (.A1(_09489_),
    .A2(_09806_),
    .B1(_09804_),
    .C1(_09801_),
    .Y(_09813_));
 sky130_fd_sc_hd__o21ai_1 _19811_ (.A1(_09510_),
    .A2(_09506_),
    .B1(_09505_),
    .Y(_09814_));
 sky130_fd_sc_hd__a21oi_2 _19812_ (.A1(_09507_),
    .A2(_09509_),
    .B1(_09504_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand3_2 _19813_ (.A(_09812_),
    .B(_09813_),
    .C(_09815_),
    .Y(_09816_));
 sky130_fd_sc_hd__a21oi_1 _19814_ (.A1(_09805_),
    .A2(_09807_),
    .B1(_09815_),
    .Y(_09817_));
 sky130_fd_sc_hd__a21oi_2 _19815_ (.A1(_09812_),
    .A2(_09813_),
    .B1(_09815_),
    .Y(_09818_));
 sky130_fd_sc_hd__nand3_1 _19816_ (.A(_09809_),
    .B(_09811_),
    .C(_09814_),
    .Y(_09819_));
 sky130_fd_sc_hd__o31a_1 _19817_ (.A1(_01901_),
    .A2(_02229_),
    .A3(_09128_),
    .B1(_09435_),
    .X(_09820_));
 sky130_fd_sc_hd__a32o_1 _19818_ (.A1(_09413_),
    .A2(_09433_),
    .A3(_09434_),
    .B1(_09438_),
    .B2(_09129_),
    .X(_09822_));
 sky130_fd_sc_hd__inv_2 _19819_ (.A(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__o2bb2ai_1 _19820_ (.A1_N(_09816_),
    .A2_N(_09819_),
    .B1(_09820_),
    .B2(_09436_),
    .Y(_09824_));
 sky130_fd_sc_hd__a31oi_1 _19821_ (.A1(_09812_),
    .A2(_09813_),
    .A3(_09815_),
    .B1(_09823_),
    .Y(_09825_));
 sky130_fd_sc_hd__a31o_1 _19822_ (.A1(_09812_),
    .A2(_09813_),
    .A3(_09815_),
    .B1(_09823_),
    .X(_09826_));
 sky130_fd_sc_hd__a21o_1 _19823_ (.A1(_09816_),
    .A2(_09819_),
    .B1(_09823_),
    .X(_09827_));
 sky130_fd_sc_hd__o211ai_1 _19824_ (.A1(_09436_),
    .A2(_09820_),
    .B1(_09819_),
    .C1(_09816_),
    .Y(_09828_));
 sky130_fd_sc_hd__a21oi_1 _19825_ (.A1(_09516_),
    .A2(_09520_),
    .B1(_09517_),
    .Y(_09829_));
 sky130_fd_sc_hd__nand3_1 _19826_ (.A(_09827_),
    .B(_09828_),
    .C(_09829_),
    .Y(_09830_));
 sky130_fd_sc_hd__o221ai_4 _19827_ (.A1(_09517_),
    .A2(_09523_),
    .B1(_09818_),
    .B2(_09826_),
    .C1(_09824_),
    .Y(_09831_));
 sky130_fd_sc_hd__nand2_1 _19828_ (.A(_09830_),
    .B(_09831_),
    .Y(_09833_));
 sky130_fd_sc_hd__o211ai_2 _19829_ (.A1(_09241_),
    .A2(_09243_),
    .B1(_09530_),
    .C1(_09234_),
    .Y(_09834_));
 sky130_fd_sc_hd__a21oi_1 _19830_ (.A1(_08939_),
    .A2(_09232_),
    .B1(_09529_),
    .Y(_09835_));
 sky130_fd_sc_hd__o21bai_1 _19831_ (.A1(_09233_),
    .A2(_09529_),
    .B1_N(_09528_),
    .Y(_09836_));
 sky130_fd_sc_hd__o21ai_4 _19832_ (.A1(_09528_),
    .A2(_09835_),
    .B1(_09834_),
    .Y(_09837_));
 sky130_fd_sc_hd__xnor2_2 _19833_ (.A(_09833_),
    .B(_09837_),
    .Y(net101));
 sky130_fd_sc_hd__a21bo_1 _19834_ (.A1(_09830_),
    .A2(_09837_),
    .B1_N(_09831_),
    .X(_09838_));
 sky130_fd_sc_hd__o22ai_2 _19835_ (.A1(_09406_),
    .A2(_09789_),
    .B1(_09630_),
    .B2(_09628_),
    .Y(_09839_));
 sky130_fd_sc_hd__a31oi_4 _19836_ (.A1(_09629_),
    .A2(_09631_),
    .A3(_09791_),
    .B1(_09792_),
    .Y(_09840_));
 sky130_fd_sc_hd__o21ai_2 _19837_ (.A1(_09676_),
    .A2(_09683_),
    .B1(_09386_),
    .Y(_09841_));
 sky130_fd_sc_hd__o21ai_1 _19838_ (.A1(_01934_),
    .A2(_08979_),
    .B1(_09663_),
    .Y(_09843_));
 sky130_fd_sc_hd__o31ai_4 _19839_ (.A1(net64),
    .A2(net34),
    .A3(net35),
    .B1(net25),
    .Y(_09844_));
 sky130_fd_sc_hd__o311a_4 _19840_ (.A1(net64),
    .A2(net34),
    .A3(net35),
    .B1(net25),
    .C1(_09658_),
    .X(_09845_));
 sky130_fd_sc_hd__a22oi_4 _19841_ (.A1(net37),
    .A2(net24),
    .B1(net25),
    .B2(net36),
    .Y(_09846_));
 sky130_fd_sc_hd__a22o_1 _19842_ (.A1(net37),
    .A2(net24),
    .B1(net25),
    .B2(net36),
    .X(_09847_));
 sky130_fd_sc_hd__nand2_1 _19843_ (.A(net37),
    .B(net25),
    .Y(_09848_));
 sky130_fd_sc_hd__and4_1 _19844_ (.A(net36),
    .B(net37),
    .C(net24),
    .D(net25),
    .X(_09849_));
 sky130_fd_sc_hd__nand4_1 _19845_ (.A(net36),
    .B(net37),
    .C(net24),
    .D(net25),
    .Y(_09850_));
 sky130_fd_sc_hd__and2_1 _19846_ (.A(net38),
    .B(net22),
    .X(_09851_));
 sky130_fd_sc_hd__a21oi_1 _19847_ (.A1(_09847_),
    .A2(_09850_),
    .B1(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__o21bai_4 _19848_ (.A1(_09846_),
    .A2(_09849_),
    .B1_N(_09851_),
    .Y(_09854_));
 sky130_fd_sc_hd__and3_1 _19849_ (.A(_09847_),
    .B(_09850_),
    .C(_09851_),
    .X(_09855_));
 sky130_fd_sc_hd__o2111ai_4 _19850_ (.A1(_09635_),
    .A2(_09848_),
    .B1(net38),
    .C1(net22),
    .D1(_09847_),
    .Y(_09856_));
 sky130_fd_sc_hd__a21oi_2 _19851_ (.A1(_09854_),
    .A2(_09856_),
    .B1(_09845_),
    .Y(_09857_));
 sky130_fd_sc_hd__o22ai_4 _19852_ (.A1(_09657_),
    .A2(_09844_),
    .B1(_09852_),
    .B2(_09855_),
    .Y(_09858_));
 sky130_fd_sc_hd__and3_2 _19853_ (.A(_09854_),
    .B(_09856_),
    .C(_09845_),
    .X(_09859_));
 sky130_fd_sc_hd__o2111ai_4 _19854_ (.A1(_09346_),
    .A2(_09649_),
    .B1(_09658_),
    .C1(_09854_),
    .D1(_09856_),
    .Y(_09860_));
 sky130_fd_sc_hd__o22ai_4 _19855_ (.A1(_08651_),
    .A2(_09339_),
    .B1(_09857_),
    .B2(_09859_),
    .Y(_09861_));
 sky130_fd_sc_hd__and3_1 _19856_ (.A(_09341_),
    .B(_09858_),
    .C(_09860_),
    .X(_09862_));
 sky130_fd_sc_hd__o2111ai_4 _19857_ (.A1(_07698_),
    .A2(_08650_),
    .B1(_09340_),
    .C1(_09858_),
    .D1(_09860_),
    .Y(_09863_));
 sky130_fd_sc_hd__o211a_1 _19858_ (.A1(_09657_),
    .A2(_09662_),
    .B1(_09861_),
    .C1(_09863_),
    .X(_09865_));
 sky130_fd_sc_hd__o211ai_4 _19859_ (.A1(_09657_),
    .A2(_09662_),
    .B1(_09861_),
    .C1(_09863_),
    .Y(_09866_));
 sky130_fd_sc_hd__a21o_1 _19860_ (.A1(_09861_),
    .A2(_09863_),
    .B1(_09843_),
    .X(_09867_));
 sky130_fd_sc_hd__nand2_1 _19861_ (.A(_09866_),
    .B(_09867_),
    .Y(_09868_));
 sky130_fd_sc_hd__a22oi_2 _19862_ (.A1(_09384_),
    .A2(_09386_),
    .B1(_09866_),
    .B2(_09867_),
    .Y(_09869_));
 sky130_fd_sc_hd__a22o_1 _19863_ (.A1(_09384_),
    .A2(_09386_),
    .B1(_09866_),
    .B2(_09867_),
    .X(_09870_));
 sky130_fd_sc_hd__o311a_2 _19864_ (.A1(_06880_),
    .A2(_07682_),
    .A3(_08959_),
    .B1(_09866_),
    .C1(_09867_),
    .X(_09871_));
 sky130_fd_sc_hd__nand3_1 _19865_ (.A(_09387_),
    .B(_09866_),
    .C(_09867_),
    .Y(_09872_));
 sky130_fd_sc_hd__a21oi_1 _19866_ (.A1(_09871_),
    .A2(_09386_),
    .B1(_09869_),
    .Y(_09873_));
 sky130_fd_sc_hd__o211ai_4 _19867_ (.A1(_09869_),
    .A2(_09871_),
    .B1(_09386_),
    .C1(_09685_),
    .Y(_09874_));
 sky130_fd_sc_hd__inv_2 _19868_ (.A(_09874_),
    .Y(_09876_));
 sky130_fd_sc_hd__and3_1 _19869_ (.A(_09841_),
    .B(_09870_),
    .C(_09872_),
    .X(_09877_));
 sky130_fd_sc_hd__nand3_2 _19870_ (.A(_09841_),
    .B(_09870_),
    .C(_09872_),
    .Y(_09878_));
 sky130_fd_sc_hd__nand2_1 _19871_ (.A(_09874_),
    .B(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__o211a_1 _19872_ (.A1(_09353_),
    .A2(_09369_),
    .B1(_09672_),
    .C1(_09355_),
    .X(_09880_));
 sky130_fd_sc_hd__nand2_1 _19873_ (.A(_09672_),
    .B(_09674_),
    .Y(_09881_));
 sky130_fd_sc_hd__o21ai_2 _19874_ (.A1(_09669_),
    .A2(_09674_),
    .B1(_09672_),
    .Y(_09882_));
 sky130_fd_sc_hd__o21ai_1 _19875_ (.A1(_09341_),
    .A2(_09668_),
    .B1(_09881_),
    .Y(_09883_));
 sky130_fd_sc_hd__o21ai_2 _19876_ (.A1(_09734_),
    .A2(_09730_),
    .B1(_09732_),
    .Y(_09884_));
 sky130_fd_sc_hd__nand2_1 _19877_ (.A(net45),
    .B(net16),
    .Y(_09885_));
 sky130_fd_sc_hd__nand2_1 _19878_ (.A(net43),
    .B(net18),
    .Y(_09887_));
 sky130_fd_sc_hd__nand4_2 _19879_ (.A(net42),
    .B(net43),
    .C(net17),
    .D(net18),
    .Y(_09888_));
 sky130_fd_sc_hd__a22oi_2 _19880_ (.A1(net43),
    .A2(net17),
    .B1(net18),
    .B2(net42),
    .Y(_09889_));
 sky130_fd_sc_hd__a22o_1 _19881_ (.A1(net43),
    .A2(net17),
    .B1(net18),
    .B2(net42),
    .X(_09890_));
 sky130_fd_sc_hd__a2bb2oi_1 _19882_ (.A1_N(_02054_),
    .A2_N(_02098_),
    .B1(_09888_),
    .B2(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__o2bb2ai_1 _19883_ (.A1_N(_09888_),
    .A2_N(_09890_),
    .B1(_02054_),
    .B2(_02098_),
    .Y(_09892_));
 sky130_fd_sc_hd__o2111a_1 _19884_ (.A1(_09729_),
    .A2(_09887_),
    .B1(net45),
    .C1(net16),
    .D1(_09890_),
    .X(_09893_));
 sky130_fd_sc_hd__o2111ai_2 _19885_ (.A1(_09729_),
    .A2(_09887_),
    .B1(net45),
    .C1(net16),
    .D1(_09890_),
    .Y(_09894_));
 sky130_fd_sc_hd__a21oi_1 _19886_ (.A1(_09892_),
    .A2(_09894_),
    .B1(_09884_),
    .Y(_09895_));
 sky130_fd_sc_hd__o21bai_2 _19887_ (.A1(_09891_),
    .A2(_09893_),
    .B1_N(_09884_),
    .Y(_09896_));
 sky130_fd_sc_hd__nand2_1 _19888_ (.A(_09892_),
    .B(_09884_),
    .Y(_09898_));
 sky130_fd_sc_hd__nand3_2 _19889_ (.A(_09892_),
    .B(_09894_),
    .C(_09884_),
    .Y(_09899_));
 sky130_fd_sc_hd__nand2_1 _19890_ (.A(net13),
    .B(net48),
    .Y(_09900_));
 sky130_fd_sc_hd__and4_1 _19891_ (.A(net14),
    .B(net46),
    .C(net15),
    .D(net47),
    .X(_09901_));
 sky130_fd_sc_hd__nand4_2 _19892_ (.A(net14),
    .B(net46),
    .C(net15),
    .D(net47),
    .Y(_09902_));
 sky130_fd_sc_hd__a22oi_1 _19893_ (.A1(net46),
    .A2(net15),
    .B1(net47),
    .B2(net14),
    .Y(_09903_));
 sky130_fd_sc_hd__a22o_1 _19894_ (.A1(net46),
    .A2(net15),
    .B1(net47),
    .B2(net14),
    .X(_09904_));
 sky130_fd_sc_hd__a22o_1 _19895_ (.A1(net13),
    .A2(net48),
    .B1(_09902_),
    .B2(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__nand4_4 _19896_ (.A(_09904_),
    .B(net48),
    .C(net13),
    .D(_09902_),
    .Y(_09906_));
 sky130_fd_sc_hd__nand2_2 _19897_ (.A(_09905_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__and4_2 _19898_ (.A(_09896_),
    .B(_09899_),
    .C(_09905_),
    .D(_09906_),
    .X(_09909_));
 sky130_fd_sc_hd__a22oi_4 _19899_ (.A1(_09896_),
    .A2(_09899_),
    .B1(_09905_),
    .B2(_09906_),
    .Y(_09910_));
 sky130_fd_sc_hd__a21oi_2 _19900_ (.A1(_09896_),
    .A2(_09899_),
    .B1(_09907_),
    .Y(_09911_));
 sky130_fd_sc_hd__and3_2 _19901_ (.A(_09896_),
    .B(_09907_),
    .C(_09899_),
    .X(_09912_));
 sky130_fd_sc_hd__o211a_1 _19902_ (.A1(_09297_),
    .A2(_09299_),
    .B1(_09303_),
    .C1(_09712_),
    .X(_09913_));
 sky130_fd_sc_hd__a21oi_1 _19903_ (.A1(_09709_),
    .A2(_09713_),
    .B1(_09710_),
    .Y(_09914_));
 sky130_fd_sc_hd__o22a_1 _19904_ (.A1(_02010_),
    .A2(_02131_),
    .B1(_09298_),
    .B2(_09701_),
    .X(_09915_));
 sky130_fd_sc_hd__and3_1 _19905_ (.A(_09699_),
    .B(net18),
    .C(net41),
    .X(_09916_));
 sky130_fd_sc_hd__a31o_1 _19906_ (.A1(_09699_),
    .A2(net18),
    .A3(net41),
    .B1(_09702_),
    .X(_09917_));
 sky130_fd_sc_hd__a21oi_2 _19907_ (.A1(_09357_),
    .A2(_09635_),
    .B1(_09633_),
    .Y(_09918_));
 sky130_fd_sc_hd__o22ai_1 _19908_ (.A1(_02218_),
    .A2(_09638_),
    .B1(_09633_),
    .B2(_09636_),
    .Y(_09920_));
 sky130_fd_sc_hd__and2_1 _19909_ (.A(net41),
    .B(net19),
    .X(_09921_));
 sky130_fd_sc_hd__nand2_2 _19910_ (.A(net39),
    .B(net21),
    .Y(_09922_));
 sky130_fd_sc_hd__a22oi_2 _19911_ (.A1(net40),
    .A2(net20),
    .B1(net21),
    .B2(net39),
    .Y(_09923_));
 sky130_fd_sc_hd__a22o_2 _19912_ (.A1(net40),
    .A2(net20),
    .B1(net21),
    .B2(net39),
    .X(_09924_));
 sky130_fd_sc_hd__nand2_4 _19913_ (.A(net40),
    .B(net21),
    .Y(_09925_));
 sky130_fd_sc_hd__o2bb2ai_1 _19914_ (.A1_N(_09701_),
    .A2_N(_09922_),
    .B1(_09925_),
    .B2(_09697_),
    .Y(_09926_));
 sky130_fd_sc_hd__o221ai_4 _19915_ (.A1(_02010_),
    .A2(_02142_),
    .B1(_09697_),
    .B2(_09925_),
    .C1(_09924_),
    .Y(_09927_));
 sky130_fd_sc_hd__nand2_2 _19916_ (.A(_09926_),
    .B(_09921_),
    .Y(_09928_));
 sky130_fd_sc_hd__o2111ai_4 _19917_ (.A1(_09697_),
    .A2(_09925_),
    .B1(net41),
    .C1(net19),
    .D1(_09924_),
    .Y(_09929_));
 sky130_fd_sc_hd__o21ai_2 _19918_ (.A1(_02010_),
    .A2(_02142_),
    .B1(_09926_),
    .Y(_09931_));
 sky130_fd_sc_hd__a2bb2oi_4 _19919_ (.A1_N(_09639_),
    .A2_N(_09918_),
    .B1(_09927_),
    .B2(_09928_),
    .Y(_09932_));
 sky130_fd_sc_hd__o211ai_4 _19920_ (.A1(_09639_),
    .A2(_09918_),
    .B1(_09929_),
    .C1(_09931_),
    .Y(_09933_));
 sky130_fd_sc_hd__a21oi_1 _19921_ (.A1(_09929_),
    .A2(_09931_),
    .B1(_09920_),
    .Y(_09934_));
 sky130_fd_sc_hd__nand3b_4 _19922_ (.A_N(_09920_),
    .B(_09927_),
    .C(_09928_),
    .Y(_09935_));
 sky130_fd_sc_hd__o21a_1 _19923_ (.A1(_09702_),
    .A2(_09916_),
    .B1(_09935_),
    .X(_09936_));
 sky130_fd_sc_hd__o21ai_1 _19924_ (.A1(_09702_),
    .A2(_09916_),
    .B1(_09935_),
    .Y(_09937_));
 sky130_fd_sc_hd__o211a_1 _19925_ (.A1(_09702_),
    .A2(_09916_),
    .B1(_09933_),
    .C1(_09935_),
    .X(_09938_));
 sky130_fd_sc_hd__o211ai_4 _19926_ (.A1(_09702_),
    .A2(_09916_),
    .B1(_09933_),
    .C1(_09935_),
    .Y(_09939_));
 sky130_fd_sc_hd__a21oi_2 _19927_ (.A1(_09933_),
    .A2(_09935_),
    .B1(_09917_),
    .Y(_09940_));
 sky130_fd_sc_hd__o22ai_4 _19928_ (.A1(_09698_),
    .A2(_09915_),
    .B1(_09932_),
    .B2(_09934_),
    .Y(_09942_));
 sky130_fd_sc_hd__o21ai_1 _19929_ (.A1(_09932_),
    .A2(_09937_),
    .B1(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__o211a_1 _19930_ (.A1(_09710_),
    .A2(_09717_),
    .B1(_09939_),
    .C1(_09942_),
    .X(_09944_));
 sky130_fd_sc_hd__o211ai_4 _19931_ (.A1(_09710_),
    .A2(_09717_),
    .B1(_09939_),
    .C1(_09942_),
    .Y(_09945_));
 sky130_fd_sc_hd__o22a_2 _19932_ (.A1(_09708_),
    .A2(_09913_),
    .B1(_09938_),
    .B2(_09940_),
    .X(_09946_));
 sky130_fd_sc_hd__o22ai_4 _19933_ (.A1(_09708_),
    .A2(_09913_),
    .B1(_09938_),
    .B2(_09940_),
    .Y(_09947_));
 sky130_fd_sc_hd__a2bb2oi_1 _19934_ (.A1_N(_09911_),
    .A2_N(_09912_),
    .B1(_09914_),
    .B2(_09943_),
    .Y(_09948_));
 sky130_fd_sc_hd__o211a_1 _19935_ (.A1(_09911_),
    .A2(_09912_),
    .B1(_09945_),
    .C1(_09947_),
    .X(_09949_));
 sky130_fd_sc_hd__o211ai_4 _19936_ (.A1(_09911_),
    .A2(_09912_),
    .B1(_09945_),
    .C1(_09947_),
    .Y(_09950_));
 sky130_fd_sc_hd__a2bb2oi_2 _19937_ (.A1_N(_09909_),
    .A2_N(_09910_),
    .B1(_09945_),
    .B2(_09947_),
    .Y(_09951_));
 sky130_fd_sc_hd__o22ai_4 _19938_ (.A1(_09909_),
    .A2(_09910_),
    .B1(_09944_),
    .B2(_09946_),
    .Y(_09953_));
 sky130_fd_sc_hd__a211oi_2 _19939_ (.A1(_09948_),
    .A2(_09945_),
    .B1(_09883_),
    .C1(_09951_),
    .Y(_09954_));
 sky130_fd_sc_hd__nand3_4 _19940_ (.A(_09882_),
    .B(_09950_),
    .C(_09953_),
    .Y(_09955_));
 sky130_fd_sc_hd__a22oi_4 _19941_ (.A1(_09670_),
    .A2(_09881_),
    .B1(_09950_),
    .B2(_09953_),
    .Y(_09956_));
 sky130_fd_sc_hd__o22ai_4 _19942_ (.A1(_09669_),
    .A2(_09880_),
    .B1(_09949_),
    .B2(_09951_),
    .Y(_09957_));
 sky130_fd_sc_hd__o211a_1 _19943_ (.A1(_09742_),
    .A2(_09761_),
    .B1(_09760_),
    .C1(_09724_),
    .X(_09958_));
 sky130_fd_sc_hd__o21ai_1 _19944_ (.A1(_09723_),
    .A2(_09763_),
    .B1(_09726_),
    .Y(_09959_));
 sky130_fd_sc_hd__a31o_1 _19945_ (.A1(_09694_),
    .A2(_09720_),
    .A3(_09721_),
    .B1(_09765_),
    .X(_09960_));
 sky130_fd_sc_hd__o2bb2ai_1 _19946_ (.A1_N(_09955_),
    .A2_N(_09957_),
    .B1(_09958_),
    .B2(_09725_),
    .Y(_09961_));
 sky130_fd_sc_hd__o2111ai_4 _19947_ (.A1(_09723_),
    .A2(_09763_),
    .B1(_09955_),
    .C1(_09957_),
    .D1(_09726_),
    .Y(_09962_));
 sky130_fd_sc_hd__a2bb2oi_1 _19948_ (.A1_N(_09723_),
    .A2_N(_09765_),
    .B1(_09955_),
    .B2(_09957_),
    .Y(_09964_));
 sky130_fd_sc_hd__o22ai_4 _19949_ (.A1(_09723_),
    .A2(_09765_),
    .B1(_09954_),
    .B2(_09956_),
    .Y(_09965_));
 sky130_fd_sc_hd__o21ai_1 _19950_ (.A1(_09725_),
    .A2(_09958_),
    .B1(_09957_),
    .Y(_09966_));
 sky130_fd_sc_hd__o311a_1 _19951_ (.A1(_09883_),
    .A2(_09949_),
    .A3(_09951_),
    .B1(_09959_),
    .C1(_09957_),
    .X(_09967_));
 sky130_fd_sc_hd__o211ai_4 _19952_ (.A1(_09725_),
    .A2(_09958_),
    .B1(_09957_),
    .C1(_09955_),
    .Y(_09968_));
 sky130_fd_sc_hd__nand2_1 _19953_ (.A(_09961_),
    .B(_09962_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand4_2 _19954_ (.A(_09874_),
    .B(_09878_),
    .C(_09965_),
    .D(_09968_),
    .Y(_09970_));
 sky130_fd_sc_hd__o2bb2ai_2 _19955_ (.A1_N(_09874_),
    .A2_N(_09878_),
    .B1(_09964_),
    .B2(_09967_),
    .Y(_09971_));
 sky130_fd_sc_hd__nand4_2 _19956_ (.A(_09874_),
    .B(_09878_),
    .C(_09961_),
    .D(_09962_),
    .Y(_09972_));
 sky130_fd_sc_hd__nand3_2 _19957_ (.A(_09879_),
    .B(_09965_),
    .C(_09968_),
    .Y(_09973_));
 sky130_fd_sc_hd__a22oi_4 _19958_ (.A1(_09686_),
    .A2(_09632_),
    .B1(_09779_),
    .B2(_09778_),
    .Y(_09975_));
 sky130_fd_sc_hd__o211a_1 _19959_ (.A1(_09687_),
    .A2(_09975_),
    .B1(_09973_),
    .C1(_09972_),
    .X(_09976_));
 sky130_fd_sc_hd__o211ai_4 _19960_ (.A1(_09687_),
    .A2(_09975_),
    .B1(_09973_),
    .C1(_09972_),
    .Y(_09977_));
 sky130_fd_sc_hd__o2111a_1 _19961_ (.A1(_09690_),
    .A2(_09782_),
    .B1(_09970_),
    .C1(_09971_),
    .D1(_09688_),
    .X(_09978_));
 sky130_fd_sc_hd__o2111ai_4 _19962_ (.A1(_09690_),
    .A2(_09782_),
    .B1(_09970_),
    .C1(_09971_),
    .D1(_09688_),
    .Y(_09979_));
 sky130_fd_sc_hd__o32a_1 _19963_ (.A1(_09256_),
    .A2(_09727_),
    .A3(_09739_),
    .B1(_09740_),
    .B2(_09754_),
    .X(_09980_));
 sky130_fd_sc_hd__o32ai_4 _19964_ (.A1(_09256_),
    .A2(_09727_),
    .A3(_09739_),
    .B1(_09740_),
    .B2(_09754_),
    .Y(_09981_));
 sky130_fd_sc_hd__o21ai_2 _19965_ (.A1(_01988_),
    .A2(_02152_),
    .B1(_09549_),
    .Y(_09982_));
 sky130_fd_sc_hd__a31o_1 _19966_ (.A1(_09547_),
    .A2(net51),
    .A3(net8),
    .B1(_09548_),
    .X(_09983_));
 sky130_fd_sc_hd__o31a_1 _19967_ (.A1(_01988_),
    .A2(_02152_),
    .A3(_09545_),
    .B1(_09549_),
    .X(_09984_));
 sky130_fd_sc_hd__a21boi_1 _19968_ (.A1(net11),
    .A2(net48),
    .B1_N(_09747_),
    .Y(_09986_));
 sky130_fd_sc_hd__nor2_1 _19969_ (.A(_09745_),
    .B(_09748_),
    .Y(_09987_));
 sky130_fd_sc_hd__o21ai_1 _19970_ (.A1(_09745_),
    .A2(_09748_),
    .B1(_09747_),
    .Y(_09988_));
 sky130_fd_sc_hd__o21a_1 _19971_ (.A1(_09745_),
    .A2(_09748_),
    .B1(_09747_),
    .X(_09989_));
 sky130_fd_sc_hd__nor2_1 _19972_ (.A(_01999_),
    .B(_02152_),
    .Y(_09990_));
 sky130_fd_sc_hd__a22oi_4 _19973_ (.A1(net11),
    .A2(net49),
    .B1(net50),
    .B2(net10),
    .Y(_09991_));
 sky130_fd_sc_hd__a22o_1 _19974_ (.A1(net11),
    .A2(net49),
    .B1(net50),
    .B2(net10),
    .X(_09992_));
 sky130_fd_sc_hd__and4_1 _19975_ (.A(net10),
    .B(net11),
    .C(net49),
    .D(net50),
    .X(_09993_));
 sky130_fd_sc_hd__nand4_4 _19976_ (.A(net10),
    .B(net11),
    .C(net49),
    .D(net50),
    .Y(_09994_));
 sky130_fd_sc_hd__o211ai_4 _19977_ (.A1(_01999_),
    .A2(_02152_),
    .B1(_09992_),
    .C1(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__o21ai_2 _19978_ (.A1(_09991_),
    .A2(_09993_),
    .B1(_09990_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand4_2 _19979_ (.A(_09992_),
    .B(_09994_),
    .C(net9),
    .D(net51),
    .Y(_09998_));
 sky130_fd_sc_hd__o22ai_4 _19980_ (.A1(_01999_),
    .A2(_02152_),
    .B1(_09991_),
    .B2(_09993_),
    .Y(_09999_));
 sky130_fd_sc_hd__a2bb2oi_4 _19981_ (.A1_N(_09746_),
    .A2_N(_09987_),
    .B1(_09995_),
    .B2(_09997_),
    .Y(_10000_));
 sky130_fd_sc_hd__nand3_4 _19982_ (.A(_09999_),
    .B(_09988_),
    .C(_09998_),
    .Y(_10001_));
 sky130_fd_sc_hd__a2bb2oi_2 _19983_ (.A1_N(_09748_),
    .A2_N(_09986_),
    .B1(_09998_),
    .B2(_09999_),
    .Y(_10002_));
 sky130_fd_sc_hd__nand3_2 _19984_ (.A(_09989_),
    .B(_09995_),
    .C(_09997_),
    .Y(_10003_));
 sky130_fd_sc_hd__nor2_2 _19985_ (.A(_09984_),
    .B(_10002_),
    .Y(_10004_));
 sky130_fd_sc_hd__and3_1 _19986_ (.A(_10003_),
    .B(_09983_),
    .C(_10001_),
    .X(_10005_));
 sky130_fd_sc_hd__nand4_4 _19987_ (.A(_09547_),
    .B(_09982_),
    .C(_10001_),
    .D(_10003_),
    .Y(_10006_));
 sky130_fd_sc_hd__a21oi_2 _19988_ (.A1(_10001_),
    .A2(_10003_),
    .B1(_09983_),
    .Y(_10008_));
 sky130_fd_sc_hd__o2bb2ai_4 _19989_ (.A1_N(_09547_),
    .A2_N(_09982_),
    .B1(_10000_),
    .B2(_10002_),
    .Y(_10009_));
 sky130_fd_sc_hd__a21oi_4 _19990_ (.A1(_10006_),
    .A2(_10009_),
    .B1(_09981_),
    .Y(_10010_));
 sky130_fd_sc_hd__o21ai_2 _19991_ (.A1(_10005_),
    .A2(_10008_),
    .B1(_09980_),
    .Y(_10011_));
 sky130_fd_sc_hd__a221oi_4 _19992_ (.A1(_10004_),
    .A2(_10001_),
    .B1(_09761_),
    .B2(_09743_),
    .C1(_10008_),
    .Y(_10012_));
 sky130_fd_sc_hd__nand3_4 _19993_ (.A(_09981_),
    .B(_10006_),
    .C(_10009_),
    .Y(_10013_));
 sky130_fd_sc_hd__o31a_2 _19994_ (.A1(_09450_),
    .A2(_09540_),
    .A3(_09556_),
    .B1(_09555_),
    .X(_10014_));
 sky130_fd_sc_hd__o21ai_1 _19995_ (.A1(_10010_),
    .A2(_10012_),
    .B1(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__o211ai_2 _19996_ (.A1(_09554_),
    .A2(_09559_),
    .B1(_10011_),
    .C1(_10013_),
    .Y(_10016_));
 sky130_fd_sc_hd__o22ai_4 _19997_ (.A1(_09554_),
    .A2(_09559_),
    .B1(_10010_),
    .B2(_10012_),
    .Y(_10017_));
 sky130_fd_sc_hd__nand4_4 _19998_ (.A(_09555_),
    .B(_09560_),
    .C(_10011_),
    .D(_10013_),
    .Y(_10019_));
 sky130_fd_sc_hd__a21o_1 _19999_ (.A1(_09537_),
    .A2(_09566_),
    .B1(_09564_),
    .X(_10020_));
 sky130_fd_sc_hd__a21oi_4 _20000_ (.A1(_09537_),
    .A2(_09566_),
    .B1(_09564_),
    .Y(_10021_));
 sky130_fd_sc_hd__and3_1 _20001_ (.A(_10017_),
    .B(_10019_),
    .C(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__nand3_2 _20002_ (.A(_10017_),
    .B(_10019_),
    .C(_10021_),
    .Y(_10023_));
 sky130_fd_sc_hd__a21oi_4 _20003_ (.A1(_10017_),
    .A2(_10019_),
    .B1(_10021_),
    .Y(_10024_));
 sky130_fd_sc_hd__nand3_4 _20004_ (.A(_10015_),
    .B(_10020_),
    .C(_10016_),
    .Y(_10025_));
 sky130_fd_sc_hd__a2bb2o_1 _20005_ (.A1_N(_09586_),
    .A2_N(_09591_),
    .B1(_09593_),
    .B2(_09600_),
    .X(_10026_));
 sky130_fd_sc_hd__o2bb2ai_1 _20006_ (.A1_N(_09582_),
    .A2_N(_09585_),
    .B1(_09583_),
    .B2(_09417_),
    .Y(_10027_));
 sky130_fd_sc_hd__nand3_1 _20007_ (.A(net7),
    .B(net8),
    .C(net53),
    .Y(_10028_));
 sky130_fd_sc_hd__and4_1 _20008_ (.A(net7),
    .B(net8),
    .C(net52),
    .D(net53),
    .X(_10030_));
 sky130_fd_sc_hd__nand4_2 _20009_ (.A(net7),
    .B(net8),
    .C(net52),
    .D(net53),
    .Y(_10031_));
 sky130_fd_sc_hd__a22o_1 _20010_ (.A1(net8),
    .A2(net52),
    .B1(net53),
    .B2(net7),
    .X(_10032_));
 sky130_fd_sc_hd__a2bb2oi_1 _20011_ (.A1_N(_01966_),
    .A2_N(_02207_),
    .B1(_10031_),
    .B2(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__o2bb2ai_1 _20012_ (.A1_N(_10031_),
    .A2_N(_10032_),
    .B1(_01966_),
    .B2(_02207_),
    .Y(_10034_));
 sky130_fd_sc_hd__o2111a_1 _20013_ (.A1(_02174_),
    .A2(_10028_),
    .B1(net54),
    .C1(net6),
    .D1(_10032_),
    .X(_10035_));
 sky130_fd_sc_hd__o2111ai_2 _20014_ (.A1(_02174_),
    .A2(_10028_),
    .B1(net54),
    .C1(net6),
    .D1(_10032_),
    .Y(_10036_));
 sky130_fd_sc_hd__o21bai_2 _20015_ (.A1(_10033_),
    .A2(_10035_),
    .B1_N(_10027_),
    .Y(_10037_));
 sky130_fd_sc_hd__a21o_1 _20016_ (.A1(_09584_),
    .A2(_09587_),
    .B1(_10033_),
    .X(_10038_));
 sky130_fd_sc_hd__nand3_1 _20017_ (.A(_10027_),
    .B(_10034_),
    .C(_10036_),
    .Y(_10039_));
 sky130_fd_sc_hd__and4_2 _20018_ (.A(_01945_),
    .B(net5),
    .C(net56),
    .D(net57),
    .X(_10041_));
 sky130_fd_sc_hd__o22a_1 _20019_ (.A1(net4),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01956_),
    .X(_10042_));
 sky130_fd_sc_hd__nor2_2 _20020_ (.A(_10041_),
    .B(_10042_),
    .Y(_10043_));
 sky130_fd_sc_hd__and3_1 _20021_ (.A(_10037_),
    .B(_10039_),
    .C(_10043_),
    .X(_10044_));
 sky130_fd_sc_hd__o211ai_1 _20022_ (.A1(_10035_),
    .A2(_10038_),
    .B1(_10043_),
    .C1(_10037_),
    .Y(_10045_));
 sky130_fd_sc_hd__a21oi_2 _20023_ (.A1(_10037_),
    .A2(_10039_),
    .B1(_10043_),
    .Y(_10046_));
 sky130_fd_sc_hd__a21o_1 _20024_ (.A1(_10037_),
    .A2(_10039_),
    .B1(_10043_),
    .X(_10047_));
 sky130_fd_sc_hd__nand3_2 _20025_ (.A(_10026_),
    .B(_10045_),
    .C(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__o221a_1 _20026_ (.A1(_09591_),
    .A2(_09586_),
    .B1(_10046_),
    .B2(_10044_),
    .C1(_09603_),
    .X(_10049_));
 sky130_fd_sc_hd__o221ai_4 _20027_ (.A1(_09591_),
    .A2(_09586_),
    .B1(_10046_),
    .B2(_10044_),
    .C1(_09603_),
    .Y(_10050_));
 sky130_fd_sc_hd__and3_1 _20028_ (.A(_10050_),
    .B(_09596_),
    .C(_10048_),
    .X(_10052_));
 sky130_fd_sc_hd__o2bb2a_1 _20029_ (.A1_N(_10048_),
    .A2_N(_10050_),
    .B1(_09594_),
    .B2(_09595_),
    .X(_10053_));
 sky130_fd_sc_hd__o311a_1 _20030_ (.A1(_01945_),
    .A2(_02229_),
    .A3(_09595_),
    .B1(_10048_),
    .C1(_10050_),
    .X(_10054_));
 sky130_fd_sc_hd__a21boi_2 _20031_ (.A1(_10048_),
    .A2(_10050_),
    .B1_N(_09596_),
    .Y(_10055_));
 sky130_fd_sc_hd__o21a_1 _20032_ (.A1(_10054_),
    .A2(_10055_),
    .B1(_10023_),
    .X(_10056_));
 sky130_fd_sc_hd__o21ai_2 _20033_ (.A1(_10054_),
    .A2(_10055_),
    .B1(_10023_),
    .Y(_10057_));
 sky130_fd_sc_hd__o2bb2ai_1 _20034_ (.A1_N(_10023_),
    .A2_N(_10025_),
    .B1(_10052_),
    .B2(_10053_),
    .Y(_10058_));
 sky130_fd_sc_hd__o211ai_2 _20035_ (.A1(_10052_),
    .A2(_10053_),
    .B1(_10023_),
    .C1(_10025_),
    .Y(_10059_));
 sky130_fd_sc_hd__o2bb2ai_1 _20036_ (.A1_N(_10023_),
    .A2_N(_10025_),
    .B1(_10054_),
    .B2(_10055_),
    .Y(_10060_));
 sky130_fd_sc_hd__a32o_1 _20037_ (.A1(_09692_),
    .A2(_09764_),
    .A3(_09767_),
    .B1(_09772_),
    .B2(_09774_),
    .X(_10061_));
 sky130_fd_sc_hd__nand3_4 _20038_ (.A(_10059_),
    .B(_10060_),
    .C(_10061_),
    .Y(_10063_));
 sky130_fd_sc_hd__inv_2 _20039_ (.A(_10063_),
    .Y(_10064_));
 sky130_fd_sc_hd__o221ai_4 _20040_ (.A1(_09771_),
    .A2(_09775_),
    .B1(_10024_),
    .B2(_10057_),
    .C1(_10058_),
    .Y(_10065_));
 sky130_fd_sc_hd__o21a_1 _20041_ (.A1(_09613_),
    .A2(_09614_),
    .B1(_09576_),
    .X(_10066_));
 sky130_fd_sc_hd__o21a_1 _20042_ (.A1(_09615_),
    .A2(_09616_),
    .B1(_09575_),
    .X(_10067_));
 sky130_fd_sc_hd__o21a_1 _20043_ (.A1(_09574_),
    .A2(_09617_),
    .B1(_09576_),
    .X(_10068_));
 sky130_fd_sc_hd__a21boi_1 _20044_ (.A1(_10063_),
    .A2(_10065_),
    .B1_N(_10068_),
    .Y(_10069_));
 sky130_fd_sc_hd__o2bb2ai_1 _20045_ (.A1_N(_10063_),
    .A2_N(_10065_),
    .B1(_10066_),
    .B2(_09574_),
    .Y(_10070_));
 sky130_fd_sc_hd__o211a_1 _20046_ (.A1(_09577_),
    .A2(_10067_),
    .B1(_10065_),
    .C1(_10063_),
    .X(_10071_));
 sky130_fd_sc_hd__o211ai_4 _20047_ (.A1(_09577_),
    .A2(_10067_),
    .B1(_10065_),
    .C1(_10063_),
    .Y(_10072_));
 sky130_fd_sc_hd__a21oi_1 _20048_ (.A1(_10063_),
    .A2(_10065_),
    .B1(_10068_),
    .Y(_10074_));
 sky130_fd_sc_hd__o2bb2ai_1 _20049_ (.A1_N(_10063_),
    .A2_N(_10065_),
    .B1(_10067_),
    .B2(_09577_),
    .Y(_10075_));
 sky130_fd_sc_hd__and3_1 _20050_ (.A(_10063_),
    .B(_10065_),
    .C(_10068_),
    .X(_10076_));
 sky130_fd_sc_hd__o2111ai_4 _20051_ (.A1(_09617_),
    .A2(_09574_),
    .B1(_09576_),
    .C1(_10063_),
    .D1(_10065_),
    .Y(_10077_));
 sky130_fd_sc_hd__nand4_1 _20052_ (.A(_09977_),
    .B(_09979_),
    .C(_10070_),
    .D(_10072_),
    .Y(_10078_));
 sky130_fd_sc_hd__o2bb2ai_1 _20053_ (.A1_N(_09977_),
    .A2_N(_09979_),
    .B1(_10069_),
    .B2(_10071_),
    .Y(_10079_));
 sky130_fd_sc_hd__nand4_2 _20054_ (.A(_09977_),
    .B(_09979_),
    .C(_10075_),
    .D(_10077_),
    .Y(_10080_));
 sky130_fd_sc_hd__o2bb2ai_2 _20055_ (.A1_N(_09977_),
    .A2_N(_09979_),
    .B1(_10074_),
    .B2(_10076_),
    .Y(_10081_));
 sky130_fd_sc_hd__a22oi_1 _20056_ (.A1(_09791_),
    .A2(_09839_),
    .B1(_10078_),
    .B2(_10079_),
    .Y(_10082_));
 sky130_fd_sc_hd__nand3_2 _20057_ (.A(_09840_),
    .B(_10080_),
    .C(_10081_),
    .Y(_10083_));
 sky130_fd_sc_hd__a21oi_4 _20058_ (.A1(_10080_),
    .A2(_10081_),
    .B1(_09840_),
    .Y(_10085_));
 sky130_fd_sc_hd__nand4_2 _20059_ (.A(_09791_),
    .B(_09839_),
    .C(_10078_),
    .D(_10079_),
    .Y(_10086_));
 sky130_fd_sc_hd__a31o_1 _20060_ (.A1(_09478_),
    .A2(_09533_),
    .A3(_09626_),
    .B1(_09622_),
    .X(_10087_));
 sky130_fd_sc_hd__a21oi_1 _20061_ (.A1(_10083_),
    .A2(_10086_),
    .B1(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__o21bai_2 _20062_ (.A1(_10082_),
    .A2(_10085_),
    .B1_N(_10087_),
    .Y(_10089_));
 sky130_fd_sc_hd__o21ai_2 _20063_ (.A1(_09622_),
    .A2(_09628_),
    .B1(_10083_),
    .Y(_10090_));
 sky130_fd_sc_hd__and3_1 _20064_ (.A(_10083_),
    .B(_10086_),
    .C(_10087_),
    .X(_10091_));
 sky130_fd_sc_hd__o211ai_2 _20065_ (.A1(_09622_),
    .A2(_09628_),
    .B1(_10083_),
    .C1(_10086_),
    .Y(_10092_));
 sky130_fd_sc_hd__o22ai_4 _20066_ (.A1(_09797_),
    .A2(_09802_),
    .B1(_09807_),
    .B2(_09800_),
    .Y(_10093_));
 sky130_fd_sc_hd__a21oi_1 _20067_ (.A1(_10089_),
    .A2(_10092_),
    .B1(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__o21bai_2 _20068_ (.A1(_10088_),
    .A2(_10091_),
    .B1_N(_10093_),
    .Y(_10095_));
 sky130_fd_sc_hd__o211a_1 _20069_ (.A1(_10085_),
    .A2(_10090_),
    .B1(_10093_),
    .C1(_10089_),
    .X(_10096_));
 sky130_fd_sc_hd__o211ai_4 _20070_ (.A1(_10085_),
    .A2(_10090_),
    .B1(_10093_),
    .C1(_10089_),
    .Y(_10097_));
 sky130_fd_sc_hd__a31o_1 _20071_ (.A1(_09578_),
    .A2(_09603_),
    .A3(_09605_),
    .B1(_09611_),
    .X(_10098_));
 sky130_fd_sc_hd__a21oi_1 _20072_ (.A1(_10095_),
    .A2(_10097_),
    .B1(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__nand3_1 _20073_ (.A(_10095_),
    .B(_10097_),
    .C(_10098_),
    .Y(_10100_));
 sky130_fd_sc_hd__o22ai_2 _20074_ (.A1(_09608_),
    .A2(_09611_),
    .B1(_10094_),
    .B2(_10096_),
    .Y(_10101_));
 sky130_fd_sc_hd__nand3b_1 _20075_ (.A_N(_10098_),
    .B(_10097_),
    .C(_10095_),
    .Y(_10102_));
 sky130_fd_sc_hd__a22oi_2 _20076_ (.A1(_09817_),
    .A2(_09811_),
    .B1(_09816_),
    .B2(_09822_),
    .Y(_10103_));
 sky130_fd_sc_hd__and3_1 _20077_ (.A(_10101_),
    .B(_10102_),
    .C(_10103_),
    .X(_10104_));
 sky130_fd_sc_hd__nand3_2 _20078_ (.A(_10101_),
    .B(_10102_),
    .C(_10103_),
    .Y(_10106_));
 sky130_fd_sc_hd__o21ai_1 _20079_ (.A1(_09818_),
    .A2(_09825_),
    .B1(_10100_),
    .Y(_10107_));
 sky130_fd_sc_hd__o21a_1 _20080_ (.A1(_10099_),
    .A2(_10107_),
    .B1(_10106_),
    .X(_10108_));
 sky130_fd_sc_hd__xor2_2 _20081_ (.A(_09838_),
    .B(_10108_),
    .X(net102));
 sky130_fd_sc_hd__a21oi_2 _20082_ (.A1(_10083_),
    .A2(_10087_),
    .B1(_10085_),
    .Y(_10109_));
 sky130_fd_sc_hd__o31a_1 _20083_ (.A1(_09574_),
    .A2(_10064_),
    .A3(_10066_),
    .B1(_10065_),
    .X(_10110_));
 sky130_fd_sc_hd__a31oi_2 _20084_ (.A1(_09979_),
    .A2(_10075_),
    .A3(_10077_),
    .B1(_09976_),
    .Y(_10111_));
 sky130_fd_sc_hd__a31oi_1 _20085_ (.A1(_09977_),
    .A2(_10070_),
    .A3(_10072_),
    .B1(_09978_),
    .Y(_10112_));
 sky130_fd_sc_hd__a31o_1 _20086_ (.A1(_09854_),
    .A2(_09856_),
    .A3(_09845_),
    .B1(_09657_),
    .X(_10113_));
 sky130_fd_sc_hd__nand2_1 _20087_ (.A(net38),
    .B(net24),
    .Y(_10114_));
 sky130_fd_sc_hd__o21ai_4 _20088_ (.A1(net36),
    .A2(net37),
    .B1(net25),
    .Y(_10116_));
 sky130_fd_sc_hd__o21a_2 _20089_ (.A1(net36),
    .A2(net37),
    .B1(net25),
    .X(_10117_));
 sky130_fd_sc_hd__and3_4 _20090_ (.A(net36),
    .B(net37),
    .C(net25),
    .X(_10118_));
 sky130_fd_sc_hd__nand3_4 _20091_ (.A(net36),
    .B(net37),
    .C(net25),
    .Y(_10119_));
 sky130_fd_sc_hd__nand3_1 _20092_ (.A(_10114_),
    .B(_10117_),
    .C(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__o21bai_1 _20093_ (.A1(_10116_),
    .A2(_10118_),
    .B1_N(_10114_),
    .Y(_10121_));
 sky130_fd_sc_hd__o2bb2a_1 _20094_ (.A1_N(net38),
    .A2_N(net24),
    .B1(_10116_),
    .B2(_10118_),
    .X(_10122_));
 sky130_fd_sc_hd__a22o_1 _20095_ (.A1(net38),
    .A2(net24),
    .B1(_10117_),
    .B2(_10119_),
    .X(_10123_));
 sky130_fd_sc_hd__nand4_4 _20096_ (.A(_10117_),
    .B(_10119_),
    .C(net38),
    .D(net24),
    .Y(_10124_));
 sky130_fd_sc_hd__nand2_1 _20097_ (.A(_10124_),
    .B(_09845_),
    .Y(_10125_));
 sky130_fd_sc_hd__and3_1 _20098_ (.A(_10123_),
    .B(_10124_),
    .C(_09845_),
    .X(_10127_));
 sky130_fd_sc_hd__o2111ai_4 _20099_ (.A1(_09346_),
    .A2(_09649_),
    .B1(_09658_),
    .C1(_10123_),
    .D1(_10124_),
    .Y(_10128_));
 sky130_fd_sc_hd__o211ai_4 _20100_ (.A1(_09657_),
    .A2(_09844_),
    .B1(_10120_),
    .C1(_10121_),
    .Y(_10129_));
 sky130_fd_sc_hd__o21ai_2 _20101_ (.A1(_10122_),
    .A2(_10125_),
    .B1(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__nand4_4 _20102_ (.A(_08652_),
    .B(_09340_),
    .C(_10128_),
    .D(_10129_),
    .Y(_10131_));
 sky130_fd_sc_hd__inv_2 _20103_ (.A(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__o21ai_2 _20104_ (.A1(_08651_),
    .A2(_09339_),
    .B1(_10130_),
    .Y(_10133_));
 sky130_fd_sc_hd__a21oi_1 _20105_ (.A1(_10131_),
    .A2(_10133_),
    .B1(_10113_),
    .Y(_10134_));
 sky130_fd_sc_hd__a21o_1 _20106_ (.A1(_10131_),
    .A2(_10133_),
    .B1(_10113_),
    .X(_10135_));
 sky130_fd_sc_hd__and3_1 _20107_ (.A(_10113_),
    .B(_10131_),
    .C(_10133_),
    .X(_10136_));
 sky130_fd_sc_hd__o211ai_4 _20108_ (.A1(_09657_),
    .A2(_09859_),
    .B1(_10131_),
    .C1(_10133_),
    .Y(_10138_));
 sky130_fd_sc_hd__o21ai_2 _20109_ (.A1(_10134_),
    .A2(_10136_),
    .B1(_09388_),
    .Y(_10139_));
 sky130_fd_sc_hd__nand4_4 _20110_ (.A(_09384_),
    .B(_09386_),
    .C(_10135_),
    .D(_10138_),
    .Y(_10140_));
 sky130_fd_sc_hd__a22oi_1 _20111_ (.A1(_08963_),
    .A2(_08006_),
    .B1(_09867_),
    .B2(_09866_),
    .Y(_10141_));
 sky130_fd_sc_hd__o21ai_1 _20112_ (.A1(_09383_),
    .A2(_09868_),
    .B1(_09386_),
    .Y(_10142_));
 sky130_fd_sc_hd__and3_1 _20113_ (.A(_10142_),
    .B(_10140_),
    .C(_10139_),
    .X(_10143_));
 sky130_fd_sc_hd__o211ai_4 _20114_ (.A1(_09385_),
    .A2(_09871_),
    .B1(_10139_),
    .C1(_10140_),
    .Y(_10144_));
 sky130_fd_sc_hd__o2bb2ai_2 _20115_ (.A1_N(_10139_),
    .A2_N(_10140_),
    .B1(_10141_),
    .B2(_09383_),
    .Y(_10145_));
 sky130_fd_sc_hd__nand2_1 _20116_ (.A(_10144_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__o31a_1 _20117_ (.A1(_09342_),
    .A2(_09857_),
    .A3(_09859_),
    .B1(_09866_),
    .X(_10147_));
 sky130_fd_sc_hd__a31o_1 _20118_ (.A1(_09341_),
    .A2(_09858_),
    .A3(_09860_),
    .B1(_09865_),
    .X(_10149_));
 sky130_fd_sc_hd__o21ai_2 _20119_ (.A1(_09885_),
    .A2(_09889_),
    .B1(_09888_),
    .Y(_10150_));
 sky130_fd_sc_hd__o22a_1 _20120_ (.A1(_09729_),
    .A2(_09887_),
    .B1(_09885_),
    .B2(_09889_),
    .X(_10151_));
 sky130_fd_sc_hd__nand2_1 _20121_ (.A(net45),
    .B(net17),
    .Y(_10152_));
 sky130_fd_sc_hd__a22oi_4 _20122_ (.A1(net43),
    .A2(net18),
    .B1(net19),
    .B2(net42),
    .Y(_10153_));
 sky130_fd_sc_hd__a22o_1 _20123_ (.A1(net43),
    .A2(net18),
    .B1(net19),
    .B2(net42),
    .X(_10154_));
 sky130_fd_sc_hd__and4_1 _20124_ (.A(net42),
    .B(net43),
    .C(net18),
    .D(net19),
    .X(_10155_));
 sky130_fd_sc_hd__nand4_2 _20125_ (.A(net42),
    .B(net43),
    .C(net18),
    .D(net19),
    .Y(_10156_));
 sky130_fd_sc_hd__nand3_2 _20126_ (.A(_10152_),
    .B(_10154_),
    .C(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__o21bai_2 _20127_ (.A1(_10153_),
    .A2(_10155_),
    .B1_N(_10152_),
    .Y(_10158_));
 sky130_fd_sc_hd__o21ai_1 _20128_ (.A1(_10153_),
    .A2(_10155_),
    .B1(_10152_),
    .Y(_10160_));
 sky130_fd_sc_hd__and4_1 _20129_ (.A(_10154_),
    .B(_10156_),
    .C(net45),
    .D(net17),
    .X(_10161_));
 sky130_fd_sc_hd__nand4_1 _20130_ (.A(_10154_),
    .B(_10156_),
    .C(net45),
    .D(net17),
    .Y(_10162_));
 sky130_fd_sc_hd__a21oi_1 _20131_ (.A1(_10160_),
    .A2(_10162_),
    .B1(_10150_),
    .Y(_10163_));
 sky130_fd_sc_hd__nand3_1 _20132_ (.A(_10151_),
    .B(_10157_),
    .C(_10158_),
    .Y(_10164_));
 sky130_fd_sc_hd__nand2_1 _20133_ (.A(_10160_),
    .B(_10150_),
    .Y(_10165_));
 sky130_fd_sc_hd__and3_1 _20134_ (.A(_10160_),
    .B(_10162_),
    .C(_10150_),
    .X(_10166_));
 sky130_fd_sc_hd__nand3_1 _20135_ (.A(_10160_),
    .B(_10162_),
    .C(_10150_),
    .Y(_10167_));
 sky130_fd_sc_hd__nand2_1 _20136_ (.A(_10164_),
    .B(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__nand2_1 _20137_ (.A(net14),
    .B(net48),
    .Y(_10169_));
 sky130_fd_sc_hd__nand4_4 _20138_ (.A(net46),
    .B(net15),
    .C(net47),
    .D(net16),
    .Y(_10171_));
 sky130_fd_sc_hd__a22oi_1 _20139_ (.A1(net15),
    .A2(net47),
    .B1(net16),
    .B2(net46),
    .Y(_10172_));
 sky130_fd_sc_hd__a22o_2 _20140_ (.A1(net15),
    .A2(net47),
    .B1(net16),
    .B2(net46),
    .X(_10173_));
 sky130_fd_sc_hd__o211ai_4 _20141_ (.A1(_02065_),
    .A2(_02109_),
    .B1(_10171_),
    .C1(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__a21o_1 _20142_ (.A1(_10171_),
    .A2(_10173_),
    .B1(_10169_),
    .X(_10175_));
 sky130_fd_sc_hd__a22o_1 _20143_ (.A1(net14),
    .A2(net48),
    .B1(_10171_),
    .B2(_10173_),
    .X(_10176_));
 sky130_fd_sc_hd__nand4_2 _20144_ (.A(_10173_),
    .B(net48),
    .C(net14),
    .D(_10171_),
    .Y(_10177_));
 sky130_fd_sc_hd__nand2_1 _20145_ (.A(_10176_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__a32oi_4 _20146_ (.A1(_10151_),
    .A2(_10157_),
    .A3(_10158_),
    .B1(_10174_),
    .B2(_10175_),
    .Y(_10179_));
 sky130_fd_sc_hd__and4_2 _20147_ (.A(_10164_),
    .B(_10167_),
    .C(_10176_),
    .D(_10177_),
    .X(_10180_));
 sky130_fd_sc_hd__and3_2 _20148_ (.A(_10168_),
    .B(_10174_),
    .C(_10175_),
    .X(_10182_));
 sky130_fd_sc_hd__and3_2 _20149_ (.A(_10178_),
    .B(_10167_),
    .C(_10164_),
    .X(_10183_));
 sky130_fd_sc_hd__a211o_1 _20150_ (.A1(_10176_),
    .A2(_10177_),
    .B1(_10163_),
    .C1(_10166_),
    .X(_10184_));
 sky130_fd_sc_hd__and3_2 _20151_ (.A(_10168_),
    .B(_10176_),
    .C(_10177_),
    .X(_10185_));
 sky130_fd_sc_hd__a22o_1 _20152_ (.A1(_10164_),
    .A2(_10167_),
    .B1(_10174_),
    .B2(_10175_),
    .X(_10186_));
 sky130_fd_sc_hd__a21o_1 _20153_ (.A1(_09935_),
    .A2(_09917_),
    .B1(_09932_),
    .X(_10187_));
 sky130_fd_sc_hd__o2bb2a_1 _20154_ (.A1_N(net38),
    .A2_N(net22),
    .B1(_09635_),
    .B2(_09848_),
    .X(_10188_));
 sky130_fd_sc_hd__o2bb2ai_1 _20155_ (.A1_N(_09851_),
    .A2_N(_09847_),
    .B1(_09635_),
    .B2(_09848_),
    .Y(_10189_));
 sky130_fd_sc_hd__nand2_1 _20156_ (.A(net40),
    .B(net22),
    .Y(_10190_));
 sky130_fd_sc_hd__nand2_4 _20157_ (.A(net39),
    .B(net22),
    .Y(_10191_));
 sky130_fd_sc_hd__and4_1 _20158_ (.A(net39),
    .B(net40),
    .C(net21),
    .D(net22),
    .X(_10193_));
 sky130_fd_sc_hd__nand4_1 _20159_ (.A(net39),
    .B(net40),
    .C(net21),
    .D(net22),
    .Y(_10194_));
 sky130_fd_sc_hd__a22oi_4 _20160_ (.A1(net40),
    .A2(net21),
    .B1(net22),
    .B2(net39),
    .Y(_10195_));
 sky130_fd_sc_hd__a22o_2 _20161_ (.A1(net40),
    .A2(net21),
    .B1(net22),
    .B2(net39),
    .X(_10196_));
 sky130_fd_sc_hd__a2bb2oi_1 _20162_ (.A1_N(_02010_),
    .A2_N(_02163_),
    .B1(_10194_),
    .B2(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__o22ai_2 _20163_ (.A1(_02010_),
    .A2(_02163_),
    .B1(_10193_),
    .B2(_10195_),
    .Y(_10198_));
 sky130_fd_sc_hd__o2111a_1 _20164_ (.A1(_09922_),
    .A2(_10190_),
    .B1(net41),
    .C1(net20),
    .D1(_10196_),
    .X(_10199_));
 sky130_fd_sc_hd__o2111ai_4 _20165_ (.A1(_09922_),
    .A2(_10190_),
    .B1(net41),
    .C1(net20),
    .D1(_10196_),
    .Y(_10200_));
 sky130_fd_sc_hd__o22ai_4 _20166_ (.A1(_09846_),
    .A2(_10188_),
    .B1(_10197_),
    .B2(_10199_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand3_4 _20167_ (.A(_10198_),
    .B(_10200_),
    .C(_10189_),
    .Y(_10202_));
 sky130_fd_sc_hd__o22a_1 _20168_ (.A1(_02010_),
    .A2(_02142_),
    .B1(_09697_),
    .B2(_09925_),
    .X(_10204_));
 sky130_fd_sc_hd__a2bb2o_1 _20169_ (.A1_N(_09697_),
    .A2_N(_09925_),
    .B1(_09921_),
    .B2(_09924_),
    .X(_10205_));
 sky130_fd_sc_hd__o2bb2ai_4 _20170_ (.A1_N(_10201_),
    .A2_N(_10202_),
    .B1(_10204_),
    .B2(_09923_),
    .Y(_10206_));
 sky130_fd_sc_hd__and3_2 _20171_ (.A(_10201_),
    .B(_10202_),
    .C(_10205_),
    .X(_10207_));
 sky130_fd_sc_hd__nand3_4 _20172_ (.A(_10201_),
    .B(_10202_),
    .C(_10205_),
    .Y(_10208_));
 sky130_fd_sc_hd__a21oi_4 _20173_ (.A1(_10206_),
    .A2(_10208_),
    .B1(_10187_),
    .Y(_10209_));
 sky130_fd_sc_hd__a21o_1 _20174_ (.A1(_10206_),
    .A2(_10208_),
    .B1(_10187_),
    .X(_10210_));
 sky130_fd_sc_hd__o21ai_2 _20175_ (.A1(_09932_),
    .A2(_09936_),
    .B1(_10206_),
    .Y(_10211_));
 sky130_fd_sc_hd__o211a_2 _20176_ (.A1(_09932_),
    .A2(_09936_),
    .B1(_10206_),
    .C1(_10208_),
    .X(_10212_));
 sky130_fd_sc_hd__nand3_1 _20177_ (.A(_10187_),
    .B(_10206_),
    .C(_10208_),
    .Y(_10213_));
 sky130_fd_sc_hd__o221ai_4 _20178_ (.A1(_10183_),
    .A2(_10185_),
    .B1(_10207_),
    .B2(_10211_),
    .C1(_10210_),
    .Y(_10215_));
 sky130_fd_sc_hd__o22ai_4 _20179_ (.A1(_10180_),
    .A2(_10182_),
    .B1(_10209_),
    .B2(_10212_),
    .Y(_10216_));
 sky130_fd_sc_hd__o22ai_4 _20180_ (.A1(_10183_),
    .A2(_10185_),
    .B1(_10209_),
    .B2(_10212_),
    .Y(_10217_));
 sky130_fd_sc_hd__o221ai_4 _20181_ (.A1(_10180_),
    .A2(_10182_),
    .B1(_10207_),
    .B2(_10211_),
    .C1(_10210_),
    .Y(_10218_));
 sky130_fd_sc_hd__o211a_1 _20182_ (.A1(_09862_),
    .A2(_09865_),
    .B1(_10215_),
    .C1(_10216_),
    .X(_10219_));
 sky130_fd_sc_hd__o211ai_4 _20183_ (.A1(_09862_),
    .A2(_09865_),
    .B1(_10215_),
    .C1(_10216_),
    .Y(_10220_));
 sky130_fd_sc_hd__nand3_2 _20184_ (.A(_10217_),
    .B(_10218_),
    .C(_10147_),
    .Y(_10221_));
 sky130_fd_sc_hd__o32a_1 _20185_ (.A1(_09938_),
    .A2(_09940_),
    .A3(_09914_),
    .B1(_09910_),
    .B2(_09909_),
    .X(_10222_));
 sky130_fd_sc_hd__o21ai_1 _20186_ (.A1(_09909_),
    .A2(_09910_),
    .B1(_09945_),
    .Y(_10223_));
 sky130_fd_sc_hd__o31a_1 _20187_ (.A1(_09911_),
    .A2(_09912_),
    .A3(_09944_),
    .B1(_09947_),
    .X(_10224_));
 sky130_fd_sc_hd__nand2_1 _20188_ (.A(_09947_),
    .B(_10223_),
    .Y(_10226_));
 sky130_fd_sc_hd__a21o_1 _20189_ (.A1(_10220_),
    .A2(_10221_),
    .B1(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__o211ai_2 _20190_ (.A1(_09946_),
    .A2(_10222_),
    .B1(_10221_),
    .C1(_10220_),
    .Y(_10228_));
 sky130_fd_sc_hd__o2bb2ai_2 _20191_ (.A1_N(_10220_),
    .A2_N(_10221_),
    .B1(_10222_),
    .B2(_09946_),
    .Y(_10229_));
 sky130_fd_sc_hd__a31oi_4 _20192_ (.A1(_10217_),
    .A2(_10218_),
    .A3(_10147_),
    .B1(_10226_),
    .Y(_10230_));
 sky130_fd_sc_hd__nand2_2 _20193_ (.A(_10230_),
    .B(_10220_),
    .Y(_10231_));
 sky130_fd_sc_hd__nand3_4 _20194_ (.A(_10146_),
    .B(_10227_),
    .C(_10228_),
    .Y(_10232_));
 sky130_fd_sc_hd__nand4_4 _20195_ (.A(_10144_),
    .B(_10145_),
    .C(_10229_),
    .D(_10231_),
    .Y(_10233_));
 sky130_fd_sc_hd__a22oi_1 _20196_ (.A1(_09841_),
    .A2(_09873_),
    .B1(_09965_),
    .B2(_09968_),
    .Y(_10234_));
 sky130_fd_sc_hd__a32o_1 _20197_ (.A1(_09841_),
    .A2(_09870_),
    .A3(_09872_),
    .B1(_09965_),
    .B2(_09968_),
    .X(_10235_));
 sky130_fd_sc_hd__a22oi_2 _20198_ (.A1(_10232_),
    .A2(_10233_),
    .B1(_10235_),
    .B2(_09874_),
    .Y(_10237_));
 sky130_fd_sc_hd__o2bb2ai_2 _20199_ (.A1_N(_10232_),
    .A2_N(_10233_),
    .B1(_10234_),
    .B2(_09876_),
    .Y(_10238_));
 sky130_fd_sc_hd__o2111a_1 _20200_ (.A1(_09877_),
    .A2(_09969_),
    .B1(_10232_),
    .C1(_10233_),
    .D1(_09874_),
    .X(_10239_));
 sky130_fd_sc_hd__o2111ai_4 _20201_ (.A1(_09877_),
    .A2(_09969_),
    .B1(_10232_),
    .C1(_10233_),
    .D1(_09874_),
    .Y(_10240_));
 sky130_fd_sc_hd__a31o_1 _20202_ (.A1(_09882_),
    .A2(_09950_),
    .A3(_09953_),
    .B1(_09959_),
    .X(_10241_));
 sky130_fd_sc_hd__nor2_1 _20203_ (.A(_09900_),
    .B(_09903_),
    .Y(_10242_));
 sky130_fd_sc_hd__o21a_1 _20204_ (.A1(_09900_),
    .A2(_09903_),
    .B1(_09902_),
    .X(_10243_));
 sky130_fd_sc_hd__nor2_1 _20205_ (.A(_02021_),
    .B(_02152_),
    .Y(_10244_));
 sky130_fd_sc_hd__a22oi_4 _20206_ (.A1(net13),
    .A2(net49),
    .B1(net50),
    .B2(net11),
    .Y(_10245_));
 sky130_fd_sc_hd__a22o_1 _20207_ (.A1(net13),
    .A2(net49),
    .B1(net50),
    .B2(net11),
    .X(_10246_));
 sky130_fd_sc_hd__and4_1 _20208_ (.A(net11),
    .B(net13),
    .C(net49),
    .D(net50),
    .X(_10248_));
 sky130_fd_sc_hd__nand4_2 _20209_ (.A(net11),
    .B(net13),
    .C(net49),
    .D(net50),
    .Y(_10249_));
 sky130_fd_sc_hd__o211ai_1 _20210_ (.A1(_02021_),
    .A2(_02152_),
    .B1(_10246_),
    .C1(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__o21ai_1 _20211_ (.A1(_10245_),
    .A2(_10248_),
    .B1(_10244_),
    .Y(_10251_));
 sky130_fd_sc_hd__o22ai_2 _20212_ (.A1(_02021_),
    .A2(_02152_),
    .B1(_10245_),
    .B2(_10248_),
    .Y(_10252_));
 sky130_fd_sc_hd__nand4_2 _20213_ (.A(_10246_),
    .B(_10249_),
    .C(net10),
    .D(net51),
    .Y(_10253_));
 sky130_fd_sc_hd__nand3_2 _20214_ (.A(_10243_),
    .B(_10250_),
    .C(_10251_),
    .Y(_10254_));
 sky130_fd_sc_hd__o211a_1 _20215_ (.A1(_09901_),
    .A2(_10242_),
    .B1(_10252_),
    .C1(_10253_),
    .X(_10255_));
 sky130_fd_sc_hd__o211ai_4 _20216_ (.A1(_09901_),
    .A2(_10242_),
    .B1(_10252_),
    .C1(_10253_),
    .Y(_10256_));
 sky130_fd_sc_hd__o21a_1 _20217_ (.A1(_01999_),
    .A2(_02152_),
    .B1(_09994_),
    .X(_10257_));
 sky130_fd_sc_hd__a31o_1 _20218_ (.A1(_09992_),
    .A2(net51),
    .A3(net9),
    .B1(_09993_),
    .X(_10259_));
 sky130_fd_sc_hd__o2bb2ai_2 _20219_ (.A1_N(_10254_),
    .A2_N(_10256_),
    .B1(_10257_),
    .B2(_09991_),
    .Y(_10260_));
 sky130_fd_sc_hd__nand2_1 _20220_ (.A(_10254_),
    .B(_10259_),
    .Y(_10261_));
 sky130_fd_sc_hd__nand3_2 _20221_ (.A(_10254_),
    .B(_10256_),
    .C(_10259_),
    .Y(_10262_));
 sky130_fd_sc_hd__o22ai_4 _20222_ (.A1(_09893_),
    .A2(_09898_),
    .B1(_09907_),
    .B2(_09895_),
    .Y(_10263_));
 sky130_fd_sc_hd__a21oi_2 _20223_ (.A1(_10260_),
    .A2(_10262_),
    .B1(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__a21o_1 _20224_ (.A1(_10260_),
    .A2(_10262_),
    .B1(_10263_),
    .X(_10265_));
 sky130_fd_sc_hd__o211a_1 _20225_ (.A1(_10255_),
    .A2(_10261_),
    .B1(_10263_),
    .C1(_10260_),
    .X(_10266_));
 sky130_fd_sc_hd__o211ai_2 _20226_ (.A1(_10255_),
    .A2(_10261_),
    .B1(_10263_),
    .C1(_10260_),
    .Y(_10267_));
 sky130_fd_sc_hd__a21oi_1 _20227_ (.A1(_10003_),
    .A2(_09983_),
    .B1(_10000_),
    .Y(_10268_));
 sky130_fd_sc_hd__o211ai_2 _20228_ (.A1(_10000_),
    .A2(_10004_),
    .B1(_10265_),
    .C1(_10267_),
    .Y(_10270_));
 sky130_fd_sc_hd__o21ai_1 _20229_ (.A1(_10264_),
    .A2(_10266_),
    .B1(_10268_),
    .Y(_10271_));
 sky130_fd_sc_hd__nand3_1 _20230_ (.A(_10265_),
    .B(_10267_),
    .C(_10268_),
    .Y(_10272_));
 sky130_fd_sc_hd__o22ai_2 _20231_ (.A1(_10000_),
    .A2(_10004_),
    .B1(_10264_),
    .B2(_10266_),
    .Y(_10273_));
 sky130_fd_sc_hd__o21ai_1 _20232_ (.A1(_10014_),
    .A2(_10010_),
    .B1(_10013_),
    .Y(_10274_));
 sky130_fd_sc_hd__o2111ai_4 _20233_ (.A1(_10014_),
    .A2(_10010_),
    .B1(_10013_),
    .C1(_10272_),
    .D1(_10273_),
    .Y(_10275_));
 sky130_fd_sc_hd__inv_2 _20234_ (.A(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__nand3_4 _20235_ (.A(_10274_),
    .B(_10271_),
    .C(_10270_),
    .Y(_10277_));
 sky130_fd_sc_hd__o2bb2ai_2 _20236_ (.A1_N(_10043_),
    .A2_N(_10037_),
    .B1(_10035_),
    .B2(_10038_),
    .Y(_10278_));
 sky130_fd_sc_hd__a31o_1 _20237_ (.A1(_10032_),
    .A2(net54),
    .A3(net6),
    .B1(_10030_),
    .X(_10279_));
 sky130_fd_sc_hd__nand2_1 _20238_ (.A(net7),
    .B(net54),
    .Y(_10281_));
 sky130_fd_sc_hd__a22oi_2 _20239_ (.A1(net9),
    .A2(net52),
    .B1(net53),
    .B2(net8),
    .Y(_10282_));
 sky130_fd_sc_hd__a22o_1 _20240_ (.A1(net9),
    .A2(net52),
    .B1(net53),
    .B2(net8),
    .X(_10283_));
 sky130_fd_sc_hd__and4_1 _20241_ (.A(net8),
    .B(net9),
    .C(net52),
    .D(net53),
    .X(_10284_));
 sky130_fd_sc_hd__nand4_2 _20242_ (.A(net8),
    .B(net9),
    .C(net52),
    .D(net53),
    .Y(_10285_));
 sky130_fd_sc_hd__o211ai_1 _20243_ (.A1(_01977_),
    .A2(_02207_),
    .B1(_10283_),
    .C1(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__o21bai_1 _20244_ (.A1(_10282_),
    .A2(_10284_),
    .B1_N(_10281_),
    .Y(_10287_));
 sky130_fd_sc_hd__and4_1 _20245_ (.A(_10283_),
    .B(_10285_),
    .C(net7),
    .D(net54),
    .X(_10288_));
 sky130_fd_sc_hd__nand4_1 _20246_ (.A(_10283_),
    .B(_10285_),
    .C(net7),
    .D(net54),
    .Y(_10289_));
 sky130_fd_sc_hd__o21ai_1 _20247_ (.A1(_10282_),
    .A2(_10284_),
    .B1(_10281_),
    .Y(_10290_));
 sky130_fd_sc_hd__o21ai_1 _20248_ (.A1(_10030_),
    .A2(_10035_),
    .B1(_10290_),
    .Y(_10292_));
 sky130_fd_sc_hd__nand3_1 _20249_ (.A(_10279_),
    .B(_10289_),
    .C(_10290_),
    .Y(_10293_));
 sky130_fd_sc_hd__nand4_2 _20250_ (.A(_10031_),
    .B(_10036_),
    .C(_10286_),
    .D(_10287_),
    .Y(_10294_));
 sky130_fd_sc_hd__and4_2 _20251_ (.A(_01956_),
    .B(net6),
    .C(net56),
    .D(net57),
    .X(_10295_));
 sky130_fd_sc_hd__or4_2 _20252_ (.A(net5),
    .B(_01966_),
    .C(_02229_),
    .D(_02240_),
    .X(_10296_));
 sky130_fd_sc_hd__o22a_1 _20253_ (.A1(net5),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01966_),
    .X(_10297_));
 sky130_fd_sc_hd__nor2_1 _20254_ (.A(_10295_),
    .B(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__o2bb2ai_1 _20255_ (.A1_N(_10293_),
    .A2_N(_10294_),
    .B1(_10295_),
    .B2(_10297_),
    .Y(_10299_));
 sky130_fd_sc_hd__nand3_1 _20256_ (.A(_10293_),
    .B(_10294_),
    .C(_10298_),
    .Y(_10300_));
 sky130_fd_sc_hd__a21oi_2 _20257_ (.A1(_10299_),
    .A2(_10300_),
    .B1(_10278_),
    .Y(_10301_));
 sky130_fd_sc_hd__a21o_1 _20258_ (.A1(_10299_),
    .A2(_10300_),
    .B1(_10278_),
    .X(_10303_));
 sky130_fd_sc_hd__and3_4 _20259_ (.A(_10278_),
    .B(_10299_),
    .C(_10300_),
    .X(_10304_));
 sky130_fd_sc_hd__o21ba_1 _20260_ (.A1(_10301_),
    .A2(_10304_),
    .B1_N(_10041_),
    .X(_10305_));
 sky130_fd_sc_hd__o21bai_2 _20261_ (.A1(_10301_),
    .A2(_10304_),
    .B1_N(_10041_),
    .Y(_10306_));
 sky130_fd_sc_hd__nand2_1 _20262_ (.A(_10303_),
    .B(_10041_),
    .Y(_10307_));
 sky130_fd_sc_hd__nor2_1 _20263_ (.A(_10304_),
    .B(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__nor3_1 _20264_ (.A(_10041_),
    .B(_10301_),
    .C(_10304_),
    .Y(_10309_));
 sky130_fd_sc_hd__o21a_1 _20265_ (.A1(_10301_),
    .A2(_10304_),
    .B1(_10041_),
    .X(_10310_));
 sky130_fd_sc_hd__o21ai_1 _20266_ (.A1(_10304_),
    .A2(_10307_),
    .B1(_10306_),
    .Y(_10311_));
 sky130_fd_sc_hd__o2bb2ai_2 _20267_ (.A1_N(_10275_),
    .A2_N(_10277_),
    .B1(_10309_),
    .B2(_10310_),
    .Y(_10312_));
 sky130_fd_sc_hd__nand3_2 _20268_ (.A(_10275_),
    .B(_10277_),
    .C(_10311_),
    .Y(_10314_));
 sky130_fd_sc_hd__o2111ai_4 _20269_ (.A1(_10304_),
    .A2(_10307_),
    .B1(_10306_),
    .C1(_10275_),
    .D1(_10277_),
    .Y(_10315_));
 sky130_fd_sc_hd__o2bb2ai_1 _20270_ (.A1_N(_10275_),
    .A2_N(_10277_),
    .B1(_10305_),
    .B2(_10308_),
    .Y(_10316_));
 sky130_fd_sc_hd__a22oi_2 _20271_ (.A1(_09955_),
    .A2(_09966_),
    .B1(_10312_),
    .B2(_10314_),
    .Y(_10317_));
 sky130_fd_sc_hd__nand4_4 _20272_ (.A(_09957_),
    .B(_10241_),
    .C(_10315_),
    .D(_10316_),
    .Y(_10318_));
 sky130_fd_sc_hd__o2111a_1 _20273_ (.A1(_09960_),
    .A2(_09956_),
    .B1(_09955_),
    .C1(_10314_),
    .D1(_10312_),
    .X(_10319_));
 sky130_fd_sc_hd__o2111ai_4 _20274_ (.A1(_09960_),
    .A2(_09956_),
    .B1(_09955_),
    .C1(_10314_),
    .D1(_10312_),
    .Y(_10320_));
 sky130_fd_sc_hd__o21a_1 _20275_ (.A1(_10052_),
    .A2(_10053_),
    .B1(_10025_),
    .X(_10321_));
 sky130_fd_sc_hd__nor2_1 _20276_ (.A(_10024_),
    .B(_10056_),
    .Y(_10322_));
 sky130_fd_sc_hd__a21oi_1 _20277_ (.A1(_10318_),
    .A2(_10320_),
    .B1(_10322_),
    .Y(_10323_));
 sky130_fd_sc_hd__o22ai_2 _20278_ (.A1(_10024_),
    .A2(_10056_),
    .B1(_10317_),
    .B2(_10319_),
    .Y(_10325_));
 sky130_fd_sc_hd__and3_1 _20279_ (.A(_10318_),
    .B(_10320_),
    .C(_10322_),
    .X(_10326_));
 sky130_fd_sc_hd__o211ai_2 _20280_ (.A1(_10022_),
    .A2(_10321_),
    .B1(_10320_),
    .C1(_10318_),
    .Y(_10327_));
 sky130_fd_sc_hd__a21boi_1 _20281_ (.A1(_10318_),
    .A2(_10320_),
    .B1_N(_10322_),
    .Y(_10328_));
 sky130_fd_sc_hd__o2bb2ai_1 _20282_ (.A1_N(_10318_),
    .A2_N(_10320_),
    .B1(_10321_),
    .B2(_10022_),
    .Y(_10329_));
 sky130_fd_sc_hd__o211a_1 _20283_ (.A1(_10024_),
    .A2(_10056_),
    .B1(_10318_),
    .C1(_10320_),
    .X(_10330_));
 sky130_fd_sc_hd__o211ai_2 _20284_ (.A1(_10024_),
    .A2(_10056_),
    .B1(_10318_),
    .C1(_10320_),
    .Y(_10331_));
 sky130_fd_sc_hd__nand4_1 _20285_ (.A(_10238_),
    .B(_10240_),
    .C(_10325_),
    .D(_10327_),
    .Y(_10332_));
 sky130_fd_sc_hd__o2bb2ai_1 _20286_ (.A1_N(_10238_),
    .A2_N(_10240_),
    .B1(_10323_),
    .B2(_10326_),
    .Y(_10333_));
 sky130_fd_sc_hd__o2bb2ai_1 _20287_ (.A1_N(_10238_),
    .A2_N(_10240_),
    .B1(_10328_),
    .B2(_10330_),
    .Y(_10334_));
 sky130_fd_sc_hd__nand4_1 _20288_ (.A(_10238_),
    .B(_10240_),
    .C(_10329_),
    .D(_10331_),
    .Y(_10336_));
 sky130_fd_sc_hd__nand3_2 _20289_ (.A(_10111_),
    .B(_10334_),
    .C(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__a21oi_1 _20290_ (.A1(_10334_),
    .A2(_10336_),
    .B1(_10111_),
    .Y(_10338_));
 sky130_fd_sc_hd__nand3_2 _20291_ (.A(_10112_),
    .B(_10332_),
    .C(_10333_),
    .Y(_10339_));
 sky130_fd_sc_hd__a22oi_2 _20292_ (.A1(_10065_),
    .A2(_10072_),
    .B1(_10337_),
    .B2(_10339_),
    .Y(_10340_));
 sky130_fd_sc_hd__a22o_1 _20293_ (.A1(_10065_),
    .A2(_10072_),
    .B1(_10337_),
    .B2(_10339_),
    .X(_10341_));
 sky130_fd_sc_hd__o2111a_1 _20294_ (.A1(_10068_),
    .A2(_10064_),
    .B1(_10065_),
    .C1(_10337_),
    .D1(_10339_),
    .X(_10342_));
 sky130_fd_sc_hd__o2111ai_2 _20295_ (.A1(_10068_),
    .A2(_10064_),
    .B1(_10065_),
    .C1(_10337_),
    .D1(_10339_),
    .Y(_10343_));
 sky130_fd_sc_hd__nor2_1 _20296_ (.A(_10340_),
    .B(_10342_),
    .Y(_10344_));
 sky130_fd_sc_hd__nand4_1 _20297_ (.A(_10086_),
    .B(_10092_),
    .C(_10341_),
    .D(_10343_),
    .Y(_10345_));
 sky130_fd_sc_hd__o2bb2a_1 _20298_ (.A1_N(_10086_),
    .A2_N(_10092_),
    .B1(_10340_),
    .B2(_10342_),
    .X(_10347_));
 sky130_fd_sc_hd__o21bai_1 _20299_ (.A1(_10340_),
    .A2(_10342_),
    .B1_N(_10109_),
    .Y(_10348_));
 sky130_fd_sc_hd__o31a_1 _20300_ (.A1(_01945_),
    .A2(_02229_),
    .A3(_09595_),
    .B1(_10048_),
    .X(_10349_));
 sky130_fd_sc_hd__o41a_1 _20301_ (.A1(net3),
    .A2(_02240_),
    .A3(_09594_),
    .A4(_10049_),
    .B1(_10048_),
    .X(_10350_));
 sky130_fd_sc_hd__o2bb2ai_1 _20302_ (.A1_N(_10345_),
    .A2_N(_10348_),
    .B1(_10349_),
    .B2(_10049_),
    .Y(_10351_));
 sky130_fd_sc_hd__a31oi_1 _20303_ (.A1(_10341_),
    .A2(_10343_),
    .A3(_10109_),
    .B1(_10350_),
    .Y(_10352_));
 sky130_fd_sc_hd__a31o_1 _20304_ (.A1(_10341_),
    .A2(_10343_),
    .A3(_10109_),
    .B1(_10350_),
    .X(_10353_));
 sky130_fd_sc_hd__a21o_1 _20305_ (.A1(_10345_),
    .A2(_10348_),
    .B1(_10350_),
    .X(_10354_));
 sky130_fd_sc_hd__o211ai_1 _20306_ (.A1(_10049_),
    .A2(_10349_),
    .B1(_10348_),
    .C1(_10345_),
    .Y(_10355_));
 sky130_fd_sc_hd__a31oi_2 _20307_ (.A1(_09607_),
    .A2(_09610_),
    .A3(_10097_),
    .B1(_10094_),
    .Y(_10356_));
 sky130_fd_sc_hd__a21oi_1 _20308_ (.A1(_10095_),
    .A2(_10098_),
    .B1(_10096_),
    .Y(_10358_));
 sky130_fd_sc_hd__nand3_2 _20309_ (.A(_10354_),
    .B(_10355_),
    .C(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__o211ai_4 _20310_ (.A1(_10347_),
    .A2(_10353_),
    .B1(_10351_),
    .C1(_10356_),
    .Y(_10360_));
 sky130_fd_sc_hd__nand2_1 _20311_ (.A(_10359_),
    .B(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__and3_1 _20312_ (.A(_10108_),
    .B(_09831_),
    .C(_09830_),
    .X(_10362_));
 sky130_fd_sc_hd__o2111ai_1 _20313_ (.A1(_10099_),
    .A2(_10107_),
    .B1(_10106_),
    .C1(_09830_),
    .D1(_09831_),
    .Y(_10363_));
 sky130_fd_sc_hd__o21a_1 _20314_ (.A1(_10099_),
    .A2(_10107_),
    .B1(_09831_),
    .X(_10364_));
 sky130_fd_sc_hd__inv_2 _20315_ (.A(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__a22oi_4 _20316_ (.A1(_10106_),
    .A2(_10365_),
    .B1(_09837_),
    .B2(_10362_),
    .Y(_10366_));
 sky130_fd_sc_hd__o2bb2ai_1 _20317_ (.A1_N(_10362_),
    .A2_N(_09837_),
    .B1(_10104_),
    .B2(_10364_),
    .Y(_10367_));
 sky130_fd_sc_hd__nand3_1 _20318_ (.A(_10359_),
    .B(_10360_),
    .C(_10367_),
    .Y(_10369_));
 sky130_fd_sc_hd__xor2_2 _20319_ (.A(_10361_),
    .B(_10366_),
    .X(net103));
 sky130_fd_sc_hd__o21ai_1 _20320_ (.A1(_10110_),
    .A2(_10338_),
    .B1(_10337_),
    .Y(_10370_));
 sky130_fd_sc_hd__a31o_1 _20321_ (.A1(_10065_),
    .A2(_10072_),
    .A3(_10337_),
    .B1(_10338_),
    .X(_10371_));
 sky130_fd_sc_hd__a21o_1 _20322_ (.A1(_10267_),
    .A2(_10268_),
    .B1(_10264_),
    .X(_10372_));
 sky130_fd_sc_hd__a21oi_1 _20323_ (.A1(_10267_),
    .A2(_10268_),
    .B1(_10264_),
    .Y(_10373_));
 sky130_fd_sc_hd__a21oi_2 _20324_ (.A1(_10254_),
    .A2(_10259_),
    .B1(_10255_),
    .Y(_10374_));
 sky130_fd_sc_hd__o21ai_1 _20325_ (.A1(_10169_),
    .A2(_10172_),
    .B1(_10171_),
    .Y(_10375_));
 sky130_fd_sc_hd__o21a_1 _20326_ (.A1(_10169_),
    .A2(_10172_),
    .B1(_10171_),
    .X(_10376_));
 sky130_fd_sc_hd__nand2_1 _20327_ (.A(net11),
    .B(net51),
    .Y(_10377_));
 sky130_fd_sc_hd__a22oi_4 _20328_ (.A1(net14),
    .A2(net49),
    .B1(net50),
    .B2(net13),
    .Y(_10379_));
 sky130_fd_sc_hd__a22o_1 _20329_ (.A1(net14),
    .A2(net49),
    .B1(net50),
    .B2(net13),
    .X(_10380_));
 sky130_fd_sc_hd__and4_1 _20330_ (.A(net13),
    .B(net14),
    .C(net49),
    .D(net50),
    .X(_10381_));
 sky130_fd_sc_hd__nand4_4 _20331_ (.A(net13),
    .B(net14),
    .C(net49),
    .D(net50),
    .Y(_10382_));
 sky130_fd_sc_hd__o211ai_1 _20332_ (.A1(_02032_),
    .A2(_02152_),
    .B1(_10380_),
    .C1(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__o21bai_1 _20333_ (.A1(_10379_),
    .A2(_10381_),
    .B1_N(_10377_),
    .Y(_10384_));
 sky130_fd_sc_hd__a22o_1 _20334_ (.A1(net11),
    .A2(net51),
    .B1(_10380_),
    .B2(_10382_),
    .X(_10385_));
 sky130_fd_sc_hd__nand4_2 _20335_ (.A(_10380_),
    .B(_10382_),
    .C(net11),
    .D(net51),
    .Y(_10386_));
 sky130_fd_sc_hd__nand3_2 _20336_ (.A(_10376_),
    .B(_10383_),
    .C(_10384_),
    .Y(_10387_));
 sky130_fd_sc_hd__nand3_4 _20337_ (.A(_10385_),
    .B(_10386_),
    .C(_10375_),
    .Y(_10388_));
 sky130_fd_sc_hd__o21a_1 _20338_ (.A1(_02021_),
    .A2(_02152_),
    .B1(_10249_),
    .X(_10390_));
 sky130_fd_sc_hd__a31o_1 _20339_ (.A1(_10246_),
    .A2(net51),
    .A3(net10),
    .B1(_10248_),
    .X(_10391_));
 sky130_fd_sc_hd__o2bb2ai_2 _20340_ (.A1_N(_10387_),
    .A2_N(_10388_),
    .B1(_10390_),
    .B2(_10245_),
    .Y(_10392_));
 sky130_fd_sc_hd__nand3_4 _20341_ (.A(_10387_),
    .B(_10388_),
    .C(_10391_),
    .Y(_10393_));
 sky130_fd_sc_hd__o22ai_2 _20342_ (.A1(_10161_),
    .A2(_10165_),
    .B1(_10178_),
    .B2(_10163_),
    .Y(_10394_));
 sky130_fd_sc_hd__a21oi_2 _20343_ (.A1(_10392_),
    .A2(_10393_),
    .B1(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__a21o_1 _20344_ (.A1(_10392_),
    .A2(_10393_),
    .B1(_10394_),
    .X(_10396_));
 sky130_fd_sc_hd__o211a_1 _20345_ (.A1(_10166_),
    .A2(_10179_),
    .B1(_10392_),
    .C1(_10393_),
    .X(_10397_));
 sky130_fd_sc_hd__o211ai_2 _20346_ (.A1(_10166_),
    .A2(_10179_),
    .B1(_10392_),
    .C1(_10393_),
    .Y(_10398_));
 sky130_fd_sc_hd__o21ai_1 _20347_ (.A1(_10395_),
    .A2(_10397_),
    .B1(_10374_),
    .Y(_10399_));
 sky130_fd_sc_hd__nand3b_1 _20348_ (.A_N(_10374_),
    .B(_10396_),
    .C(_10398_),
    .Y(_10401_));
 sky130_fd_sc_hd__nand3_1 _20349_ (.A(_10396_),
    .B(_10398_),
    .C(_10374_),
    .Y(_10402_));
 sky130_fd_sc_hd__o2bb2ai_2 _20350_ (.A1_N(_10256_),
    .A2_N(_10262_),
    .B1(_10395_),
    .B2(_10397_),
    .Y(_10403_));
 sky130_fd_sc_hd__nand3_4 _20351_ (.A(_10372_),
    .B(_10402_),
    .C(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__inv_2 _20352_ (.A(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__nand3_4 _20353_ (.A(_10373_),
    .B(_10399_),
    .C(_10401_),
    .Y(_10406_));
 sky130_fd_sc_hd__o2bb2ai_2 _20354_ (.A1_N(_10298_),
    .A2_N(_10294_),
    .B1(_10288_),
    .B2(_10292_),
    .Y(_10407_));
 sky130_fd_sc_hd__o21ai_1 _20355_ (.A1(_01977_),
    .A2(_02207_),
    .B1(_10285_),
    .Y(_10408_));
 sky130_fd_sc_hd__o31a_1 _20356_ (.A1(_01977_),
    .A2(_02207_),
    .A3(_10282_),
    .B1(_10285_),
    .X(_10409_));
 sky130_fd_sc_hd__nand2_1 _20357_ (.A(net8),
    .B(net54),
    .Y(_10410_));
 sky130_fd_sc_hd__a22oi_2 _20358_ (.A1(net10),
    .A2(net52),
    .B1(net53),
    .B2(net9),
    .Y(_10412_));
 sky130_fd_sc_hd__a22o_1 _20359_ (.A1(net10),
    .A2(net52),
    .B1(net53),
    .B2(net9),
    .X(_10413_));
 sky130_fd_sc_hd__nand2_1 _20360_ (.A(net10),
    .B(net53),
    .Y(_10414_));
 sky130_fd_sc_hd__and4_1 _20361_ (.A(net9),
    .B(net10),
    .C(net52),
    .D(net53),
    .X(_10415_));
 sky130_fd_sc_hd__nand4_1 _20362_ (.A(net9),
    .B(net10),
    .C(net52),
    .D(net53),
    .Y(_10416_));
 sky130_fd_sc_hd__o211ai_1 _20363_ (.A1(_01988_),
    .A2(_02207_),
    .B1(_10413_),
    .C1(_10416_),
    .Y(_10417_));
 sky130_fd_sc_hd__a21o_1 _20364_ (.A1(_10413_),
    .A2(_10416_),
    .B1(_10410_),
    .X(_10418_));
 sky130_fd_sc_hd__nand4_1 _20365_ (.A(_10413_),
    .B(_10416_),
    .C(net8),
    .D(net54),
    .Y(_10419_));
 sky130_fd_sc_hd__o21ai_2 _20366_ (.A1(_10412_),
    .A2(_10415_),
    .B1(_10410_),
    .Y(_10420_));
 sky130_fd_sc_hd__nand4_4 _20367_ (.A(_10283_),
    .B(_10408_),
    .C(_10419_),
    .D(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__nand3_2 _20368_ (.A(_10409_),
    .B(_10417_),
    .C(_10418_),
    .Y(_10423_));
 sky130_fd_sc_hd__nand2_1 _20369_ (.A(_01966_),
    .B(net57),
    .Y(_10424_));
 sky130_fd_sc_hd__and4_1 _20370_ (.A(_01966_),
    .B(net7),
    .C(net56),
    .D(net57),
    .X(_10425_));
 sky130_fd_sc_hd__or4_2 _20371_ (.A(net6),
    .B(_01977_),
    .C(_02229_),
    .D(_02240_),
    .X(_10426_));
 sky130_fd_sc_hd__o22a_1 _20372_ (.A1(net6),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_01977_),
    .X(_10427_));
 sky130_fd_sc_hd__a22o_1 _20373_ (.A1(net7),
    .A2(net56),
    .B1(_01966_),
    .B2(net57),
    .X(_10428_));
 sky130_fd_sc_hd__o2bb2ai_2 _20374_ (.A1_N(_10421_),
    .A2_N(_10423_),
    .B1(_10425_),
    .B2(_10427_),
    .Y(_10429_));
 sky130_fd_sc_hd__nand4_4 _20375_ (.A(_10421_),
    .B(_10423_),
    .C(_10426_),
    .D(_10428_),
    .Y(_10430_));
 sky130_fd_sc_hd__a21oi_2 _20376_ (.A1(_10429_),
    .A2(_10430_),
    .B1(_10407_),
    .Y(_10431_));
 sky130_fd_sc_hd__a21o_1 _20377_ (.A1(_10429_),
    .A2(_10430_),
    .B1(_10407_),
    .X(_10432_));
 sky130_fd_sc_hd__and3_1 _20378_ (.A(_10407_),
    .B(_10429_),
    .C(_10430_),
    .X(_10434_));
 sky130_fd_sc_hd__nand3_2 _20379_ (.A(_10407_),
    .B(_10429_),
    .C(_10430_),
    .Y(_10435_));
 sky130_fd_sc_hd__a21oi_1 _20380_ (.A1(_10432_),
    .A2(_10435_),
    .B1(_10295_),
    .Y(_10436_));
 sky130_fd_sc_hd__o21ai_1 _20381_ (.A1(_10431_),
    .A2(_10434_),
    .B1(_10296_),
    .Y(_10437_));
 sky130_fd_sc_hd__nand2_1 _20382_ (.A(_10432_),
    .B(_10295_),
    .Y(_10438_));
 sky130_fd_sc_hd__and3_1 _20383_ (.A(_10432_),
    .B(_10435_),
    .C(_10295_),
    .X(_10439_));
 sky130_fd_sc_hd__and3_1 _20384_ (.A(_10296_),
    .B(_10432_),
    .C(_10435_),
    .X(_10440_));
 sky130_fd_sc_hd__a21oi_1 _20385_ (.A1(_10432_),
    .A2(_10435_),
    .B1(_10296_),
    .Y(_10441_));
 sky130_fd_sc_hd__o21ai_2 _20386_ (.A1(_10434_),
    .A2(_10438_),
    .B1(_10437_),
    .Y(_10442_));
 sky130_fd_sc_hd__o2111ai_2 _20387_ (.A1(_10434_),
    .A2(_10438_),
    .B1(_10437_),
    .C1(_10404_),
    .D1(_10406_),
    .Y(_10443_));
 sky130_fd_sc_hd__o2bb2ai_1 _20388_ (.A1_N(_10404_),
    .A2_N(_10406_),
    .B1(_10436_),
    .B2(_10439_),
    .Y(_10445_));
 sky130_fd_sc_hd__o2bb2ai_1 _20389_ (.A1_N(_10404_),
    .A2_N(_10406_),
    .B1(_10440_),
    .B2(_10441_),
    .Y(_10446_));
 sky130_fd_sc_hd__o211ai_1 _20390_ (.A1(_10436_),
    .A2(_10439_),
    .B1(_10404_),
    .C1(_10406_),
    .Y(_10447_));
 sky130_fd_sc_hd__a32oi_2 _20391_ (.A1(_10149_),
    .A2(_10215_),
    .A3(_10216_),
    .B1(_10221_),
    .B2(_10224_),
    .Y(_10448_));
 sky130_fd_sc_hd__nand3_2 _20392_ (.A(_10446_),
    .B(_10448_),
    .C(_10447_),
    .Y(_10449_));
 sky130_fd_sc_hd__inv_2 _20393_ (.A(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__o211a_1 _20394_ (.A1(_10219_),
    .A2(_10230_),
    .B1(_10443_),
    .C1(_10445_),
    .X(_10451_));
 sky130_fd_sc_hd__o211ai_2 _20395_ (.A1(_10219_),
    .A2(_10230_),
    .B1(_10443_),
    .C1(_10445_),
    .Y(_10452_));
 sky130_fd_sc_hd__o21a_1 _20396_ (.A1(_10305_),
    .A2(_10308_),
    .B1(_10277_),
    .X(_10453_));
 sky130_fd_sc_hd__nand2_1 _20397_ (.A(_10277_),
    .B(_10315_),
    .Y(_10454_));
 sky130_fd_sc_hd__a21oi_1 _20398_ (.A1(_10449_),
    .A2(_10452_),
    .B1(_10454_),
    .Y(_10456_));
 sky130_fd_sc_hd__o2bb2ai_1 _20399_ (.A1_N(_10449_),
    .A2_N(_10452_),
    .B1(_10453_),
    .B2(_10276_),
    .Y(_10457_));
 sky130_fd_sc_hd__nand2_1 _20400_ (.A(_10449_),
    .B(_10454_),
    .Y(_10458_));
 sky130_fd_sc_hd__and3_1 _20401_ (.A(_10449_),
    .B(_10452_),
    .C(_10454_),
    .X(_10459_));
 sky130_fd_sc_hd__o21ai_1 _20402_ (.A1(_10451_),
    .A2(_10458_),
    .B1(_10457_),
    .Y(_10460_));
 sky130_fd_sc_hd__a31oi_2 _20403_ (.A1(_10145_),
    .A2(_10229_),
    .A3(_10231_),
    .B1(_10143_),
    .Y(_10461_));
 sky130_fd_sc_hd__a31o_1 _20404_ (.A1(_10145_),
    .A2(_10229_),
    .A3(_10231_),
    .B1(_10143_),
    .X(_10462_));
 sky130_fd_sc_hd__o211ai_2 _20405_ (.A1(_08959_),
    .A2(_08004_),
    .B1(_10138_),
    .C1(_10135_),
    .Y(_10463_));
 sky130_fd_sc_hd__o21ai_1 _20406_ (.A1(_08007_),
    .A2(_08962_),
    .B1(_10463_),
    .Y(_10464_));
 sky130_fd_sc_hd__a31o_1 _20407_ (.A1(_10123_),
    .A2(_10124_),
    .A3(_09845_),
    .B1(_09657_),
    .X(_10465_));
 sky130_fd_sc_hd__and2_1 _20408_ (.A(net38),
    .B(net25),
    .X(_10467_));
 sky130_fd_sc_hd__nand2_2 _20409_ (.A(net38),
    .B(net25),
    .Y(_10468_));
 sky130_fd_sc_hd__nor3_2 _20410_ (.A(_10116_),
    .B(_10468_),
    .C(_10118_),
    .Y(_10469_));
 sky130_fd_sc_hd__nand4_4 _20411_ (.A(_10117_),
    .B(_10119_),
    .C(net38),
    .D(net25),
    .Y(_10470_));
 sky130_fd_sc_hd__a21oi_1 _20412_ (.A1(_10117_),
    .A2(_10119_),
    .B1(_10467_),
    .Y(_10471_));
 sky130_fd_sc_hd__o2bb2ai_4 _20413_ (.A1_N(net38),
    .A2_N(net25),
    .B1(_10116_),
    .B2(_10118_),
    .Y(_10472_));
 sky130_fd_sc_hd__a21oi_4 _20414_ (.A1(_10470_),
    .A2(_10472_),
    .B1(_09845_),
    .Y(_10473_));
 sky130_fd_sc_hd__o22ai_2 _20415_ (.A1(_09657_),
    .A2(_09844_),
    .B1(_10469_),
    .B2(_10471_),
    .Y(_10474_));
 sky130_fd_sc_hd__nand2_1 _20416_ (.A(_10472_),
    .B(_09845_),
    .Y(_10475_));
 sky130_fd_sc_hd__and3_2 _20417_ (.A(_10472_),
    .B(_09845_),
    .C(_10470_),
    .X(_10476_));
 sky130_fd_sc_hd__o2111ai_4 _20418_ (.A1(_09346_),
    .A2(_09649_),
    .B1(_09658_),
    .C1(_10470_),
    .D1(_10472_),
    .Y(_10478_));
 sky130_fd_sc_hd__o22ai_4 _20419_ (.A1(_08651_),
    .A2(_09339_),
    .B1(_10473_),
    .B2(_10476_),
    .Y(_10479_));
 sky130_fd_sc_hd__o211ai_4 _20420_ (.A1(_10469_),
    .A2(_10475_),
    .B1(_08652_),
    .C1(_09340_),
    .Y(_10480_));
 sky130_fd_sc_hd__and3_4 _20421_ (.A(_09341_),
    .B(_10474_),
    .C(_10478_),
    .X(_10481_));
 sky130_fd_sc_hd__nand4_4 _20422_ (.A(_08652_),
    .B(_09340_),
    .C(_10474_),
    .D(_10478_),
    .Y(_10482_));
 sky130_fd_sc_hd__o211a_2 _20423_ (.A1(_09657_),
    .A2(_10127_),
    .B1(_10479_),
    .C1(_10482_),
    .X(_10483_));
 sky130_fd_sc_hd__o221ai_4 _20424_ (.A1(_09657_),
    .A2(_10127_),
    .B1(_10473_),
    .B2(_10480_),
    .C1(_10479_),
    .Y(_10484_));
 sky130_fd_sc_hd__a21oi_1 _20425_ (.A1(_10479_),
    .A2(_10482_),
    .B1(_10465_),
    .Y(_10485_));
 sky130_fd_sc_hd__a21o_1 _20426_ (.A1(_10479_),
    .A2(_10482_),
    .B1(_10465_),
    .X(_10486_));
 sky130_fd_sc_hd__o211ai_4 _20427_ (.A1(_09383_),
    .A2(_09385_),
    .B1(_10484_),
    .C1(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__o21ai_2 _20428_ (.A1(_10483_),
    .A2(_10485_),
    .B1(_09387_),
    .Y(_10489_));
 sky130_fd_sc_hd__a22o_1 _20429_ (.A1(_09384_),
    .A2(_09386_),
    .B1(_10484_),
    .B2(_10486_),
    .X(_10490_));
 sky130_fd_sc_hd__nand4_1 _20430_ (.A(_09384_),
    .B(_09386_),
    .C(_10484_),
    .D(_10486_),
    .Y(_10491_));
 sky130_fd_sc_hd__a21oi_1 _20431_ (.A1(_10490_),
    .A2(_10491_),
    .B1(_10464_),
    .Y(_10492_));
 sky130_fd_sc_hd__nand4_4 _20432_ (.A(_09386_),
    .B(_10140_),
    .C(_10487_),
    .D(_10489_),
    .Y(_10493_));
 sky130_fd_sc_hd__a22oi_4 _20433_ (.A1(_09386_),
    .A2(_10463_),
    .B1(_10487_),
    .B2(_10489_),
    .Y(_10494_));
 sky130_fd_sc_hd__nand3_2 _20434_ (.A(_10464_),
    .B(_10490_),
    .C(_10491_),
    .Y(_10495_));
 sky130_fd_sc_hd__nand2_1 _20435_ (.A(_10493_),
    .B(_10495_),
    .Y(_10496_));
 sky130_fd_sc_hd__o31a_2 _20436_ (.A1(_08651_),
    .A2(_09339_),
    .A3(_10130_),
    .B1(_10138_),
    .X(_10497_));
 sky130_fd_sc_hd__o21ai_1 _20437_ (.A1(_09342_),
    .A2(_10130_),
    .B1(_10138_),
    .Y(_10498_));
 sky130_fd_sc_hd__nand2_1 _20438_ (.A(net46),
    .B(net17),
    .Y(_10500_));
 sky130_fd_sc_hd__and4_1 _20439_ (.A(net46),
    .B(net47),
    .C(net16),
    .D(net17),
    .X(_10501_));
 sky130_fd_sc_hd__nand4_1 _20440_ (.A(net46),
    .B(net47),
    .C(net16),
    .D(net17),
    .Y(_10502_));
 sky130_fd_sc_hd__a22o_1 _20441_ (.A1(net47),
    .A2(net16),
    .B1(net17),
    .B2(net46),
    .X(_10503_));
 sky130_fd_sc_hd__a22o_1 _20442_ (.A1(net15),
    .A2(net48),
    .B1(_10502_),
    .B2(_10503_),
    .X(_10504_));
 sky130_fd_sc_hd__nand4_1 _20443_ (.A(_10503_),
    .B(net48),
    .C(net15),
    .D(_10502_),
    .Y(_10505_));
 sky130_fd_sc_hd__nand2_2 _20444_ (.A(_10504_),
    .B(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__o21ai_1 _20445_ (.A1(_10152_),
    .A2(_10153_),
    .B1(_10156_),
    .Y(_10507_));
 sky130_fd_sc_hd__o21a_1 _20446_ (.A1(_10152_),
    .A2(_10153_),
    .B1(_10156_),
    .X(_10508_));
 sky130_fd_sc_hd__nand2_1 _20447_ (.A(net45),
    .B(net18),
    .Y(_10509_));
 sky130_fd_sc_hd__nand2_1 _20448_ (.A(net42),
    .B(net20),
    .Y(_10511_));
 sky130_fd_sc_hd__and4_2 _20449_ (.A(net42),
    .B(net43),
    .C(net19),
    .D(net20),
    .X(_10512_));
 sky130_fd_sc_hd__nand4_2 _20450_ (.A(net42),
    .B(net43),
    .C(net19),
    .D(net20),
    .Y(_10513_));
 sky130_fd_sc_hd__a22oi_4 _20451_ (.A1(net43),
    .A2(net19),
    .B1(net20),
    .B2(net42),
    .Y(_10514_));
 sky130_fd_sc_hd__a22o_1 _20452_ (.A1(net43),
    .A2(net19),
    .B1(net20),
    .B2(net42),
    .X(_10515_));
 sky130_fd_sc_hd__o211ai_1 _20453_ (.A1(_02054_),
    .A2(_02131_),
    .B1(_10513_),
    .C1(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__a21o_1 _20454_ (.A1(_10513_),
    .A2(_10515_),
    .B1(_10509_),
    .X(_10517_));
 sky130_fd_sc_hd__o22ai_4 _20455_ (.A1(_02054_),
    .A2(_02131_),
    .B1(_10512_),
    .B2(_10514_),
    .Y(_10518_));
 sky130_fd_sc_hd__nand4_2 _20456_ (.A(_10515_),
    .B(net18),
    .C(net45),
    .D(_10513_),
    .Y(_10519_));
 sky130_fd_sc_hd__nand2_1 _20457_ (.A(_10518_),
    .B(_10519_),
    .Y(_10520_));
 sky130_fd_sc_hd__and3_1 _20458_ (.A(_10518_),
    .B(_10519_),
    .C(_10507_),
    .X(_10522_));
 sky130_fd_sc_hd__nand3_2 _20459_ (.A(_10518_),
    .B(_10519_),
    .C(_10507_),
    .Y(_10523_));
 sky130_fd_sc_hd__a21oi_1 _20460_ (.A1(_10518_),
    .A2(_10519_),
    .B1(_10507_),
    .Y(_10524_));
 sky130_fd_sc_hd__nand3_2 _20461_ (.A(_10508_),
    .B(_10516_),
    .C(_10517_),
    .Y(_10525_));
 sky130_fd_sc_hd__a21oi_4 _20462_ (.A1(_10523_),
    .A2(_10525_),
    .B1(_10506_),
    .Y(_10526_));
 sky130_fd_sc_hd__and3_2 _20463_ (.A(_10525_),
    .B(_10506_),
    .C(_10523_),
    .X(_10527_));
 sky130_fd_sc_hd__a21oi_2 _20464_ (.A1(_10520_),
    .A2(_10508_),
    .B1(_10506_),
    .Y(_10528_));
 sky130_fd_sc_hd__and4_2 _20465_ (.A(_10504_),
    .B(_10505_),
    .C(_10523_),
    .D(_10525_),
    .X(_10529_));
 sky130_fd_sc_hd__o2bb2a_2 _20466_ (.A1_N(_10504_),
    .A2_N(_10505_),
    .B1(_10522_),
    .B2(_10524_),
    .X(_10530_));
 sky130_fd_sc_hd__a21o_1 _20467_ (.A1(_10523_),
    .A2(_10528_),
    .B1(_10530_),
    .X(_10531_));
 sky130_fd_sc_hd__nand2_2 _20468_ (.A(_10202_),
    .B(_10208_),
    .Y(_10533_));
 sky130_fd_sc_hd__o22a_1 _20469_ (.A1(_02010_),
    .A2(_02163_),
    .B1(_09925_),
    .B2(_10191_),
    .X(_10534_));
 sky130_fd_sc_hd__and3_1 _20470_ (.A(_10196_),
    .B(net20),
    .C(net41),
    .X(_10535_));
 sky130_fd_sc_hd__a31o_1 _20471_ (.A1(_10196_),
    .A2(net20),
    .A3(net41),
    .B1(_10193_),
    .X(_10536_));
 sky130_fd_sc_hd__o32a_2 _20472_ (.A1(_02010_),
    .A2(_02163_),
    .A3(_10195_),
    .B1(_10190_),
    .B2(_09922_),
    .X(_10537_));
 sky130_fd_sc_hd__a21oi_1 _20473_ (.A1(net38),
    .A2(net24),
    .B1(_10118_),
    .Y(_10538_));
 sky130_fd_sc_hd__o2111a_1 _20474_ (.A1(net36),
    .A2(net37),
    .B1(net38),
    .C1(net24),
    .D1(net25),
    .X(_10539_));
 sky130_fd_sc_hd__o21a_1 _20475_ (.A1(_10114_),
    .A2(_10116_),
    .B1(_10119_),
    .X(_10540_));
 sky130_fd_sc_hd__and2_1 _20476_ (.A(net41),
    .B(net21),
    .X(_10541_));
 sky130_fd_sc_hd__nand2_2 _20477_ (.A(net40),
    .B(net24),
    .Y(_10542_));
 sky130_fd_sc_hd__and4_1 _20478_ (.A(net39),
    .B(net40),
    .C(net22),
    .D(net24),
    .X(_10544_));
 sky130_fd_sc_hd__nand4_1 _20479_ (.A(net39),
    .B(net40),
    .C(net22),
    .D(net24),
    .Y(_10545_));
 sky130_fd_sc_hd__a22oi_4 _20480_ (.A1(net40),
    .A2(net22),
    .B1(net24),
    .B2(net39),
    .Y(_10546_));
 sky130_fd_sc_hd__a22o_2 _20481_ (.A1(net40),
    .A2(net22),
    .B1(net24),
    .B2(net39),
    .X(_10547_));
 sky130_fd_sc_hd__o221ai_4 _20482_ (.A1(_02010_),
    .A2(_02185_),
    .B1(_10191_),
    .B2(_10542_),
    .C1(_10547_),
    .Y(_10548_));
 sky130_fd_sc_hd__o21ai_1 _20483_ (.A1(_10544_),
    .A2(_10546_),
    .B1(_10541_),
    .Y(_10549_));
 sky130_fd_sc_hd__a2bb2oi_1 _20484_ (.A1_N(_02010_),
    .A2_N(_02185_),
    .B1(_10545_),
    .B2(_10547_),
    .Y(_10550_));
 sky130_fd_sc_hd__o2bb2ai_2 _20485_ (.A1_N(_10545_),
    .A2_N(_10547_),
    .B1(_02010_),
    .B2(_02185_),
    .Y(_10551_));
 sky130_fd_sc_hd__o211a_1 _20486_ (.A1(_10191_),
    .A2(_10542_),
    .B1(_10541_),
    .C1(_10547_),
    .X(_10552_));
 sky130_fd_sc_hd__o2111ai_4 _20487_ (.A1(_10191_),
    .A2(_10542_),
    .B1(net41),
    .C1(net21),
    .D1(_10547_),
    .Y(_10553_));
 sky130_fd_sc_hd__o211a_1 _20488_ (.A1(_10118_),
    .A2(_10539_),
    .B1(_10551_),
    .C1(_10553_),
    .X(_10555_));
 sky130_fd_sc_hd__o211ai_4 _20489_ (.A1(_10118_),
    .A2(_10539_),
    .B1(_10551_),
    .C1(_10553_),
    .Y(_10556_));
 sky130_fd_sc_hd__o22a_1 _20490_ (.A1(_10116_),
    .A2(_10538_),
    .B1(_10550_),
    .B2(_10552_),
    .X(_10557_));
 sky130_fd_sc_hd__o22ai_2 _20491_ (.A1(_10116_),
    .A2(_10538_),
    .B1(_10550_),
    .B2(_10552_),
    .Y(_10558_));
 sky130_fd_sc_hd__a31oi_4 _20492_ (.A1(_10540_),
    .A2(_10548_),
    .A3(_10549_),
    .B1(_10537_),
    .Y(_10559_));
 sky130_fd_sc_hd__o211a_1 _20493_ (.A1(_10193_),
    .A2(_10535_),
    .B1(_10556_),
    .C1(_10558_),
    .X(_10560_));
 sky130_fd_sc_hd__nand2_2 _20494_ (.A(_10559_),
    .B(_10556_),
    .Y(_10561_));
 sky130_fd_sc_hd__a2bb2oi_2 _20495_ (.A1_N(_10195_),
    .A2_N(_10534_),
    .B1(_10556_),
    .B2(_10558_),
    .Y(_10562_));
 sky130_fd_sc_hd__o22ai_4 _20496_ (.A1(_10195_),
    .A2(_10534_),
    .B1(_10555_),
    .B2(_10557_),
    .Y(_10563_));
 sky130_fd_sc_hd__a221oi_4 _20497_ (.A1(_10559_),
    .A2(_10556_),
    .B1(_10208_),
    .B2(_10202_),
    .C1(_10562_),
    .Y(_10564_));
 sky130_fd_sc_hd__nand3_4 _20498_ (.A(_10533_),
    .B(_10561_),
    .C(_10563_),
    .Y(_10566_));
 sky130_fd_sc_hd__a21oi_4 _20499_ (.A1(_10561_),
    .A2(_10563_),
    .B1(_10533_),
    .Y(_10567_));
 sky130_fd_sc_hd__o211ai_4 _20500_ (.A1(_10560_),
    .A2(_10562_),
    .B1(_10202_),
    .C1(_10208_),
    .Y(_10568_));
 sky130_fd_sc_hd__o22ai_4 _20501_ (.A1(_10526_),
    .A2(_10527_),
    .B1(_10564_),
    .B2(_10567_),
    .Y(_10569_));
 sky130_fd_sc_hd__o211ai_4 _20502_ (.A1(_10529_),
    .A2(_10530_),
    .B1(_10566_),
    .C1(_10568_),
    .Y(_10570_));
 sky130_fd_sc_hd__o211ai_4 _20503_ (.A1(_10526_),
    .A2(_10527_),
    .B1(_10566_),
    .C1(_10568_),
    .Y(_10571_));
 sky130_fd_sc_hd__o22ai_4 _20504_ (.A1(_10529_),
    .A2(_10530_),
    .B1(_10564_),
    .B2(_10567_),
    .Y(_10572_));
 sky130_fd_sc_hd__and3_1 _20505_ (.A(_10569_),
    .B(_10570_),
    .C(_10497_),
    .X(_10573_));
 sky130_fd_sc_hd__nand3_4 _20506_ (.A(_10569_),
    .B(_10570_),
    .C(_10497_),
    .Y(_10574_));
 sky130_fd_sc_hd__and3_1 _20507_ (.A(_10498_),
    .B(_10571_),
    .C(_10572_),
    .X(_10575_));
 sky130_fd_sc_hd__o211ai_4 _20508_ (.A1(_10132_),
    .A2(_10136_),
    .B1(_10571_),
    .C1(_10572_),
    .Y(_10577_));
 sky130_fd_sc_hd__and3_1 _20509_ (.A(_10184_),
    .B(_10186_),
    .C(_10213_),
    .X(_10578_));
 sky130_fd_sc_hd__a21oi_2 _20510_ (.A1(_10184_),
    .A2(_10186_),
    .B1(_10209_),
    .Y(_10579_));
 sky130_fd_sc_hd__o31a_1 _20511_ (.A1(_10183_),
    .A2(_10185_),
    .A3(_10212_),
    .B1(_10210_),
    .X(_10580_));
 sky130_fd_sc_hd__a31o_1 _20512_ (.A1(_10184_),
    .A2(_10186_),
    .A3(_10213_),
    .B1(_10209_),
    .X(_10581_));
 sky130_fd_sc_hd__o2bb2ai_4 _20513_ (.A1_N(_10574_),
    .A2_N(_10577_),
    .B1(_10578_),
    .B2(_10209_),
    .Y(_10582_));
 sky130_fd_sc_hd__a31oi_4 _20514_ (.A1(_10569_),
    .A2(_10570_),
    .A3(_10497_),
    .B1(_10581_),
    .Y(_10583_));
 sky130_fd_sc_hd__o211ai_4 _20515_ (.A1(_10212_),
    .A2(_10579_),
    .B1(_10577_),
    .C1(_10574_),
    .Y(_10584_));
 sky130_fd_sc_hd__o211ai_2 _20516_ (.A1(_10209_),
    .A2(_10578_),
    .B1(_10577_),
    .C1(_10574_),
    .Y(_10585_));
 sky130_fd_sc_hd__o2bb2ai_1 _20517_ (.A1_N(_10574_),
    .A2_N(_10577_),
    .B1(_10579_),
    .B2(_10212_),
    .Y(_10586_));
 sky130_fd_sc_hd__a22oi_4 _20518_ (.A1(_10493_),
    .A2(_10495_),
    .B1(_10582_),
    .B2(_10584_),
    .Y(_10588_));
 sky130_fd_sc_hd__a22o_1 _20519_ (.A1(_10493_),
    .A2(_10495_),
    .B1(_10582_),
    .B2(_10584_),
    .X(_10589_));
 sky130_fd_sc_hd__a211oi_1 _20520_ (.A1(_10583_),
    .A2(_10577_),
    .B1(_10494_),
    .C1(_10492_),
    .Y(_10590_));
 sky130_fd_sc_hd__a21oi_2 _20521_ (.A1(_10585_),
    .A2(_10586_),
    .B1(_10496_),
    .Y(_10591_));
 sky130_fd_sc_hd__a21o_1 _20522_ (.A1(_10585_),
    .A2(_10586_),
    .B1(_10496_),
    .X(_10592_));
 sky130_fd_sc_hd__a221oi_2 _20523_ (.A1(_10590_),
    .A2(_10582_),
    .B1(_10233_),
    .B2(_10144_),
    .C1(_10588_),
    .Y(_10593_));
 sky130_fd_sc_hd__nand3_2 _20524_ (.A(_10462_),
    .B(_10589_),
    .C(_10592_),
    .Y(_10594_));
 sky130_fd_sc_hd__o21a_1 _20525_ (.A1(_10588_),
    .A2(_10591_),
    .B1(_10461_),
    .X(_10595_));
 sky130_fd_sc_hd__o21ai_2 _20526_ (.A1(_10588_),
    .A2(_10591_),
    .B1(_10461_),
    .Y(_10596_));
 sky130_fd_sc_hd__a21o_1 _20527_ (.A1(_10594_),
    .A2(_10596_),
    .B1(_10460_),
    .X(_10597_));
 sky130_fd_sc_hd__o211ai_2 _20528_ (.A1(_10456_),
    .A2(_10459_),
    .B1(_10594_),
    .C1(_10596_),
    .Y(_10599_));
 sky130_fd_sc_hd__o22ai_2 _20529_ (.A1(_10456_),
    .A2(_10459_),
    .B1(_10593_),
    .B2(_10595_),
    .Y(_10600_));
 sky130_fd_sc_hd__o2111ai_2 _20530_ (.A1(_10458_),
    .A2(_10451_),
    .B1(_10457_),
    .C1(_10594_),
    .D1(_10596_),
    .Y(_10601_));
 sky130_fd_sc_hd__a31oi_2 _20531_ (.A1(_10240_),
    .A2(_10325_),
    .A3(_10327_),
    .B1(_10237_),
    .Y(_10602_));
 sky130_fd_sc_hd__a31oi_2 _20532_ (.A1(_10238_),
    .A2(_10329_),
    .A3(_10331_),
    .B1(_10239_),
    .Y(_10603_));
 sky130_fd_sc_hd__nand3_2 _20533_ (.A(_10597_),
    .B(_10599_),
    .C(_10603_),
    .Y(_10604_));
 sky130_fd_sc_hd__inv_2 _20534_ (.A(_10604_),
    .Y(_10605_));
 sky130_fd_sc_hd__and3_1 _20535_ (.A(_10600_),
    .B(_10602_),
    .C(_10601_),
    .X(_10606_));
 sky130_fd_sc_hd__nand3_2 _20536_ (.A(_10600_),
    .B(_10602_),
    .C(_10601_),
    .Y(_10607_));
 sky130_fd_sc_hd__a31o_1 _20537_ (.A1(_10025_),
    .A2(_10057_),
    .A3(_10318_),
    .B1(_10319_),
    .X(_10608_));
 sky130_fd_sc_hd__inv_2 _20538_ (.A(_10608_),
    .Y(_10610_));
 sky130_fd_sc_hd__a21o_1 _20539_ (.A1(_10604_),
    .A2(_10607_),
    .B1(_10610_),
    .X(_10611_));
 sky130_fd_sc_hd__a31oi_2 _20540_ (.A1(_10597_),
    .A2(_10599_),
    .A3(_10603_),
    .B1(_10608_),
    .Y(_10612_));
 sky130_fd_sc_hd__o211ai_2 _20541_ (.A1(_10317_),
    .A2(_10330_),
    .B1(_10604_),
    .C1(_10607_),
    .Y(_10613_));
 sky130_fd_sc_hd__a22o_1 _20542_ (.A1(_10318_),
    .A2(_10331_),
    .B1(_10604_),
    .B2(_10607_),
    .X(_10614_));
 sky130_fd_sc_hd__o2111ai_1 _20543_ (.A1(_10322_),
    .A2(_10319_),
    .B1(_10318_),
    .C1(_10607_),
    .D1(_10604_),
    .Y(_10615_));
 sky130_fd_sc_hd__nand2_1 _20544_ (.A(_10611_),
    .B(_10613_),
    .Y(_10616_));
 sky130_fd_sc_hd__nand3_2 _20545_ (.A(_10371_),
    .B(_10614_),
    .C(_10615_),
    .Y(_10617_));
 sky130_fd_sc_hd__and3_1 _20546_ (.A(_10611_),
    .B(_10613_),
    .C(_10370_),
    .X(_10618_));
 sky130_fd_sc_hd__nand3_2 _20547_ (.A(_10611_),
    .B(_10613_),
    .C(_10370_),
    .Y(_10619_));
 sky130_fd_sc_hd__nor2_1 _20548_ (.A(_10041_),
    .B(_10304_),
    .Y(_10621_));
 sky130_fd_sc_hd__a21o_1 _20549_ (.A1(_10303_),
    .A2(_10041_),
    .B1(_10304_),
    .X(_10622_));
 sky130_fd_sc_hd__a21oi_2 _20550_ (.A1(_10617_),
    .A2(_10619_),
    .B1(_10622_),
    .Y(_10623_));
 sky130_fd_sc_hd__o2bb2ai_1 _20551_ (.A1_N(_10617_),
    .A2_N(_10619_),
    .B1(_10621_),
    .B2(_10301_),
    .Y(_10624_));
 sky130_fd_sc_hd__and3_1 _20552_ (.A(_10617_),
    .B(_10619_),
    .C(_10622_),
    .X(_10625_));
 sky130_fd_sc_hd__nand3_2 _20553_ (.A(_10617_),
    .B(_10619_),
    .C(_10622_),
    .Y(_10626_));
 sky130_fd_sc_hd__o21ai_1 _20554_ (.A1(_10109_),
    .A2(_10344_),
    .B1(_10353_),
    .Y(_10627_));
 sky130_fd_sc_hd__o21a_1 _20555_ (.A1(_10109_),
    .A2(_10344_),
    .B1(_10353_),
    .X(_10628_));
 sky130_fd_sc_hd__a21oi_1 _20556_ (.A1(_10624_),
    .A2(_10626_),
    .B1(_10627_),
    .Y(_10629_));
 sky130_fd_sc_hd__o21ai_2 _20557_ (.A1(_10623_),
    .A2(_10625_),
    .B1(_10628_),
    .Y(_10630_));
 sky130_fd_sc_hd__o21ai_2 _20558_ (.A1(_10347_),
    .A2(_10352_),
    .B1(_10626_),
    .Y(_10632_));
 sky130_fd_sc_hd__nand3_1 _20559_ (.A(_10624_),
    .B(_10627_),
    .C(_10626_),
    .Y(_10633_));
 sky130_fd_sc_hd__o21ai_1 _20560_ (.A1(_10623_),
    .A2(_10632_),
    .B1(_10630_),
    .Y(_10634_));
 sky130_fd_sc_hd__a21oi_1 _20561_ (.A1(_10360_),
    .A2(_10369_),
    .B1(_10634_),
    .Y(_10635_));
 sky130_fd_sc_hd__and3_1 _20562_ (.A(_10360_),
    .B(_10369_),
    .C(_10634_),
    .X(_10636_));
 sky130_fd_sc_hd__nor2_1 _20563_ (.A(_10635_),
    .B(_10636_),
    .Y(net104));
 sky130_fd_sc_hd__and3_1 _20564_ (.A(_10277_),
    .B(_10315_),
    .C(_10452_),
    .X(_10637_));
 sky130_fd_sc_hd__a31o_1 _20565_ (.A1(_10277_),
    .A2(_10315_),
    .A3(_10452_),
    .B1(_10450_),
    .X(_10638_));
 sky130_fd_sc_hd__o211ai_1 _20566_ (.A1(_10458_),
    .A2(_10451_),
    .B1(_10457_),
    .C1(_10596_),
    .Y(_10639_));
 sky130_fd_sc_hd__a21oi_1 _20567_ (.A1(_10460_),
    .A2(_10594_),
    .B1(_10595_),
    .Y(_10640_));
 sky130_fd_sc_hd__o21ai_2 _20568_ (.A1(_10374_),
    .A2(_10395_),
    .B1(_10398_),
    .Y(_10642_));
 sky130_fd_sc_hd__o21a_1 _20569_ (.A1(_10374_),
    .A2(_10395_),
    .B1(_10398_),
    .X(_10643_));
 sky130_fd_sc_hd__a21boi_2 _20570_ (.A1(_10387_),
    .A2(_10391_),
    .B1_N(_10388_),
    .Y(_10644_));
 sky130_fd_sc_hd__a31o_1 _20571_ (.A1(_10503_),
    .A2(net48),
    .A3(net15),
    .B1(_10501_),
    .X(_10645_));
 sky130_fd_sc_hd__a31oi_4 _20572_ (.A1(_10503_),
    .A2(net48),
    .A3(net15),
    .B1(_10501_),
    .Y(_10646_));
 sky130_fd_sc_hd__nand2_1 _20573_ (.A(net13),
    .B(net51),
    .Y(_10647_));
 sky130_fd_sc_hd__nand2_1 _20574_ (.A(net15),
    .B(net49),
    .Y(_10648_));
 sky130_fd_sc_hd__a22oi_1 _20575_ (.A1(net15),
    .A2(net49),
    .B1(net50),
    .B2(net14),
    .Y(_10649_));
 sky130_fd_sc_hd__a22o_2 _20576_ (.A1(net15),
    .A2(net49),
    .B1(net50),
    .B2(net14),
    .X(_10650_));
 sky130_fd_sc_hd__and4_1 _20577_ (.A(net14),
    .B(net15),
    .C(net49),
    .D(net50),
    .X(_10651_));
 sky130_fd_sc_hd__nand4_4 _20578_ (.A(net14),
    .B(net15),
    .C(net49),
    .D(net50),
    .Y(_10653_));
 sky130_fd_sc_hd__o211ai_4 _20579_ (.A1(_02043_),
    .A2(_02152_),
    .B1(_10650_),
    .C1(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__a21o_1 _20580_ (.A1(_10650_),
    .A2(_10653_),
    .B1(_10647_),
    .X(_10655_));
 sky130_fd_sc_hd__a22o_1 _20581_ (.A1(net13),
    .A2(net51),
    .B1(_10650_),
    .B2(_10653_),
    .X(_10656_));
 sky130_fd_sc_hd__nand4_1 _20582_ (.A(_10650_),
    .B(_10653_),
    .C(net13),
    .D(net51),
    .Y(_10657_));
 sky130_fd_sc_hd__nand3_4 _20583_ (.A(_10646_),
    .B(_10654_),
    .C(_10655_),
    .Y(_10658_));
 sky130_fd_sc_hd__inv_2 _20584_ (.A(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__a21oi_4 _20585_ (.A1(_10654_),
    .A2(_10655_),
    .B1(_10646_),
    .Y(_10660_));
 sky130_fd_sc_hd__nand3_2 _20586_ (.A(_10645_),
    .B(_10656_),
    .C(_10657_),
    .Y(_10661_));
 sky130_fd_sc_hd__o21a_1 _20587_ (.A1(_02032_),
    .A2(_02152_),
    .B1(_10382_),
    .X(_10662_));
 sky130_fd_sc_hd__and3_1 _20588_ (.A(_10380_),
    .B(net51),
    .C(net11),
    .X(_10664_));
 sky130_fd_sc_hd__o2bb2ai_2 _20589_ (.A1_N(_10658_),
    .A2_N(_10661_),
    .B1(_10662_),
    .B2(_10379_),
    .Y(_10665_));
 sky130_fd_sc_hd__o21a_1 _20590_ (.A1(_10381_),
    .A2(_10664_),
    .B1(_10658_),
    .X(_10666_));
 sky130_fd_sc_hd__o21ai_2 _20591_ (.A1(_10381_),
    .A2(_10664_),
    .B1(_10658_),
    .Y(_10667_));
 sky130_fd_sc_hd__o2111ai_4 _20592_ (.A1(_10377_),
    .A2(_10379_),
    .B1(_10382_),
    .C1(_10658_),
    .D1(_10661_),
    .Y(_10668_));
 sky130_fd_sc_hd__o2bb2ai_2 _20593_ (.A1_N(_10658_),
    .A2_N(_10661_),
    .B1(_10664_),
    .B2(_10381_),
    .Y(_10669_));
 sky130_fd_sc_hd__o21a_1 _20594_ (.A1(_10506_),
    .A2(_10524_),
    .B1(_10523_),
    .X(_10670_));
 sky130_fd_sc_hd__nand3_1 _20595_ (.A(_10670_),
    .B(_10669_),
    .C(_10668_),
    .Y(_10671_));
 sky130_fd_sc_hd__o221a_1 _20596_ (.A1(_10660_),
    .A2(_10667_),
    .B1(_10522_),
    .B2(_10528_),
    .C1(_10665_),
    .X(_10672_));
 sky130_fd_sc_hd__o221ai_4 _20597_ (.A1(_10660_),
    .A2(_10667_),
    .B1(_10522_),
    .B2(_10528_),
    .C1(_10665_),
    .Y(_10673_));
 sky130_fd_sc_hd__a22o_1 _20598_ (.A1(_10388_),
    .A2(_10393_),
    .B1(_10671_),
    .B2(_10673_),
    .X(_10675_));
 sky130_fd_sc_hd__nand4_2 _20599_ (.A(_10388_),
    .B(_10393_),
    .C(_10671_),
    .D(_10673_),
    .Y(_10676_));
 sky130_fd_sc_hd__a21bo_1 _20600_ (.A1(_10671_),
    .A2(_10673_),
    .B1_N(_10644_),
    .X(_10677_));
 sky130_fd_sc_hd__a31oi_4 _20601_ (.A1(_10670_),
    .A2(_10669_),
    .A3(_10668_),
    .B1(_10644_),
    .Y(_10678_));
 sky130_fd_sc_hd__nand2_1 _20602_ (.A(_10678_),
    .B(_10673_),
    .Y(_10679_));
 sky130_fd_sc_hd__nand3_4 _20603_ (.A(_10643_),
    .B(_10675_),
    .C(_10676_),
    .Y(_10680_));
 sky130_fd_sc_hd__inv_2 _20604_ (.A(_10680_),
    .Y(_10681_));
 sky130_fd_sc_hd__and3_2 _20605_ (.A(_10677_),
    .B(_10679_),
    .C(_10642_),
    .X(_10682_));
 sky130_fd_sc_hd__nand3_4 _20606_ (.A(_10677_),
    .B(_10679_),
    .C(_10642_),
    .Y(_10683_));
 sky130_fd_sc_hd__nand2_1 _20607_ (.A(_10421_),
    .B(_10430_),
    .Y(_10684_));
 sky130_fd_sc_hd__a22o_1 _20608_ (.A1(net8),
    .A2(net56),
    .B1(_01977_),
    .B2(net57),
    .X(_10686_));
 sky130_fd_sc_hd__nand2_1 _20609_ (.A(_01977_),
    .B(net8),
    .Y(_10687_));
 sky130_fd_sc_hd__and3_1 _20610_ (.A(_01977_),
    .B(net8),
    .C(net56),
    .X(_10688_));
 sky130_fd_sc_hd__or4_2 _20611_ (.A(net7),
    .B(_01988_),
    .C(_02229_),
    .D(_02240_),
    .X(_10689_));
 sky130_fd_sc_hd__o31a_1 _20612_ (.A1(_02229_),
    .A2(_02240_),
    .A3(_10687_),
    .B1(_10686_),
    .X(_10690_));
 sky130_fd_sc_hd__nor2_1 _20613_ (.A(_10410_),
    .B(_10412_),
    .Y(_10691_));
 sky130_fd_sc_hd__o32a_1 _20614_ (.A1(_01999_),
    .A2(_02174_),
    .A3(_10414_),
    .B1(_10412_),
    .B2(_10410_),
    .X(_10692_));
 sky130_fd_sc_hd__nand2_1 _20615_ (.A(net9),
    .B(net54),
    .Y(_10693_));
 sky130_fd_sc_hd__nand2_2 _20616_ (.A(net11),
    .B(net52),
    .Y(_10694_));
 sky130_fd_sc_hd__a22oi_2 _20617_ (.A1(net11),
    .A2(net52),
    .B1(net53),
    .B2(net10),
    .Y(_10695_));
 sky130_fd_sc_hd__a22o_1 _20618_ (.A1(net11),
    .A2(net52),
    .B1(net53),
    .B2(net10),
    .X(_10697_));
 sky130_fd_sc_hd__nand2_1 _20619_ (.A(net11),
    .B(net53),
    .Y(_10698_));
 sky130_fd_sc_hd__and4_1 _20620_ (.A(net10),
    .B(net11),
    .C(net52),
    .D(net53),
    .X(_10699_));
 sky130_fd_sc_hd__nand4_2 _20621_ (.A(net10),
    .B(net11),
    .C(net52),
    .D(net53),
    .Y(_10700_));
 sky130_fd_sc_hd__o211ai_1 _20622_ (.A1(_01999_),
    .A2(_02207_),
    .B1(_10697_),
    .C1(_10700_),
    .Y(_10701_));
 sky130_fd_sc_hd__a21o_1 _20623_ (.A1(_10697_),
    .A2(_10700_),
    .B1(_10693_),
    .X(_10702_));
 sky130_fd_sc_hd__o21ai_1 _20624_ (.A1(_10695_),
    .A2(_10699_),
    .B1(_10693_),
    .Y(_10703_));
 sky130_fd_sc_hd__and4_1 _20625_ (.A(_10697_),
    .B(_10700_),
    .C(net9),
    .D(net54),
    .X(_10704_));
 sky130_fd_sc_hd__nand4_1 _20626_ (.A(_10697_),
    .B(_10700_),
    .C(net9),
    .D(net54),
    .Y(_10705_));
 sky130_fd_sc_hd__nand3_2 _20627_ (.A(_10692_),
    .B(_10701_),
    .C(_10702_),
    .Y(_10706_));
 sky130_fd_sc_hd__o21ai_2 _20628_ (.A1(_10415_),
    .A2(_10691_),
    .B1(_10703_),
    .Y(_10708_));
 sky130_fd_sc_hd__o211ai_2 _20629_ (.A1(_10415_),
    .A2(_10691_),
    .B1(_10703_),
    .C1(_10705_),
    .Y(_10709_));
 sky130_fd_sc_hd__a21oi_1 _20630_ (.A1(_10706_),
    .A2(_10709_),
    .B1(_10690_),
    .Y(_10710_));
 sky130_fd_sc_hd__a22o_1 _20631_ (.A1(_10686_),
    .A2(_10689_),
    .B1(_10706_),
    .B2(_10709_),
    .X(_10711_));
 sky130_fd_sc_hd__and3_1 _20632_ (.A(_10706_),
    .B(_10709_),
    .C(_10690_),
    .X(_10712_));
 sky130_fd_sc_hd__o2111ai_4 _20633_ (.A1(_10704_),
    .A2(_10708_),
    .B1(_10706_),
    .C1(_10686_),
    .D1(_10689_),
    .Y(_10713_));
 sky130_fd_sc_hd__o211ai_4 _20634_ (.A1(_10710_),
    .A2(_10712_),
    .B1(_10421_),
    .C1(_10430_),
    .Y(_10714_));
 sky130_fd_sc_hd__nand3_2 _20635_ (.A(_10684_),
    .B(_10711_),
    .C(_10713_),
    .Y(_10715_));
 sky130_fd_sc_hd__nand2_1 _20636_ (.A(_10714_),
    .B(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__o31a_1 _20637_ (.A1(_01977_),
    .A2(_02229_),
    .A3(_10424_),
    .B1(_10716_),
    .X(_10717_));
 sky130_fd_sc_hd__and3_1 _20638_ (.A(_10714_),
    .B(_10715_),
    .C(_10425_),
    .X(_10719_));
 sky130_fd_sc_hd__o311a_1 _20639_ (.A1(_01977_),
    .A2(_02229_),
    .A3(_10424_),
    .B1(_10714_),
    .C1(_10715_),
    .X(_10720_));
 sky130_fd_sc_hd__a41o_1 _20640_ (.A1(_01966_),
    .A2(net7),
    .A3(net56),
    .A4(net57),
    .B1(_10716_),
    .X(_10721_));
 sky130_fd_sc_hd__a21oi_2 _20641_ (.A1(_10714_),
    .A2(_10715_),
    .B1(_10426_),
    .Y(_10722_));
 sky130_fd_sc_hd__a21o_1 _20642_ (.A1(_10714_),
    .A2(_10715_),
    .B1(_10426_),
    .X(_10723_));
 sky130_fd_sc_hd__o2bb2ai_2 _20643_ (.A1_N(_10680_),
    .A2_N(_10683_),
    .B1(_10717_),
    .B2(_10719_),
    .Y(_10724_));
 sky130_fd_sc_hd__o21a_1 _20644_ (.A1(_10720_),
    .A2(_10722_),
    .B1(_10680_),
    .X(_10725_));
 sky130_fd_sc_hd__o211ai_2 _20645_ (.A1(_10720_),
    .A2(_10722_),
    .B1(_10680_),
    .C1(_10683_),
    .Y(_10726_));
 sky130_fd_sc_hd__nand4_2 _20646_ (.A(_10680_),
    .B(_10683_),
    .C(_10721_),
    .D(_10723_),
    .Y(_10727_));
 sky130_fd_sc_hd__o2bb2ai_1 _20647_ (.A1_N(_10680_),
    .A2_N(_10683_),
    .B1(_10720_),
    .B2(_10722_),
    .Y(_10728_));
 sky130_fd_sc_hd__a31oi_2 _20648_ (.A1(_10498_),
    .A2(_10571_),
    .A3(_10572_),
    .B1(_10580_),
    .Y(_10730_));
 sky130_fd_sc_hd__o211ai_4 _20649_ (.A1(_10573_),
    .A2(_10730_),
    .B1(_10728_),
    .C1(_10727_),
    .Y(_10731_));
 sky130_fd_sc_hd__inv_2 _20650_ (.A(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__o211ai_4 _20651_ (.A1(_10575_),
    .A2(_10583_),
    .B1(_10724_),
    .C1(_10726_),
    .Y(_10733_));
 sky130_fd_sc_hd__o21a_1 _20652_ (.A1(_10436_),
    .A2(_10439_),
    .B1(_10406_),
    .X(_10734_));
 sky130_fd_sc_hd__a32o_1 _20653_ (.A1(_10372_),
    .A2(_10402_),
    .A3(_10403_),
    .B1(_10406_),
    .B2(_10442_),
    .X(_10735_));
 sky130_fd_sc_hd__nand3b_1 _20654_ (.A_N(_10735_),
    .B(_10733_),
    .C(_10731_),
    .Y(_10736_));
 sky130_fd_sc_hd__o2bb2ai_2 _20655_ (.A1_N(_10731_),
    .A2_N(_10733_),
    .B1(_10734_),
    .B2(_10405_),
    .Y(_10737_));
 sky130_fd_sc_hd__a21oi_1 _20656_ (.A1(_10731_),
    .A2(_10733_),
    .B1(_10735_),
    .Y(_10738_));
 sky130_fd_sc_hd__and3_1 _20657_ (.A(_10731_),
    .B(_10733_),
    .C(_10735_),
    .X(_10739_));
 sky130_fd_sc_hd__o2111ai_1 _20658_ (.A1(_10442_),
    .A2(_10405_),
    .B1(_10406_),
    .C1(_10731_),
    .D1(_10733_),
    .Y(_10741_));
 sky130_fd_sc_hd__a31oi_2 _20659_ (.A1(_10493_),
    .A2(_10582_),
    .A3(_10584_),
    .B1(_10494_),
    .Y(_10742_));
 sky130_fd_sc_hd__a31o_1 _20660_ (.A1(_10493_),
    .A2(_10582_),
    .A3(_10584_),
    .B1(_10494_),
    .X(_10743_));
 sky130_fd_sc_hd__o2bb2ai_2 _20661_ (.A1_N(_08963_),
    .A2_N(_08006_),
    .B1(_10485_),
    .B2(_10483_),
    .Y(_10744_));
 sky130_fd_sc_hd__a31o_2 _20662_ (.A1(_10472_),
    .A2(_09845_),
    .A3(_10470_),
    .B1(_09657_),
    .X(_10745_));
 sky130_fd_sc_hd__a21oi_4 _20663_ (.A1(_10479_),
    .A2(_10482_),
    .B1(_10745_),
    .Y(_10746_));
 sky130_fd_sc_hd__a21o_4 _20664_ (.A1(_10479_),
    .A2(_10482_),
    .B1(_10745_),
    .X(_10747_));
 sky130_fd_sc_hd__o221a_4 _20665_ (.A1(_09657_),
    .A2(_10476_),
    .B1(_10473_),
    .B2(_10480_),
    .C1(_10479_),
    .X(_10748_));
 sky130_fd_sc_hd__o211ai_4 _20666_ (.A1(_09657_),
    .A2(_10476_),
    .B1(_10479_),
    .C1(_10482_),
    .Y(_10749_));
 sky130_fd_sc_hd__nor2_8 _20667_ (.A(_10746_),
    .B(_10748_),
    .Y(_10750_));
 sky130_fd_sc_hd__nand2_4 _20668_ (.A(_10747_),
    .B(_10749_),
    .Y(_10752_));
 sky130_fd_sc_hd__o21ai_2 _20669_ (.A1(_10746_),
    .A2(_10748_),
    .B1(_09388_),
    .Y(_10753_));
 sky130_fd_sc_hd__nand4_4 _20670_ (.A(_09384_),
    .B(_09386_),
    .C(_10747_),
    .D(_10749_),
    .Y(_10754_));
 sky130_fd_sc_hd__and4_1 _20671_ (.A(_09384_),
    .B(_10744_),
    .C(_10753_),
    .D(_10754_),
    .X(_10755_));
 sky130_fd_sc_hd__nand4_4 _20672_ (.A(_09384_),
    .B(_10744_),
    .C(_10753_),
    .D(_10754_),
    .Y(_10756_));
 sky130_fd_sc_hd__a22oi_2 _20673_ (.A1(_09384_),
    .A2(_10744_),
    .B1(_10753_),
    .B2(_10754_),
    .Y(_10757_));
 sky130_fd_sc_hd__a22o_1 _20674_ (.A1(_09384_),
    .A2(_10744_),
    .B1(_10753_),
    .B2(_10754_),
    .X(_10758_));
 sky130_fd_sc_hd__o31a_1 _20675_ (.A1(_10526_),
    .A2(_10527_),
    .A3(_10564_),
    .B1(_10568_),
    .X(_10759_));
 sky130_fd_sc_hd__o31a_1 _20676_ (.A1(_09342_),
    .A2(_10473_),
    .A3(_10476_),
    .B1(_10484_),
    .X(_10760_));
 sky130_fd_sc_hd__o21a_1 _20677_ (.A1(_02054_),
    .A2(_02131_),
    .B1(_10513_),
    .X(_10761_));
 sky130_fd_sc_hd__nor2_1 _20678_ (.A(_10509_),
    .B(_10514_),
    .Y(_10763_));
 sky130_fd_sc_hd__a31o_1 _20679_ (.A1(_10515_),
    .A2(net18),
    .A3(net45),
    .B1(_10512_),
    .X(_10764_));
 sky130_fd_sc_hd__nand2_1 _20680_ (.A(net43),
    .B(net21),
    .Y(_10765_));
 sky130_fd_sc_hd__nand2_2 _20681_ (.A(net42),
    .B(net21),
    .Y(_10766_));
 sky130_fd_sc_hd__nand4_4 _20682_ (.A(net42),
    .B(net43),
    .C(net20),
    .D(net21),
    .Y(_10767_));
 sky130_fd_sc_hd__a22oi_2 _20683_ (.A1(net43),
    .A2(net20),
    .B1(net21),
    .B2(net42),
    .Y(_10768_));
 sky130_fd_sc_hd__a22o_1 _20684_ (.A1(net43),
    .A2(net20),
    .B1(net21),
    .B2(net42),
    .X(_10769_));
 sky130_fd_sc_hd__a22oi_2 _20685_ (.A1(net45),
    .A2(net19),
    .B1(_10767_),
    .B2(_10769_),
    .Y(_10770_));
 sky130_fd_sc_hd__o2bb2ai_2 _20686_ (.A1_N(_10767_),
    .A2_N(_10769_),
    .B1(_02054_),
    .B2(_02142_),
    .Y(_10771_));
 sky130_fd_sc_hd__o2111a_4 _20687_ (.A1(_10511_),
    .A2(_10765_),
    .B1(net45),
    .C1(net19),
    .D1(_10769_),
    .X(_10772_));
 sky130_fd_sc_hd__o22ai_4 _20688_ (.A1(_10514_),
    .A2(_10761_),
    .B1(_10770_),
    .B2(_10772_),
    .Y(_10774_));
 sky130_fd_sc_hd__o21ai_4 _20689_ (.A1(_10512_),
    .A2(_10763_),
    .B1(_10771_),
    .Y(_10775_));
 sky130_fd_sc_hd__nand3b_1 _20690_ (.A_N(_10772_),
    .B(_10764_),
    .C(_10771_),
    .Y(_10776_));
 sky130_fd_sc_hd__a22oi_4 _20691_ (.A1(net47),
    .A2(net17),
    .B1(net18),
    .B2(net46),
    .Y(_10777_));
 sky130_fd_sc_hd__a22o_1 _20692_ (.A1(net47),
    .A2(net17),
    .B1(net18),
    .B2(net46),
    .X(_10778_));
 sky130_fd_sc_hd__nand2_1 _20693_ (.A(net47),
    .B(net18),
    .Y(_10779_));
 sky130_fd_sc_hd__nand4_4 _20694_ (.A(net46),
    .B(net47),
    .C(net17),
    .D(net18),
    .Y(_10780_));
 sky130_fd_sc_hd__a22oi_4 _20695_ (.A1(net16),
    .A2(net48),
    .B1(_10778_),
    .B2(_10780_),
    .Y(_10781_));
 sky130_fd_sc_hd__a22o_1 _20696_ (.A1(net16),
    .A2(net48),
    .B1(_10778_),
    .B2(_10780_),
    .X(_10782_));
 sky130_fd_sc_hd__o2111a_1 _20697_ (.A1(_10500_),
    .A2(_10779_),
    .B1(net16),
    .C1(net48),
    .D1(_10778_),
    .X(_10783_));
 sky130_fd_sc_hd__or4b_2 _20698_ (.A(_02098_),
    .B(_02109_),
    .C(_10777_),
    .D_N(_10780_),
    .X(_10785_));
 sky130_fd_sc_hd__nor2_1 _20699_ (.A(_10781_),
    .B(_10783_),
    .Y(_10786_));
 sky130_fd_sc_hd__o221ai_4 _20700_ (.A1(_10781_),
    .A2(_10783_),
    .B1(_10772_),
    .B2(_10775_),
    .C1(_10774_),
    .Y(_10787_));
 sky130_fd_sc_hd__a21bo_1 _20701_ (.A1(_10774_),
    .A2(_10776_),
    .B1_N(_10786_),
    .X(_10788_));
 sky130_fd_sc_hd__o2111ai_4 _20702_ (.A1(_10772_),
    .A2(_10775_),
    .B1(_10782_),
    .C1(_10785_),
    .D1(_10774_),
    .Y(_10789_));
 sky130_fd_sc_hd__a22o_1 _20703_ (.A1(_10774_),
    .A2(_10776_),
    .B1(_10782_),
    .B2(_10785_),
    .X(_10790_));
 sky130_fd_sc_hd__a21oi_1 _20704_ (.A1(_10558_),
    .A2(_10536_),
    .B1(_10555_),
    .Y(_10791_));
 sky130_fd_sc_hd__o21ai_2 _20705_ (.A1(_10537_),
    .A2(_10557_),
    .B1(_10556_),
    .Y(_10792_));
 sky130_fd_sc_hd__o22a_1 _20706_ (.A1(_02010_),
    .A2(_02185_),
    .B1(_10191_),
    .B2(_10542_),
    .X(_10793_));
 sky130_fd_sc_hd__and3_1 _20707_ (.A(_10547_),
    .B(net21),
    .C(net41),
    .X(_10794_));
 sky130_fd_sc_hd__a31o_1 _20708_ (.A1(_10547_),
    .A2(net21),
    .A3(net41),
    .B1(_10544_),
    .X(_10796_));
 sky130_fd_sc_hd__o32a_1 _20709_ (.A1(_02010_),
    .A2(_02185_),
    .A3(_10546_),
    .B1(_10542_),
    .B2(_10191_),
    .X(_10797_));
 sky130_fd_sc_hd__o21a_4 _20710_ (.A1(_10468_),
    .A2(_10116_),
    .B1(_10119_),
    .X(_10798_));
 sky130_fd_sc_hd__o21ai_4 _20711_ (.A1(_10468_),
    .A2(_10116_),
    .B1(_10119_),
    .Y(_10799_));
 sky130_fd_sc_hd__nand2_2 _20712_ (.A(net41),
    .B(net22),
    .Y(_10800_));
 sky130_fd_sc_hd__a22oi_4 _20713_ (.A1(net40),
    .A2(net24),
    .B1(net25),
    .B2(net39),
    .Y(_10801_));
 sky130_fd_sc_hd__a22o_2 _20714_ (.A1(net40),
    .A2(net24),
    .B1(net25),
    .B2(net39),
    .X(_10802_));
 sky130_fd_sc_hd__and3_4 _20715_ (.A(net39),
    .B(net40),
    .C(net25),
    .X(_10803_));
 sky130_fd_sc_hd__nand3_4 _20716_ (.A(net39),
    .B(net40),
    .C(net25),
    .Y(_10804_));
 sky130_fd_sc_hd__and4_2 _20717_ (.A(net39),
    .B(net40),
    .C(net24),
    .D(net25),
    .X(_10805_));
 sky130_fd_sc_hd__o21bai_4 _20718_ (.A1(_10801_),
    .A2(_10805_),
    .B1_N(_10800_),
    .Y(_10807_));
 sky130_fd_sc_hd__o221ai_4 _20719_ (.A1(_02010_),
    .A2(_02196_),
    .B1(_02218_),
    .B2(_10804_),
    .C1(_10802_),
    .Y(_10808_));
 sky130_fd_sc_hd__o2111ai_4 _20720_ (.A1(_02218_),
    .A2(_10804_),
    .B1(net41),
    .C1(net22),
    .D1(_10802_),
    .Y(_10809_));
 sky130_fd_sc_hd__o21ai_4 _20721_ (.A1(_10801_),
    .A2(_10805_),
    .B1(_10800_),
    .Y(_10810_));
 sky130_fd_sc_hd__a21oi_4 _20722_ (.A1(_10807_),
    .A2(_10808_),
    .B1(_10798_),
    .Y(_10811_));
 sky130_fd_sc_hd__a22o_1 _20723_ (.A1(_10119_),
    .A2(_10470_),
    .B1(_10807_),
    .B2(_10808_),
    .X(_10812_));
 sky130_fd_sc_hd__a21oi_4 _20724_ (.A1(_10809_),
    .A2(_10810_),
    .B1(_10799_),
    .Y(_10813_));
 sky130_fd_sc_hd__nand4_1 _20725_ (.A(_10119_),
    .B(_10470_),
    .C(_10807_),
    .D(_10808_),
    .Y(_10814_));
 sky130_fd_sc_hd__o22ai_1 _20726_ (.A1(_10544_),
    .A2(_10794_),
    .B1(_10811_),
    .B2(_10813_),
    .Y(_10815_));
 sky130_fd_sc_hd__o211ai_1 _20727_ (.A1(_10546_),
    .A2(_10793_),
    .B1(_10812_),
    .C1(_10814_),
    .Y(_10816_));
 sky130_fd_sc_hd__a31oi_2 _20728_ (.A1(_10798_),
    .A2(_10807_),
    .A3(_10808_),
    .B1(_10797_),
    .Y(_10818_));
 sky130_fd_sc_hd__a31o_1 _20729_ (.A1(_10798_),
    .A2(_10807_),
    .A3(_10808_),
    .B1(_10797_),
    .X(_10819_));
 sky130_fd_sc_hd__o22ai_2 _20730_ (.A1(_10546_),
    .A2(_10793_),
    .B1(_10811_),
    .B2(_10813_),
    .Y(_10820_));
 sky130_fd_sc_hd__o211a_1 _20731_ (.A1(_10811_),
    .A2(_10819_),
    .B1(_10820_),
    .C1(_10792_),
    .X(_10821_));
 sky130_fd_sc_hd__o211ai_4 _20732_ (.A1(_10811_),
    .A2(_10819_),
    .B1(_10820_),
    .C1(_10792_),
    .Y(_10822_));
 sky130_fd_sc_hd__nand3_2 _20733_ (.A(_10815_),
    .B(_10816_),
    .C(_10791_),
    .Y(_10823_));
 sky130_fd_sc_hd__nand4_2 _20734_ (.A(_10787_),
    .B(_10788_),
    .C(_10822_),
    .D(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__a22o_1 _20735_ (.A1(_10787_),
    .A2(_10788_),
    .B1(_10822_),
    .B2(_10823_),
    .X(_10825_));
 sky130_fd_sc_hd__and3_1 _20736_ (.A(_10789_),
    .B(_10790_),
    .C(_10823_),
    .X(_10826_));
 sky130_fd_sc_hd__nand4_2 _20737_ (.A(_10789_),
    .B(_10790_),
    .C(_10822_),
    .D(_10823_),
    .Y(_10827_));
 sky130_fd_sc_hd__a22o_1 _20738_ (.A1(_10789_),
    .A2(_10790_),
    .B1(_10822_),
    .B2(_10823_),
    .X(_10829_));
 sky130_fd_sc_hd__o211a_1 _20739_ (.A1(_10481_),
    .A2(_10483_),
    .B1(_10827_),
    .C1(_10829_),
    .X(_10830_));
 sky130_fd_sc_hd__o211ai_4 _20740_ (.A1(_10481_),
    .A2(_10483_),
    .B1(_10827_),
    .C1(_10829_),
    .Y(_10831_));
 sky130_fd_sc_hd__nand3_4 _20741_ (.A(_10825_),
    .B(_10760_),
    .C(_10824_),
    .Y(_10832_));
 sky130_fd_sc_hd__inv_2 _20742_ (.A(_10832_),
    .Y(_10833_));
 sky130_fd_sc_hd__o2111ai_4 _20743_ (.A1(_10531_),
    .A2(_10567_),
    .B1(_10831_),
    .C1(_10832_),
    .D1(_10566_),
    .Y(_10834_));
 sky130_fd_sc_hd__a21bo_1 _20744_ (.A1(_10831_),
    .A2(_10832_),
    .B1_N(_10759_),
    .X(_10835_));
 sky130_fd_sc_hd__o311a_2 _20745_ (.A1(_10526_),
    .A2(_10527_),
    .A3(_10564_),
    .B1(_10568_),
    .C1(_10832_),
    .X(_10836_));
 sky130_fd_sc_hd__nand3_2 _20746_ (.A(_10831_),
    .B(_10832_),
    .C(_10759_),
    .Y(_10837_));
 sky130_fd_sc_hd__a21oi_1 _20747_ (.A1(_10831_),
    .A2(_10832_),
    .B1(_10759_),
    .Y(_10838_));
 sky130_fd_sc_hd__a21o_1 _20748_ (.A1(_10831_),
    .A2(_10832_),
    .B1(_10759_),
    .X(_10840_));
 sky130_fd_sc_hd__nand4_2 _20749_ (.A(_10756_),
    .B(_10758_),
    .C(_10834_),
    .D(_10835_),
    .Y(_10841_));
 sky130_fd_sc_hd__o211ai_2 _20750_ (.A1(_10755_),
    .A2(_10757_),
    .B1(_10837_),
    .C1(_10840_),
    .Y(_10842_));
 sky130_fd_sc_hd__nand4_4 _20751_ (.A(_10756_),
    .B(_10758_),
    .C(_10837_),
    .D(_10840_),
    .Y(_10843_));
 sky130_fd_sc_hd__o211ai_2 _20752_ (.A1(_10755_),
    .A2(_10757_),
    .B1(_10834_),
    .C1(_10835_),
    .Y(_10844_));
 sky130_fd_sc_hd__a21oi_2 _20753_ (.A1(_10841_),
    .A2(_10842_),
    .B1(_10742_),
    .Y(_10845_));
 sky130_fd_sc_hd__o211ai_1 _20754_ (.A1(_10494_),
    .A2(_10591_),
    .B1(_10843_),
    .C1(_10844_),
    .Y(_10846_));
 sky130_fd_sc_hd__a21oi_1 _20755_ (.A1(_10843_),
    .A2(_10844_),
    .B1(_10743_),
    .Y(_10847_));
 sky130_fd_sc_hd__nand3_1 _20756_ (.A(_10742_),
    .B(_10841_),
    .C(_10842_),
    .Y(_10848_));
 sky130_fd_sc_hd__o22ai_1 _20757_ (.A1(_10738_),
    .A2(_10739_),
    .B1(_10845_),
    .B2(_10847_),
    .Y(_10849_));
 sky130_fd_sc_hd__nand4b_1 _20758_ (.A_N(_10738_),
    .B(_10741_),
    .C(_10846_),
    .D(_10848_),
    .Y(_10851_));
 sky130_fd_sc_hd__o2bb2ai_1 _20759_ (.A1_N(_10736_),
    .A2_N(_10737_),
    .B1(_10845_),
    .B2(_10847_),
    .Y(_10852_));
 sky130_fd_sc_hd__nand4_1 _20760_ (.A(_10736_),
    .B(_10737_),
    .C(_10846_),
    .D(_10848_),
    .Y(_10853_));
 sky130_fd_sc_hd__a22oi_1 _20761_ (.A1(_10594_),
    .A2(_10639_),
    .B1(_10849_),
    .B2(_10851_),
    .Y(_10854_));
 sky130_fd_sc_hd__nand3_1 _20762_ (.A(_10640_),
    .B(_10852_),
    .C(_10853_),
    .Y(_10855_));
 sky130_fd_sc_hd__a21oi_1 _20763_ (.A1(_10852_),
    .A2(_10853_),
    .B1(_10640_),
    .Y(_10856_));
 sky130_fd_sc_hd__a21o_1 _20764_ (.A1(_10852_),
    .A2(_10853_),
    .B1(_10640_),
    .X(_10857_));
 sky130_fd_sc_hd__o211a_1 _20765_ (.A1(_10451_),
    .A2(_10459_),
    .B1(_10855_),
    .C1(_10857_),
    .X(_10858_));
 sky130_fd_sc_hd__o211ai_2 _20766_ (.A1(_10451_),
    .A2(_10459_),
    .B1(_10855_),
    .C1(_10857_),
    .Y(_10859_));
 sky130_fd_sc_hd__o22ai_2 _20767_ (.A1(_10450_),
    .A2(_10637_),
    .B1(_10854_),
    .B2(_10856_),
    .Y(_10860_));
 sky130_fd_sc_hd__o211a_1 _20768_ (.A1(_10322_),
    .A2(_10319_),
    .B1(_10318_),
    .C1(_10607_),
    .X(_10862_));
 sky130_fd_sc_hd__o2bb2ai_2 _20769_ (.A1_N(_10859_),
    .A2_N(_10860_),
    .B1(_10862_),
    .B2(_10605_),
    .Y(_10863_));
 sky130_fd_sc_hd__o21ai_1 _20770_ (.A1(_10606_),
    .A2(_10612_),
    .B1(_10860_),
    .Y(_10864_));
 sky130_fd_sc_hd__o211ai_2 _20771_ (.A1(_10606_),
    .A2(_10612_),
    .B1(_10859_),
    .C1(_10860_),
    .Y(_10865_));
 sky130_fd_sc_hd__o21ai_2 _20772_ (.A1(_10296_),
    .A2(_10431_),
    .B1(_10435_),
    .Y(_10866_));
 sky130_fd_sc_hd__a21o_1 _20773_ (.A1(_10863_),
    .A2(_10865_),
    .B1(_10866_),
    .X(_10867_));
 sky130_fd_sc_hd__o211ai_1 _20774_ (.A1(_10858_),
    .A2(_10864_),
    .B1(_10866_),
    .C1(_10863_),
    .Y(_10868_));
 sky130_fd_sc_hd__a22o_1 _20775_ (.A1(_10435_),
    .A2(_10438_),
    .B1(_10863_),
    .B2(_10865_),
    .X(_10869_));
 sky130_fd_sc_hd__o2111ai_2 _20776_ (.A1(_10296_),
    .A2(_10431_),
    .B1(_10435_),
    .C1(_10863_),
    .D1(_10865_),
    .Y(_10870_));
 sky130_fd_sc_hd__nand2_1 _20777_ (.A(_10869_),
    .B(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__a21oi_1 _20778_ (.A1(_10617_),
    .A2(_10622_),
    .B1(_10618_),
    .Y(_10873_));
 sky130_fd_sc_hd__o21ai_1 _20779_ (.A1(_10371_),
    .A2(_10616_),
    .B1(_10626_),
    .Y(_10874_));
 sky130_fd_sc_hd__nand3_1 _20780_ (.A(_10869_),
    .B(_10873_),
    .C(_10870_),
    .Y(_10875_));
 sky130_fd_sc_hd__nand3_1 _20781_ (.A(_10867_),
    .B(_10868_),
    .C(_10874_),
    .Y(_10876_));
 sky130_fd_sc_hd__nand2_1 _20782_ (.A(_10875_),
    .B(_10876_),
    .Y(_10877_));
 sky130_fd_sc_hd__o2111ai_4 _20783_ (.A1(_10632_),
    .A2(_10623_),
    .B1(_10360_),
    .C1(_10359_),
    .D1(_10630_),
    .Y(_10878_));
 sky130_fd_sc_hd__o31a_1 _20784_ (.A1(_10623_),
    .A2(_10628_),
    .A3(_10625_),
    .B1(_10360_),
    .X(_10879_));
 sky130_fd_sc_hd__a21o_1 _20785_ (.A1(_10360_),
    .A2(_10633_),
    .B1(_10629_),
    .X(_10880_));
 sky130_fd_sc_hd__o21ai_1 _20786_ (.A1(_10878_),
    .A2(_10366_),
    .B1(_10880_),
    .Y(_10881_));
 sky130_fd_sc_hd__xnor2_2 _20787_ (.A(_10877_),
    .B(_10881_),
    .Y(net105));
 sky130_fd_sc_hd__nand2_1 _20788_ (.A(_10758_),
    .B(_10837_),
    .Y(_10883_));
 sky130_fd_sc_hd__o21bai_1 _20789_ (.A1(_10838_),
    .A2(_10883_),
    .B1_N(_10755_),
    .Y(_10884_));
 sky130_fd_sc_hd__a21oi_4 _20790_ (.A1(_10747_),
    .A2(_10749_),
    .B1(_09384_),
    .Y(_10885_));
 sky130_fd_sc_hd__a211o_4 _20791_ (.A1(_10747_),
    .A2(_10749_),
    .B1(_08004_),
    .C1(_08959_),
    .X(_10886_));
 sky130_fd_sc_hd__and3_4 _20792_ (.A(_10747_),
    .B(_10749_),
    .C(_09385_),
    .X(_10887_));
 sky130_fd_sc_hd__nand4_4 _20793_ (.A(_10747_),
    .B(_08006_),
    .C(_08963_),
    .D(_10749_),
    .Y(_10888_));
 sky130_fd_sc_hd__a21oi_4 _20794_ (.A1(_09385_),
    .A2(_10750_),
    .B1(_10885_),
    .Y(_10889_));
 sky130_fd_sc_hd__o21ai_4 _20795_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .Y(_10890_));
 sky130_fd_sc_hd__a31o_1 _20796_ (.A1(_10789_),
    .A2(_10790_),
    .A3(_10823_),
    .B1(_10821_),
    .X(_10891_));
 sky130_fd_sc_hd__a21boi_4 _20797_ (.A1(_10479_),
    .A2(_10745_),
    .B1_N(_10482_),
    .Y(_10892_));
 sky130_fd_sc_hd__o2bb2ai_4 _20798_ (.A1_N(_10479_),
    .A2_N(_10745_),
    .B1(_10480_),
    .B2(_10473_),
    .Y(_10894_));
 sky130_fd_sc_hd__nand2_1 _20799_ (.A(net48),
    .B(net17),
    .Y(_10895_));
 sky130_fd_sc_hd__nand4_2 _20800_ (.A(net46),
    .B(net47),
    .C(net18),
    .D(net19),
    .Y(_10896_));
 sky130_fd_sc_hd__a22oi_1 _20801_ (.A1(net47),
    .A2(net18),
    .B1(net19),
    .B2(net46),
    .Y(_10897_));
 sky130_fd_sc_hd__a22o_1 _20802_ (.A1(net47),
    .A2(net18),
    .B1(net19),
    .B2(net46),
    .X(_10898_));
 sky130_fd_sc_hd__a22oi_1 _20803_ (.A1(net48),
    .A2(net17),
    .B1(_10896_),
    .B2(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__a22o_1 _20804_ (.A1(net48),
    .A2(net17),
    .B1(_10896_),
    .B2(_10898_),
    .X(_10900_));
 sky130_fd_sc_hd__and4_1 _20805_ (.A(_10898_),
    .B(net17),
    .C(net48),
    .D(_10896_),
    .X(_10901_));
 sky130_fd_sc_hd__nand4_1 _20806_ (.A(_10898_),
    .B(net17),
    .C(net48),
    .D(_10896_),
    .Y(_10902_));
 sky130_fd_sc_hd__nor2_1 _20807_ (.A(_10899_),
    .B(_10901_),
    .Y(_10903_));
 sky130_fd_sc_hd__nand2_1 _20808_ (.A(_10900_),
    .B(_10902_),
    .Y(_10905_));
 sky130_fd_sc_hd__o31ai_4 _20809_ (.A1(_02054_),
    .A2(_02142_),
    .A3(_10768_),
    .B1(_10767_),
    .Y(_10906_));
 sky130_fd_sc_hd__and2_1 _20810_ (.A(net45),
    .B(net20),
    .X(_10907_));
 sky130_fd_sc_hd__nand2_2 _20811_ (.A(net43),
    .B(net22),
    .Y(_10908_));
 sky130_fd_sc_hd__nand4_1 _20812_ (.A(net42),
    .B(net43),
    .C(net21),
    .D(net22),
    .Y(_10909_));
 sky130_fd_sc_hd__a22o_2 _20813_ (.A1(net43),
    .A2(net21),
    .B1(net22),
    .B2(net42),
    .X(_10910_));
 sky130_fd_sc_hd__o211a_1 _20814_ (.A1(_10766_),
    .A2(_10908_),
    .B1(_10907_),
    .C1(_10910_),
    .X(_10911_));
 sky130_fd_sc_hd__o2111ai_4 _20815_ (.A1(_10766_),
    .A2(_10908_),
    .B1(net45),
    .C1(net20),
    .D1(_10910_),
    .Y(_10912_));
 sky130_fd_sc_hd__a21oi_1 _20816_ (.A1(_10909_),
    .A2(_10910_),
    .B1(_10907_),
    .Y(_10913_));
 sky130_fd_sc_hd__o2bb2ai_1 _20817_ (.A1_N(_10909_),
    .A2_N(_10910_),
    .B1(_02054_),
    .B2(_02163_),
    .Y(_10914_));
 sky130_fd_sc_hd__and3_1 _20818_ (.A(_10906_),
    .B(_10912_),
    .C(_10914_),
    .X(_10916_));
 sky130_fd_sc_hd__nand3_2 _20819_ (.A(_10906_),
    .B(_10912_),
    .C(_10914_),
    .Y(_10917_));
 sky130_fd_sc_hd__a21oi_1 _20820_ (.A1(_10912_),
    .A2(_10914_),
    .B1(_10906_),
    .Y(_10918_));
 sky130_fd_sc_hd__o21bai_1 _20821_ (.A1(_10911_),
    .A2(_10913_),
    .B1_N(_10906_),
    .Y(_10919_));
 sky130_fd_sc_hd__nor2_1 _20822_ (.A(_10905_),
    .B(_10918_),
    .Y(_10920_));
 sky130_fd_sc_hd__nand2_1 _20823_ (.A(_10919_),
    .B(_10903_),
    .Y(_10921_));
 sky130_fd_sc_hd__a21oi_1 _20824_ (.A1(_10917_),
    .A2(_10919_),
    .B1(_10903_),
    .Y(_10922_));
 sky130_fd_sc_hd__a22o_1 _20825_ (.A1(_10900_),
    .A2(_10902_),
    .B1(_10917_),
    .B2(_10919_),
    .X(_10923_));
 sky130_fd_sc_hd__a21oi_1 _20826_ (.A1(_10917_),
    .A2(_10920_),
    .B1(_10922_),
    .Y(_10924_));
 sky130_fd_sc_hd__a31oi_4 _20827_ (.A1(_10799_),
    .A2(_10809_),
    .A3(_10810_),
    .B1(_10796_),
    .Y(_10925_));
 sky130_fd_sc_hd__nor2_1 _20828_ (.A(_02010_),
    .B(_02218_),
    .Y(_10927_));
 sky130_fd_sc_hd__o21ai_2 _20829_ (.A1(net39),
    .A2(net40),
    .B1(net25),
    .Y(_10928_));
 sky130_fd_sc_hd__o21a_4 _20830_ (.A1(net39),
    .A2(net40),
    .B1(net25),
    .X(_10929_));
 sky130_fd_sc_hd__o2bb2ai_2 _20831_ (.A1_N(_10804_),
    .A2_N(_10929_),
    .B1(_02010_),
    .B2(_02218_),
    .Y(_10930_));
 sky130_fd_sc_hd__and3_1 _20832_ (.A(_10929_),
    .B(net24),
    .C(net41),
    .X(_10931_));
 sky130_fd_sc_hd__o2111ai_4 _20833_ (.A1(net39),
    .A2(net40),
    .B1(net41),
    .C1(net24),
    .D1(net25),
    .Y(_10932_));
 sky130_fd_sc_hd__o211ai_2 _20834_ (.A1(_02010_),
    .A2(_02218_),
    .B1(_10804_),
    .C1(_10929_),
    .Y(_10933_));
 sky130_fd_sc_hd__o21ai_1 _20835_ (.A1(_10803_),
    .A2(_10928_),
    .B1(_10927_),
    .Y(_10934_));
 sky130_fd_sc_hd__nand3_4 _20836_ (.A(_10934_),
    .B(_10798_),
    .C(_10933_),
    .Y(_10935_));
 sky130_fd_sc_hd__o211a_1 _20837_ (.A1(_10932_),
    .A2(_10803_),
    .B1(_10799_),
    .C1(_10930_),
    .X(_10936_));
 sky130_fd_sc_hd__o211ai_4 _20838_ (.A1(_10932_),
    .A2(_10803_),
    .B1(_10799_),
    .C1(_10930_),
    .Y(_10938_));
 sky130_fd_sc_hd__and3_1 _20839_ (.A(_10802_),
    .B(net22),
    .C(net41),
    .X(_10939_));
 sky130_fd_sc_hd__a31o_1 _20840_ (.A1(_10802_),
    .A2(net22),
    .A3(net41),
    .B1(_10805_),
    .X(_10940_));
 sky130_fd_sc_hd__o211a_1 _20841_ (.A1(_10805_),
    .A2(_10939_),
    .B1(_10938_),
    .C1(_10935_),
    .X(_10941_));
 sky130_fd_sc_hd__o211ai_2 _20842_ (.A1(_10805_),
    .A2(_10939_),
    .B1(_10938_),
    .C1(_10935_),
    .Y(_10942_));
 sky130_fd_sc_hd__a21oi_2 _20843_ (.A1(_10935_),
    .A2(_10938_),
    .B1(_10940_),
    .Y(_10943_));
 sky130_fd_sc_hd__a21o_1 _20844_ (.A1(_10935_),
    .A2(_10938_),
    .B1(_10940_),
    .X(_10944_));
 sky130_fd_sc_hd__o211a_1 _20845_ (.A1(_10811_),
    .A2(_10818_),
    .B1(_10942_),
    .C1(_10944_),
    .X(_10945_));
 sky130_fd_sc_hd__o211ai_4 _20846_ (.A1(_10811_),
    .A2(_10818_),
    .B1(_10942_),
    .C1(_10944_),
    .Y(_10946_));
 sky130_fd_sc_hd__o22ai_4 _20847_ (.A1(_10813_),
    .A2(_10925_),
    .B1(_10941_),
    .B2(_10943_),
    .Y(_10947_));
 sky130_fd_sc_hd__o2111a_2 _20848_ (.A1(_10916_),
    .A2(_10921_),
    .B1(_10923_),
    .C1(_10946_),
    .D1(_10947_),
    .X(_10949_));
 sky130_fd_sc_hd__o2111ai_2 _20849_ (.A1(_10916_),
    .A2(_10921_),
    .B1(_10923_),
    .C1(_10946_),
    .D1(_10947_),
    .Y(_10950_));
 sky130_fd_sc_hd__a21oi_2 _20850_ (.A1(_10946_),
    .A2(_10947_),
    .B1(_10924_),
    .Y(_10951_));
 sky130_fd_sc_hd__a21o_1 _20851_ (.A1(_10946_),
    .A2(_10947_),
    .B1(_10924_),
    .X(_10952_));
 sky130_fd_sc_hd__nor3_2 _20852_ (.A(_10892_),
    .B(_10949_),
    .C(_10951_),
    .Y(_10953_));
 sky130_fd_sc_hd__o211ai_2 _20853_ (.A1(_10481_),
    .A2(_10748_),
    .B1(_10950_),
    .C1(_10952_),
    .Y(_10954_));
 sky130_fd_sc_hd__o21a_1 _20854_ (.A1(_10949_),
    .A2(_10951_),
    .B1(_10892_),
    .X(_10955_));
 sky130_fd_sc_hd__o21ai_2 _20855_ (.A1(_10949_),
    .A2(_10951_),
    .B1(_10892_),
    .Y(_10956_));
 sky130_fd_sc_hd__o21ai_2 _20856_ (.A1(_10953_),
    .A2(_10955_),
    .B1(_10891_),
    .Y(_10957_));
 sky130_fd_sc_hd__nand3b_2 _20857_ (.A_N(_10891_),
    .B(_10954_),
    .C(_10956_),
    .Y(_10958_));
 sky130_fd_sc_hd__o21a_1 _20858_ (.A1(_10821_),
    .A2(_10826_),
    .B1(_10956_),
    .X(_10960_));
 sky130_fd_sc_hd__o211ai_2 _20859_ (.A1(_10821_),
    .A2(_10826_),
    .B1(_10954_),
    .C1(_10956_),
    .Y(_10961_));
 sky130_fd_sc_hd__a21o_1 _20860_ (.A1(_10954_),
    .A2(_10956_),
    .B1(_10891_),
    .X(_10962_));
 sky130_fd_sc_hd__and3_1 _20861_ (.A(_10962_),
    .B(_10889_),
    .C(_10961_),
    .X(_10963_));
 sky130_fd_sc_hd__o2111ai_1 _20862_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .C1(_10961_),
    .D1(_10962_),
    .Y(_10964_));
 sky130_fd_sc_hd__o211ai_2 _20863_ (.A1(_10885_),
    .A2(_10887_),
    .B1(_10957_),
    .C1(_10958_),
    .Y(_10965_));
 sky130_fd_sc_hd__nand3_1 _20864_ (.A(_10957_),
    .B(_10958_),
    .C(_10889_),
    .Y(_10966_));
 sky130_fd_sc_hd__o211ai_2 _20865_ (.A1(_10885_),
    .A2(_10887_),
    .B1(_10961_),
    .C1(_10962_),
    .Y(_10967_));
 sky130_fd_sc_hd__nand4_4 _20866_ (.A(_10756_),
    .B(_10843_),
    .C(_10966_),
    .D(_10967_),
    .Y(_10968_));
 sky130_fd_sc_hd__inv_2 _20867_ (.A(_10968_),
    .Y(_10969_));
 sky130_fd_sc_hd__nand2_2 _20868_ (.A(_10884_),
    .B(_10965_),
    .Y(_10971_));
 sky130_fd_sc_hd__nand3_1 _20869_ (.A(_10884_),
    .B(_10964_),
    .C(_10965_),
    .Y(_10972_));
 sky130_fd_sc_hd__nand2_1 _20870_ (.A(_10968_),
    .B(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__o22a_1 _20871_ (.A1(_02098_),
    .A2(_02109_),
    .B1(_10500_),
    .B2(_10779_),
    .X(_10974_));
 sky130_fd_sc_hd__o31ai_2 _20872_ (.A1(_02098_),
    .A2(_02109_),
    .A3(_10777_),
    .B1(_10780_),
    .Y(_10975_));
 sky130_fd_sc_hd__nand2_2 _20873_ (.A(net16),
    .B(net50),
    .Y(_10976_));
 sky130_fd_sc_hd__nand2_1 _20874_ (.A(net16),
    .B(net49),
    .Y(_10977_));
 sky130_fd_sc_hd__and4_1 _20875_ (.A(net15),
    .B(net16),
    .C(net49),
    .D(net50),
    .X(_10978_));
 sky130_fd_sc_hd__nand4_1 _20876_ (.A(net15),
    .B(net16),
    .C(net49),
    .D(net50),
    .Y(_10979_));
 sky130_fd_sc_hd__a22oi_1 _20877_ (.A1(net16),
    .A2(net49),
    .B1(net50),
    .B2(net15),
    .Y(_10980_));
 sky130_fd_sc_hd__a22o_2 _20878_ (.A1(net16),
    .A2(net49),
    .B1(net50),
    .B2(net15),
    .X(_10982_));
 sky130_fd_sc_hd__a2bb2oi_2 _20879_ (.A1_N(_02065_),
    .A2_N(_02152_),
    .B1(_10979_),
    .B2(_10982_),
    .Y(_10983_));
 sky130_fd_sc_hd__a22o_1 _20880_ (.A1(net14),
    .A2(net51),
    .B1(_10979_),
    .B2(_10982_),
    .X(_10984_));
 sky130_fd_sc_hd__o2111a_1 _20881_ (.A1(_10648_),
    .A2(_10976_),
    .B1(net14),
    .C1(net51),
    .D1(_10982_),
    .X(_10985_));
 sky130_fd_sc_hd__o2111ai_4 _20882_ (.A1(_10648_),
    .A2(_10976_),
    .B1(net14),
    .C1(net51),
    .D1(_10982_),
    .Y(_10986_));
 sky130_fd_sc_hd__o22ai_4 _20883_ (.A1(_10777_),
    .A2(_10974_),
    .B1(_10983_),
    .B2(_10985_),
    .Y(_10987_));
 sky130_fd_sc_hd__nand3_4 _20884_ (.A(_10984_),
    .B(_10986_),
    .C(_10975_),
    .Y(_10988_));
 sky130_fd_sc_hd__and3_1 _20885_ (.A(_10650_),
    .B(net51),
    .C(net13),
    .X(_10989_));
 sky130_fd_sc_hd__a31o_1 _20886_ (.A1(_10650_),
    .A2(net51),
    .A3(net13),
    .B1(_10651_),
    .X(_10990_));
 sky130_fd_sc_hd__a21o_1 _20887_ (.A1(_10987_),
    .A2(_10988_),
    .B1(_10990_),
    .X(_10991_));
 sky130_fd_sc_hd__o21ai_2 _20888_ (.A1(_10651_),
    .A2(_10989_),
    .B1(_10987_),
    .Y(_10993_));
 sky130_fd_sc_hd__o211ai_2 _20889_ (.A1(_10651_),
    .A2(_10989_),
    .B1(_10988_),
    .C1(_10987_),
    .Y(_10994_));
 sky130_fd_sc_hd__o2111ai_1 _20890_ (.A1(_10647_),
    .A2(_10649_),
    .B1(_10653_),
    .C1(_10987_),
    .D1(_10988_),
    .Y(_10995_));
 sky130_fd_sc_hd__o2bb2ai_1 _20891_ (.A1_N(_10987_),
    .A2_N(_10988_),
    .B1(_10989_),
    .B2(_10651_),
    .Y(_10996_));
 sky130_fd_sc_hd__o2bb2ai_1 _20892_ (.A1_N(_10786_),
    .A2_N(_10774_),
    .B1(_10772_),
    .B2(_10775_),
    .Y(_10997_));
 sky130_fd_sc_hd__a2bb2oi_1 _20893_ (.A1_N(_10772_),
    .A2_N(_10775_),
    .B1(_10786_),
    .B2(_10774_),
    .Y(_10998_));
 sky130_fd_sc_hd__nand3_2 _20894_ (.A(_10995_),
    .B(_10996_),
    .C(_10998_),
    .Y(_10999_));
 sky130_fd_sc_hd__nand3_4 _20895_ (.A(_10991_),
    .B(_10997_),
    .C(_10994_),
    .Y(_11000_));
 sky130_fd_sc_hd__o311a_1 _20896_ (.A1(_02032_),
    .A2(_02152_),
    .A3(_10379_),
    .B1(_10382_),
    .C1(_10661_),
    .X(_11001_));
 sky130_fd_sc_hd__o2bb2ai_4 _20897_ (.A1_N(_10999_),
    .A2_N(_11000_),
    .B1(_11001_),
    .B2(_10659_),
    .Y(_11002_));
 sky130_fd_sc_hd__o211ai_4 _20898_ (.A1(_10660_),
    .A2(_10666_),
    .B1(_10999_),
    .C1(_11000_),
    .Y(_11004_));
 sky130_fd_sc_hd__a32oi_2 _20899_ (.A1(_10668_),
    .A2(_10669_),
    .A3(_10670_),
    .B1(_10673_),
    .B2(_10644_),
    .Y(_11005_));
 sky130_fd_sc_hd__a21oi_2 _20900_ (.A1(_11002_),
    .A2(_11004_),
    .B1(_11005_),
    .Y(_11006_));
 sky130_fd_sc_hd__a21o_2 _20901_ (.A1(_11002_),
    .A2(_11004_),
    .B1(_11005_),
    .X(_11007_));
 sky130_fd_sc_hd__o211a_4 _20902_ (.A1(_10672_),
    .A2(_10678_),
    .B1(_11002_),
    .C1(_11004_),
    .X(_11008_));
 sky130_fd_sc_hd__o211ai_4 _20903_ (.A1(_10672_),
    .A2(_10678_),
    .B1(_11002_),
    .C1(_11004_),
    .Y(_11009_));
 sky130_fd_sc_hd__o2bb2a_1 _20904_ (.A1_N(_10690_),
    .A2_N(_10706_),
    .B1(_10708_),
    .B2(_10704_),
    .X(_11010_));
 sky130_fd_sc_hd__a2bb2o_1 _20905_ (.A1_N(_10704_),
    .A2_N(_10708_),
    .B1(_10706_),
    .B2(_10690_),
    .X(_11011_));
 sky130_fd_sc_hd__a22o_1 _20906_ (.A1(net9),
    .A2(net56),
    .B1(_01988_),
    .B2(net57),
    .X(_11012_));
 sky130_fd_sc_hd__nand4_4 _20907_ (.A(_01988_),
    .B(net9),
    .C(net56),
    .D(net57),
    .Y(_11013_));
 sky130_fd_sc_hd__nand2_1 _20908_ (.A(_11012_),
    .B(_11013_),
    .Y(_11015_));
 sky130_fd_sc_hd__nand2_1 _20909_ (.A(net10),
    .B(net54),
    .Y(_11016_));
 sky130_fd_sc_hd__nand2_1 _20910_ (.A(net13),
    .B(net53),
    .Y(_11017_));
 sky130_fd_sc_hd__nand4_1 _20911_ (.A(net11),
    .B(net13),
    .C(net52),
    .D(net53),
    .Y(_11018_));
 sky130_fd_sc_hd__nand2_1 _20912_ (.A(net13),
    .B(net52),
    .Y(_11019_));
 sky130_fd_sc_hd__a22oi_1 _20913_ (.A1(net13),
    .A2(net52),
    .B1(net53),
    .B2(net11),
    .Y(_11020_));
 sky130_fd_sc_hd__a22o_1 _20914_ (.A1(net13),
    .A2(net52),
    .B1(net53),
    .B2(net11),
    .X(_11021_));
 sky130_fd_sc_hd__o2bb2ai_1 _20915_ (.A1_N(_10698_),
    .A2_N(_11019_),
    .B1(_11017_),
    .B2(_10694_),
    .Y(_11022_));
 sky130_fd_sc_hd__o21ai_2 _20916_ (.A1(_02021_),
    .A2(_02207_),
    .B1(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__o2111ai_4 _20917_ (.A1(_10694_),
    .A2(_11017_),
    .B1(net10),
    .C1(net54),
    .D1(_11021_),
    .Y(_11024_));
 sky130_fd_sc_hd__o22a_1 _20918_ (.A1(_01999_),
    .A2(_02207_),
    .B1(_10414_),
    .B2(_10694_),
    .X(_11026_));
 sky130_fd_sc_hd__a21o_1 _20919_ (.A1(_10414_),
    .A2(_10694_),
    .B1(_10693_),
    .X(_11027_));
 sky130_fd_sc_hd__o21ai_1 _20920_ (.A1(_10693_),
    .A2(_10695_),
    .B1(_10700_),
    .Y(_11028_));
 sky130_fd_sc_hd__a21oi_1 _20921_ (.A1(_11023_),
    .A2(_11024_),
    .B1(_11028_),
    .Y(_11029_));
 sky130_fd_sc_hd__o2bb2ai_2 _20922_ (.A1_N(_11023_),
    .A2_N(_11024_),
    .B1(_11026_),
    .B2(_10695_),
    .Y(_11030_));
 sky130_fd_sc_hd__a22oi_1 _20923_ (.A1(_11016_),
    .A2(_11022_),
    .B1(_11027_),
    .B2(_10700_),
    .Y(_11031_));
 sky130_fd_sc_hd__and3_1 _20924_ (.A(_11023_),
    .B(_11028_),
    .C(_11024_),
    .X(_11032_));
 sky130_fd_sc_hd__nand3_2 _20925_ (.A(_11023_),
    .B(_11024_),
    .C(_11028_),
    .Y(_11033_));
 sky130_fd_sc_hd__a22oi_1 _20926_ (.A1(_11012_),
    .A2(_11013_),
    .B1(_11030_),
    .B2(_11033_),
    .Y(_11034_));
 sky130_fd_sc_hd__a22o_1 _20927_ (.A1(_11012_),
    .A2(_11013_),
    .B1(_11030_),
    .B2(_11033_),
    .X(_11035_));
 sky130_fd_sc_hd__a211oi_2 _20928_ (.A1(_11031_),
    .A2(_11024_),
    .B1(_11015_),
    .C1(_11029_),
    .Y(_11037_));
 sky130_fd_sc_hd__nand4_4 _20929_ (.A(_11012_),
    .B(_11013_),
    .C(_11030_),
    .D(_11033_),
    .Y(_11038_));
 sky130_fd_sc_hd__nand2_1 _20930_ (.A(_11035_),
    .B(_11038_),
    .Y(_11039_));
 sky130_fd_sc_hd__o221a_1 _20931_ (.A1(_10704_),
    .A2(_10708_),
    .B1(_11034_),
    .B2(_11037_),
    .C1(_10713_),
    .X(_11040_));
 sky130_fd_sc_hd__o21ai_1 _20932_ (.A1(_11034_),
    .A2(_11037_),
    .B1(_11010_),
    .Y(_11041_));
 sky130_fd_sc_hd__nand3_4 _20933_ (.A(_11011_),
    .B(_11035_),
    .C(_11038_),
    .Y(_11042_));
 sky130_fd_sc_hd__a22oi_2 _20934_ (.A1(net57),
    .A2(_10688_),
    .B1(_11041_),
    .B2(_11042_),
    .Y(_11043_));
 sky130_fd_sc_hd__a21oi_1 _20935_ (.A1(_11039_),
    .A2(_11010_),
    .B1(_10689_),
    .Y(_11044_));
 sky130_fd_sc_hd__or4_1 _20936_ (.A(_02229_),
    .B(_02240_),
    .C(_10687_),
    .D(_11040_),
    .X(_11045_));
 sky130_fd_sc_hd__a21oi_4 _20937_ (.A1(_11044_),
    .A2(_11042_),
    .B1(_11043_),
    .Y(_11046_));
 sky130_fd_sc_hd__o21bai_4 _20938_ (.A1(_11006_),
    .A2(_11008_),
    .B1_N(_11046_),
    .Y(_11048_));
 sky130_fd_sc_hd__and3_2 _20939_ (.A(_11007_),
    .B(_11046_),
    .C(_11009_),
    .X(_11049_));
 sky130_fd_sc_hd__nand3_4 _20940_ (.A(_11007_),
    .B(_11009_),
    .C(_11046_),
    .Y(_11050_));
 sky130_fd_sc_hd__o211a_1 _20941_ (.A1(_10531_),
    .A2(_10567_),
    .B1(_10831_),
    .C1(_10566_),
    .X(_11051_));
 sky130_fd_sc_hd__o2bb2a_1 _20942_ (.A1_N(_11048_),
    .A2_N(_11050_),
    .B1(_11051_),
    .B2(_10833_),
    .X(_11052_));
 sky130_fd_sc_hd__o2bb2ai_4 _20943_ (.A1_N(_11048_),
    .A2_N(_11050_),
    .B1(_11051_),
    .B2(_10833_),
    .Y(_11053_));
 sky130_fd_sc_hd__o21ai_2 _20944_ (.A1(_10830_),
    .A2(_10836_),
    .B1(_11048_),
    .Y(_11054_));
 sky130_fd_sc_hd__o211ai_4 _20945_ (.A1(_10830_),
    .A2(_10836_),
    .B1(_11048_),
    .C1(_11050_),
    .Y(_11055_));
 sky130_fd_sc_hd__inv_2 _20946_ (.A(_11055_),
    .Y(_11056_));
 sky130_fd_sc_hd__and3_1 _20947_ (.A(_10683_),
    .B(_10721_),
    .C(_10723_),
    .X(_11057_));
 sky130_fd_sc_hd__a31o_1 _20948_ (.A1(_10683_),
    .A2(_10721_),
    .A3(_10723_),
    .B1(_10681_),
    .X(_11059_));
 sky130_fd_sc_hd__a21boi_2 _20949_ (.A1(_11053_),
    .A2(_11055_),
    .B1_N(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__o2bb2ai_1 _20950_ (.A1_N(_11053_),
    .A2_N(_11055_),
    .B1(_11057_),
    .B2(_10681_),
    .Y(_11061_));
 sky130_fd_sc_hd__o221a_1 _20951_ (.A1(_10682_),
    .A2(_10725_),
    .B1(_11049_),
    .B2(_11054_),
    .C1(_11053_),
    .X(_11062_));
 sky130_fd_sc_hd__o221ai_4 _20952_ (.A1(_10682_),
    .A2(_10725_),
    .B1(_11049_),
    .B2(_11054_),
    .C1(_11053_),
    .Y(_11063_));
 sky130_fd_sc_hd__a22o_1 _20953_ (.A1(_10968_),
    .A2(_10972_),
    .B1(_11061_),
    .B2(_11063_),
    .X(_11064_));
 sky130_fd_sc_hd__o2111ai_1 _20954_ (.A1(_10963_),
    .A2(_10971_),
    .B1(_11061_),
    .C1(_11063_),
    .D1(_10968_),
    .Y(_11065_));
 sky130_fd_sc_hd__o221ai_2 _20955_ (.A1(_10971_),
    .A2(_10963_),
    .B1(_11062_),
    .B2(_11060_),
    .C1(_10968_),
    .Y(_11066_));
 sky130_fd_sc_hd__nand3_1 _20956_ (.A(_10973_),
    .B(_11061_),
    .C(_11063_),
    .Y(_11067_));
 sky130_fd_sc_hd__a31o_1 _20957_ (.A1(_10736_),
    .A2(_10737_),
    .A3(_10848_),
    .B1(_10845_),
    .X(_11068_));
 sky130_fd_sc_hd__a31oi_1 _20958_ (.A1(_10736_),
    .A2(_10737_),
    .A3(_10848_),
    .B1(_10845_),
    .Y(_11070_));
 sky130_fd_sc_hd__nand3_2 _20959_ (.A(_11066_),
    .B(_11067_),
    .C(_11070_),
    .Y(_11071_));
 sky130_fd_sc_hd__and3_1 _20960_ (.A(_11064_),
    .B(_11068_),
    .C(_11065_),
    .X(_11072_));
 sky130_fd_sc_hd__nand3_1 _20961_ (.A(_11064_),
    .B(_11068_),
    .C(_11065_),
    .Y(_11073_));
 sky130_fd_sc_hd__o211a_1 _20962_ (.A1(_10442_),
    .A2(_10405_),
    .B1(_10406_),
    .C1(_10733_),
    .X(_11074_));
 sky130_fd_sc_hd__o21ai_1 _20963_ (.A1(_10735_),
    .A2(_10732_),
    .B1(_10733_),
    .Y(_11075_));
 sky130_fd_sc_hd__o2bb2ai_2 _20964_ (.A1_N(_11071_),
    .A2_N(_11073_),
    .B1(_11074_),
    .B2(_10732_),
    .Y(_11076_));
 sky130_fd_sc_hd__nand2_1 _20965_ (.A(_11071_),
    .B(_11075_),
    .Y(_11077_));
 sky130_fd_sc_hd__nand3_1 _20966_ (.A(_11071_),
    .B(_11073_),
    .C(_11075_),
    .Y(_11078_));
 sky130_fd_sc_hd__o21ai_2 _20967_ (.A1(_10638_),
    .A2(_10856_),
    .B1(_10855_),
    .Y(_11079_));
 sky130_fd_sc_hd__a21oi_1 _20968_ (.A1(_11076_),
    .A2(_11078_),
    .B1(_11079_),
    .Y(_11081_));
 sky130_fd_sc_hd__a21o_1 _20969_ (.A1(_11076_),
    .A2(_11078_),
    .B1(_11079_),
    .X(_11082_));
 sky130_fd_sc_hd__o211a_1 _20970_ (.A1(_11072_),
    .A2(_11077_),
    .B1(_11079_),
    .C1(_11076_),
    .X(_11083_));
 sky130_fd_sc_hd__o211ai_1 _20971_ (.A1(_11072_),
    .A2(_11077_),
    .B1(_11079_),
    .C1(_11076_),
    .Y(_11084_));
 sky130_fd_sc_hd__a32o_1 _20972_ (.A1(_10684_),
    .A2(_10711_),
    .A3(_10713_),
    .B1(_10714_),
    .B2(_10425_),
    .X(_11085_));
 sky130_fd_sc_hd__o21bai_1 _20973_ (.A1(_11081_),
    .A2(_11083_),
    .B1_N(_11085_),
    .Y(_11086_));
 sky130_fd_sc_hd__nand3_1 _20974_ (.A(_11082_),
    .B(_11084_),
    .C(_11085_),
    .Y(_11087_));
 sky130_fd_sc_hd__o21ai_1 _20975_ (.A1(_11081_),
    .A2(_11083_),
    .B1(_11085_),
    .Y(_11088_));
 sky130_fd_sc_hd__nand3b_1 _20976_ (.A_N(_11085_),
    .B(_11084_),
    .C(_11082_),
    .Y(_11089_));
 sky130_fd_sc_hd__o2bb2ai_1 _20977_ (.A1_N(_10866_),
    .A2_N(_10863_),
    .B1(_10858_),
    .B2(_10864_),
    .Y(_11090_));
 sky130_fd_sc_hd__a21boi_1 _20978_ (.A1(_10863_),
    .A2(_10866_),
    .B1_N(_10865_),
    .Y(_11092_));
 sky130_fd_sc_hd__nand3_1 _20979_ (.A(_11088_),
    .B(_11089_),
    .C(_11092_),
    .Y(_11093_));
 sky130_fd_sc_hd__a21oi_1 _20980_ (.A1(_11088_),
    .A2(_11089_),
    .B1(_11092_),
    .Y(_11094_));
 sky130_fd_sc_hd__nand3_1 _20981_ (.A(_11086_),
    .B(_11087_),
    .C(_11090_),
    .Y(_11095_));
 sky130_fd_sc_hd__and2_1 _20982_ (.A(_11093_),
    .B(_11095_),
    .X(_11096_));
 sky130_fd_sc_hd__o221ai_2 _20983_ (.A1(_10629_),
    .A2(_10879_),
    .B1(_10878_),
    .B2(_10366_),
    .C1(_10876_),
    .Y(_11097_));
 sky130_fd_sc_hd__o311a_1 _20984_ (.A1(_10618_),
    .A2(_10625_),
    .A3(_10871_),
    .B1(_11096_),
    .C1(_11097_),
    .X(_11098_));
 sky130_fd_sc_hd__a21oi_1 _20985_ (.A1(_10875_),
    .A2(_11097_),
    .B1(_11096_),
    .Y(_11099_));
 sky130_fd_sc_hd__nor2_1 _20986_ (.A(_11098_),
    .B(_11099_),
    .Y(net106));
 sky130_fd_sc_hd__a31o_1 _20987_ (.A1(_11076_),
    .A2(_11079_),
    .A3(_11078_),
    .B1(_11085_),
    .X(_11100_));
 sky130_fd_sc_hd__a21o_1 _20988_ (.A1(_11071_),
    .A2(_11075_),
    .B1(_11072_),
    .X(_11102_));
 sky130_fd_sc_hd__o22a_1 _20989_ (.A1(_10681_),
    .A2(_11057_),
    .B1(_11049_),
    .B2(_11054_),
    .X(_11103_));
 sky130_fd_sc_hd__o311a_1 _20990_ (.A1(_10682_),
    .A2(_10720_),
    .A3(_10722_),
    .B1(_11053_),
    .C1(_10680_),
    .X(_11104_));
 sky130_fd_sc_hd__o31a_1 _20991_ (.A1(_10682_),
    .A2(_10725_),
    .A3(_11056_),
    .B1(_11053_),
    .X(_11105_));
 sky130_fd_sc_hd__o41a_1 _20992_ (.A1(_10813_),
    .A2(_10925_),
    .A3(_10941_),
    .A4(_10943_),
    .B1(_10950_),
    .X(_11106_));
 sky130_fd_sc_hd__o221ai_4 _20993_ (.A1(_10800_),
    .A2(_10801_),
    .B1(_10804_),
    .B2(_02218_),
    .C1(_10938_),
    .Y(_11107_));
 sky130_fd_sc_hd__a21o_1 _20994_ (.A1(_10935_),
    .A2(_10940_),
    .B1(_10936_),
    .X(_11108_));
 sky130_fd_sc_hd__a31o_1 _20995_ (.A1(_10929_),
    .A2(net24),
    .A3(net41),
    .B1(_10803_),
    .X(_11109_));
 sky130_fd_sc_hd__nor2_1 _20996_ (.A(_02010_),
    .B(_02251_),
    .Y(_11110_));
 sky130_fd_sc_hd__nand2_2 _20997_ (.A(net41),
    .B(net25),
    .Y(_11111_));
 sky130_fd_sc_hd__o2bb2ai_2 _20998_ (.A1_N(_10804_),
    .A2_N(_10929_),
    .B1(_02010_),
    .B2(_02251_),
    .Y(_11113_));
 sky130_fd_sc_hd__nand4_2 _20999_ (.A(_10929_),
    .B(net25),
    .C(net41),
    .D(_10804_),
    .Y(_11114_));
 sky130_fd_sc_hd__o21bai_1 _21000_ (.A1(_10803_),
    .A2(_10928_),
    .B1_N(_11111_),
    .Y(_11115_));
 sky130_fd_sc_hd__o211ai_1 _21001_ (.A1(_02010_),
    .A2(_02251_),
    .B1(_10804_),
    .C1(_10929_),
    .Y(_11116_));
 sky130_fd_sc_hd__nand3_4 _21002_ (.A(_10799_),
    .B(_11113_),
    .C(_11114_),
    .Y(_11117_));
 sky130_fd_sc_hd__a21oi_1 _21003_ (.A1(_11113_),
    .A2(_11114_),
    .B1(_10799_),
    .Y(_11118_));
 sky130_fd_sc_hd__nand3_2 _21004_ (.A(_11115_),
    .B(_11116_),
    .C(_10798_),
    .Y(_11119_));
 sky130_fd_sc_hd__o211a_1 _21005_ (.A1(_10803_),
    .A2(_10931_),
    .B1(_11117_),
    .C1(_11119_),
    .X(_11120_));
 sky130_fd_sc_hd__o211ai_4 _21006_ (.A1(_10803_),
    .A2(_10931_),
    .B1(_11117_),
    .C1(_11119_),
    .Y(_11121_));
 sky130_fd_sc_hd__a21oi_1 _21007_ (.A1(_11117_),
    .A2(_11119_),
    .B1(_11109_),
    .Y(_11122_));
 sky130_fd_sc_hd__a21o_1 _21008_ (.A1(_11117_),
    .A2(_11119_),
    .B1(_11109_),
    .X(_11124_));
 sky130_fd_sc_hd__nand3_4 _21009_ (.A(_11124_),
    .B(_11108_),
    .C(_11121_),
    .Y(_11125_));
 sky130_fd_sc_hd__o2bb2ai_2 _21010_ (.A1_N(_10935_),
    .A2_N(_11107_),
    .B1(_11120_),
    .B2(_11122_),
    .Y(_11126_));
 sky130_fd_sc_hd__nand2_1 _21011_ (.A(net48),
    .B(net18),
    .Y(_11127_));
 sky130_fd_sc_hd__nand4_2 _21012_ (.A(net46),
    .B(net47),
    .C(net19),
    .D(net20),
    .Y(_11128_));
 sky130_fd_sc_hd__a22oi_1 _21013_ (.A1(net47),
    .A2(net19),
    .B1(net20),
    .B2(net46),
    .Y(_11129_));
 sky130_fd_sc_hd__a22o_1 _21014_ (.A1(net47),
    .A2(net19),
    .B1(net20),
    .B2(net46),
    .X(_11130_));
 sky130_fd_sc_hd__nand4_1 _21015_ (.A(_11130_),
    .B(net18),
    .C(net48),
    .D(_11128_),
    .Y(_11131_));
 sky130_fd_sc_hd__o2bb2ai_1 _21016_ (.A1_N(_11128_),
    .A2_N(_11130_),
    .B1(_02109_),
    .B2(_02131_),
    .Y(_11132_));
 sky130_fd_sc_hd__and2_1 _21017_ (.A(_11131_),
    .B(_11132_),
    .X(_11133_));
 sky130_fd_sc_hd__nand2_1 _21018_ (.A(_11131_),
    .B(_11132_),
    .Y(_11135_));
 sky130_fd_sc_hd__a22oi_4 _21019_ (.A1(net43),
    .A2(net22),
    .B1(net24),
    .B2(net42),
    .Y(_11136_));
 sky130_fd_sc_hd__a22o_1 _21020_ (.A1(net43),
    .A2(net22),
    .B1(net24),
    .B2(net42),
    .X(_11137_));
 sky130_fd_sc_hd__and4_1 _21021_ (.A(net42),
    .B(net43),
    .C(net22),
    .D(net24),
    .X(_11138_));
 sky130_fd_sc_hd__nand4_1 _21022_ (.A(net42),
    .B(net43),
    .C(net22),
    .D(net24),
    .Y(_11139_));
 sky130_fd_sc_hd__o22ai_4 _21023_ (.A1(_02054_),
    .A2(_02185_),
    .B1(_11136_),
    .B2(_11138_),
    .Y(_11140_));
 sky130_fd_sc_hd__nand4_2 _21024_ (.A(_11137_),
    .B(_11139_),
    .C(net45),
    .D(net21),
    .Y(_11141_));
 sky130_fd_sc_hd__nand2_1 _21025_ (.A(_11140_),
    .B(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__o2bb2a_1 _21026_ (.A1_N(_10907_),
    .A2_N(_10910_),
    .B1(_10908_),
    .B2(_10766_),
    .X(_11143_));
 sky130_fd_sc_hd__o2bb2ai_1 _21027_ (.A1_N(_10907_),
    .A2_N(_10910_),
    .B1(_10908_),
    .B2(_10766_),
    .Y(_11144_));
 sky130_fd_sc_hd__o2bb2ai_1 _21028_ (.A1_N(_11140_),
    .A2_N(_11141_),
    .B1(_10766_),
    .B2(_10908_),
    .Y(_11146_));
 sky130_fd_sc_hd__a21o_1 _21029_ (.A1(_11140_),
    .A2(_11141_),
    .B1(_11144_),
    .X(_11147_));
 sky130_fd_sc_hd__and3_1 _21030_ (.A(_11140_),
    .B(_11141_),
    .C(_11144_),
    .X(_11148_));
 sky130_fd_sc_hd__nand3_1 _21031_ (.A(_11140_),
    .B(_11141_),
    .C(_11144_),
    .Y(_11149_));
 sky130_fd_sc_hd__a21oi_1 _21032_ (.A1(_11142_),
    .A2(_11143_),
    .B1(_11135_),
    .Y(_11150_));
 sky130_fd_sc_hd__o2bb2ai_1 _21033_ (.A1_N(_11135_),
    .A2_N(_11149_),
    .B1(_10911_),
    .B2(_11146_),
    .Y(_11151_));
 sky130_fd_sc_hd__a21oi_1 _21034_ (.A1(_11147_),
    .A2(_11149_),
    .B1(_11133_),
    .Y(_11152_));
 sky130_fd_sc_hd__and3_1 _21035_ (.A(_11147_),
    .B(_11149_),
    .C(_11133_),
    .X(_11153_));
 sky130_fd_sc_hd__a21oi_1 _21036_ (.A1(_11147_),
    .A2(_11149_),
    .B1(_11135_),
    .Y(_11154_));
 sky130_fd_sc_hd__and3_1 _21037_ (.A(_11135_),
    .B(_11147_),
    .C(_11149_),
    .X(_11155_));
 sky130_fd_sc_hd__o2bb2ai_4 _21038_ (.A1_N(_11125_),
    .A2_N(_11126_),
    .B1(_11152_),
    .B2(_11153_),
    .Y(_11157_));
 sky130_fd_sc_hd__o211ai_4 _21039_ (.A1(_11154_),
    .A2(_11155_),
    .B1(_11125_),
    .C1(_11126_),
    .Y(_11158_));
 sky130_fd_sc_hd__nand2_1 _21040_ (.A(_11157_),
    .B(_11158_),
    .Y(_11159_));
 sky130_fd_sc_hd__a21oi_2 _21041_ (.A1(_11157_),
    .A2(_11158_),
    .B1(_10894_),
    .Y(_11160_));
 sky130_fd_sc_hd__and3_1 _21042_ (.A(_10894_),
    .B(_11157_),
    .C(_11158_),
    .X(_11161_));
 sky130_fd_sc_hd__o211ai_4 _21043_ (.A1(_10481_),
    .A2(_10748_),
    .B1(_11157_),
    .C1(_11158_),
    .Y(_11162_));
 sky130_fd_sc_hd__o21ai_1 _21044_ (.A1(_11160_),
    .A2(_11161_),
    .B1(_11106_),
    .Y(_11163_));
 sky130_fd_sc_hd__o2bb2ai_2 _21045_ (.A1_N(_10892_),
    .A2_N(_11159_),
    .B1(_10949_),
    .B2(_10945_),
    .Y(_11164_));
 sky130_fd_sc_hd__o22ai_2 _21046_ (.A1(_10945_),
    .A2(_10949_),
    .B1(_11160_),
    .B2(_11161_),
    .Y(_11165_));
 sky130_fd_sc_hd__nand3b_1 _21047_ (.A_N(_11160_),
    .B(_11162_),
    .C(_11106_),
    .Y(_11166_));
 sky130_fd_sc_hd__o211ai_4 _21048_ (.A1(_10885_),
    .A2(_10887_),
    .B1(_11165_),
    .C1(_11166_),
    .Y(_11168_));
 sky130_fd_sc_hd__o211ai_4 _21049_ (.A1(_11161_),
    .A2(_11164_),
    .B1(_10889_),
    .C1(_11163_),
    .Y(_11169_));
 sky130_fd_sc_hd__nand2_1 _21050_ (.A(_11168_),
    .B(_11169_),
    .Y(_11170_));
 sky130_fd_sc_hd__nand3_2 _21051_ (.A(_10888_),
    .B(_10957_),
    .C(_10958_),
    .Y(_11171_));
 sky130_fd_sc_hd__o21ai_1 _21052_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_11171_),
    .Y(_11172_));
 sky130_fd_sc_hd__a22oi_2 _21053_ (.A1(_11168_),
    .A2(_11169_),
    .B1(_11171_),
    .B2(_10886_),
    .Y(_11173_));
 sky130_fd_sc_hd__a22o_2 _21054_ (.A1(_11168_),
    .A2(_11169_),
    .B1(_11171_),
    .B2(_10886_),
    .X(_11174_));
 sky130_fd_sc_hd__o2111a_1 _21055_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_11168_),
    .C1(_11169_),
    .D1(_11171_),
    .X(_11175_));
 sky130_fd_sc_hd__o2111ai_2 _21056_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_11168_),
    .C1(_11169_),
    .D1(_11171_),
    .Y(_11176_));
 sky130_fd_sc_hd__a21oi_2 _21057_ (.A1(_11007_),
    .A2(_11046_),
    .B1(_11008_),
    .Y(_11177_));
 sky130_fd_sc_hd__nand2_2 _21058_ (.A(_11000_),
    .B(_11004_),
    .Y(_11179_));
 sky130_fd_sc_hd__o31a_1 _21059_ (.A1(_10899_),
    .A2(_10901_),
    .A3(_10918_),
    .B1(_10917_),
    .X(_11180_));
 sky130_fd_sc_hd__o21ai_2 _21060_ (.A1(_10905_),
    .A2(_10918_),
    .B1(_10917_),
    .Y(_11181_));
 sky130_fd_sc_hd__nand2_2 _21061_ (.A(net17),
    .B(net50),
    .Y(_11182_));
 sky130_fd_sc_hd__nand2_1 _21062_ (.A(net17),
    .B(net49),
    .Y(_11183_));
 sky130_fd_sc_hd__and4_2 _21063_ (.A(net16),
    .B(net17),
    .C(net49),
    .D(net50),
    .X(_11184_));
 sky130_fd_sc_hd__a22o_1 _21064_ (.A1(net17),
    .A2(net49),
    .B1(net50),
    .B2(net16),
    .X(_11185_));
 sky130_fd_sc_hd__nand3_1 _21065_ (.A(_11183_),
    .B(net50),
    .C(net16),
    .Y(_11186_));
 sky130_fd_sc_hd__nand3_1 _21066_ (.A(_10976_),
    .B(net49),
    .C(net17),
    .Y(_11187_));
 sky130_fd_sc_hd__o2111a_1 _21067_ (.A1(_10977_),
    .A2(_11182_),
    .B1(net15),
    .C1(net51),
    .D1(_11185_),
    .X(_11188_));
 sky130_fd_sc_hd__o2111ai_4 _21068_ (.A1(_10977_),
    .A2(_11182_),
    .B1(net15),
    .C1(net51),
    .D1(_11185_),
    .Y(_11190_));
 sky130_fd_sc_hd__o211ai_2 _21069_ (.A1(_02076_),
    .A2(_02152_),
    .B1(_11186_),
    .C1(_11187_),
    .Y(_11191_));
 sky130_fd_sc_hd__o21ai_2 _21070_ (.A1(_10895_),
    .A2(_10897_),
    .B1(_10896_),
    .Y(_11192_));
 sky130_fd_sc_hd__nand3_2 _21071_ (.A(_11190_),
    .B(_11191_),
    .C(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__inv_2 _21072_ (.A(_11193_),
    .Y(_11194_));
 sky130_fd_sc_hd__a21oi_1 _21073_ (.A1(_11190_),
    .A2(_11191_),
    .B1(_11192_),
    .Y(_11195_));
 sky130_fd_sc_hd__a21o_1 _21074_ (.A1(_11190_),
    .A2(_11191_),
    .B1(_11192_),
    .X(_11196_));
 sky130_fd_sc_hd__o32a_1 _21075_ (.A1(_02076_),
    .A2(_02120_),
    .A3(_10976_),
    .B1(_02152_),
    .B2(_02065_),
    .X(_11197_));
 sky130_fd_sc_hd__a31o_1 _21076_ (.A1(_10982_),
    .A2(net51),
    .A3(net14),
    .B1(_10978_),
    .X(_11198_));
 sky130_fd_sc_hd__o2bb2ai_2 _21077_ (.A1_N(_11193_),
    .A2_N(_11196_),
    .B1(_11197_),
    .B2(_10980_),
    .Y(_11199_));
 sky130_fd_sc_hd__nand2_1 _21078_ (.A(_11193_),
    .B(_11198_),
    .Y(_11201_));
 sky130_fd_sc_hd__and3_2 _21079_ (.A(_11193_),
    .B(_11196_),
    .C(_11198_),
    .X(_11202_));
 sky130_fd_sc_hd__nand3_1 _21080_ (.A(_11193_),
    .B(_11196_),
    .C(_11198_),
    .Y(_11203_));
 sky130_fd_sc_hd__o21ai_1 _21081_ (.A1(_11195_),
    .A2(_11201_),
    .B1(_11199_),
    .Y(_11204_));
 sky130_fd_sc_hd__a21oi_2 _21082_ (.A1(_11199_),
    .A2(_11203_),
    .B1(_11181_),
    .Y(_11205_));
 sky130_fd_sc_hd__a21o_1 _21083_ (.A1(_11199_),
    .A2(_11203_),
    .B1(_11181_),
    .X(_11206_));
 sky130_fd_sc_hd__o21ai_2 _21084_ (.A1(_10916_),
    .A2(_10920_),
    .B1(_11199_),
    .Y(_11207_));
 sky130_fd_sc_hd__o211a_2 _21085_ (.A1(_11195_),
    .A2(_11201_),
    .B1(_11199_),
    .C1(_11181_),
    .X(_11208_));
 sky130_fd_sc_hd__nand2_1 _21086_ (.A(_10988_),
    .B(_10993_),
    .Y(_11209_));
 sky130_fd_sc_hd__o41a_2 _21087_ (.A1(_10777_),
    .A2(_10974_),
    .A3(_10983_),
    .A4(_10985_),
    .B1(_10993_),
    .X(_11210_));
 sky130_fd_sc_hd__o21ai_2 _21088_ (.A1(_11205_),
    .A2(_11208_),
    .B1(_11210_),
    .Y(_11212_));
 sky130_fd_sc_hd__a22oi_2 _21089_ (.A1(_10988_),
    .A2(_10993_),
    .B1(_11204_),
    .B2(_11180_),
    .Y(_11213_));
 sky130_fd_sc_hd__a22o_1 _21090_ (.A1(_10988_),
    .A2(_10993_),
    .B1(_11204_),
    .B2(_11180_),
    .X(_11214_));
 sky130_fd_sc_hd__o211ai_1 _21091_ (.A1(_11202_),
    .A2(_11207_),
    .B1(_11209_),
    .C1(_11206_),
    .Y(_11215_));
 sky130_fd_sc_hd__a21oi_1 _21092_ (.A1(_11212_),
    .A2(_11215_),
    .B1(_11179_),
    .Y(_11216_));
 sky130_fd_sc_hd__a21o_1 _21093_ (.A1(_11212_),
    .A2(_11215_),
    .B1(_11179_),
    .X(_11217_));
 sky130_fd_sc_hd__o211a_1 _21094_ (.A1(_11208_),
    .A2(_11214_),
    .B1(_11212_),
    .C1(_11179_),
    .X(_11218_));
 sky130_fd_sc_hd__o211ai_2 _21095_ (.A1(_11208_),
    .A2(_11214_),
    .B1(_11212_),
    .C1(_11179_),
    .Y(_11219_));
 sky130_fd_sc_hd__and4_2 _21096_ (.A(_01999_),
    .B(net10),
    .C(net56),
    .D(net57),
    .X(_11220_));
 sky130_fd_sc_hd__or4_1 _21097_ (.A(net9),
    .B(_02021_),
    .C(_02229_),
    .D(_02240_),
    .X(_11221_));
 sky130_fd_sc_hd__o22a_1 _21098_ (.A1(net9),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02021_),
    .X(_11223_));
 sky130_fd_sc_hd__nor2_1 _21099_ (.A(_11220_),
    .B(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__o21ai_1 _21100_ (.A1(_11016_),
    .A2(_11020_),
    .B1(_11018_),
    .Y(_11225_));
 sky130_fd_sc_hd__and2_1 _21101_ (.A(net11),
    .B(net54),
    .X(_11226_));
 sky130_fd_sc_hd__nand2_1 _21102_ (.A(net14),
    .B(net53),
    .Y(_11227_));
 sky130_fd_sc_hd__nand4_2 _21103_ (.A(net13),
    .B(net14),
    .C(net52),
    .D(net53),
    .Y(_11228_));
 sky130_fd_sc_hd__nand2_1 _21104_ (.A(net14),
    .B(net52),
    .Y(_11229_));
 sky130_fd_sc_hd__a22o_1 _21105_ (.A1(net14),
    .A2(net52),
    .B1(net53),
    .B2(net13),
    .X(_11230_));
 sky130_fd_sc_hd__a22oi_2 _21106_ (.A1(net11),
    .A2(net54),
    .B1(_11228_),
    .B2(_11230_),
    .Y(_11231_));
 sky130_fd_sc_hd__a22o_1 _21107_ (.A1(net11),
    .A2(net54),
    .B1(_11228_),
    .B2(_11230_),
    .X(_11232_));
 sky130_fd_sc_hd__o211a_1 _21108_ (.A1(_11019_),
    .A2(_11227_),
    .B1(_11226_),
    .C1(_11230_),
    .X(_11234_));
 sky130_fd_sc_hd__o2111ai_2 _21109_ (.A1(_11019_),
    .A2(_11227_),
    .B1(net11),
    .C1(net54),
    .D1(_11230_),
    .Y(_11235_));
 sky130_fd_sc_hd__o21bai_2 _21110_ (.A1(_11231_),
    .A2(_11234_),
    .B1_N(_11225_),
    .Y(_11236_));
 sky130_fd_sc_hd__a21o_1 _21111_ (.A1(_11018_),
    .A2(_11024_),
    .B1(_11231_),
    .X(_11237_));
 sky130_fd_sc_hd__nand3_1 _21112_ (.A(_11225_),
    .B(_11232_),
    .C(_11235_),
    .Y(_11238_));
 sky130_fd_sc_hd__o211ai_1 _21113_ (.A1(_11234_),
    .A2(_11237_),
    .B1(_11236_),
    .C1(_11224_),
    .Y(_11239_));
 sky130_fd_sc_hd__a2bb2o_1 _21114_ (.A1_N(_11220_),
    .A2_N(_11223_),
    .B1(_11236_),
    .B2(_11238_),
    .X(_11240_));
 sky130_fd_sc_hd__a21bo_1 _21115_ (.A1(_11236_),
    .A2(_11238_),
    .B1_N(_11224_),
    .X(_11241_));
 sky130_fd_sc_hd__o221ai_2 _21116_ (.A1(_11220_),
    .A2(_11223_),
    .B1(_11234_),
    .B2(_11237_),
    .C1(_11236_),
    .Y(_11242_));
 sky130_fd_sc_hd__nand4_2 _21117_ (.A(_11033_),
    .B(_11038_),
    .C(_11241_),
    .D(_11242_),
    .Y(_11243_));
 sky130_fd_sc_hd__inv_2 _21118_ (.A(_11243_),
    .Y(_11245_));
 sky130_fd_sc_hd__o211ai_2 _21119_ (.A1(_11032_),
    .A2(_11037_),
    .B1(_11239_),
    .C1(_11240_),
    .Y(_11246_));
 sky130_fd_sc_hd__nand3_1 _21120_ (.A(_11013_),
    .B(_11243_),
    .C(_11246_),
    .Y(_11247_));
 sky130_fd_sc_hd__a21o_1 _21121_ (.A1(_11243_),
    .A2(_11246_),
    .B1(_11013_),
    .X(_11248_));
 sky130_fd_sc_hd__nand2_2 _21122_ (.A(_11247_),
    .B(_11248_),
    .Y(_11249_));
 sky130_fd_sc_hd__o21bai_4 _21123_ (.A1(_11216_),
    .A2(_11218_),
    .B1_N(_11249_),
    .Y(_11250_));
 sky130_fd_sc_hd__nand3_4 _21124_ (.A(_11217_),
    .B(_11249_),
    .C(_11219_),
    .Y(_11251_));
 sky130_fd_sc_hd__nor2_1 _21125_ (.A(_10891_),
    .B(_10953_),
    .Y(_11252_));
 sky130_fd_sc_hd__a21o_1 _21126_ (.A1(_10956_),
    .A2(_10891_),
    .B1(_10953_),
    .X(_11253_));
 sky130_fd_sc_hd__a21oi_4 _21127_ (.A1(_11250_),
    .A2(_11251_),
    .B1(_11253_),
    .Y(_11254_));
 sky130_fd_sc_hd__o2bb2ai_1 _21128_ (.A1_N(_11250_),
    .A2_N(_11251_),
    .B1(_11252_),
    .B2(_10955_),
    .Y(_11256_));
 sky130_fd_sc_hd__o211a_1 _21129_ (.A1(_10953_),
    .A2(_10960_),
    .B1(_11250_),
    .C1(_11251_),
    .X(_11257_));
 sky130_fd_sc_hd__o211ai_4 _21130_ (.A1(_10953_),
    .A2(_10960_),
    .B1(_11250_),
    .C1(_11251_),
    .Y(_11258_));
 sky130_fd_sc_hd__o211ai_2 _21131_ (.A1(_11008_),
    .A2(_11049_),
    .B1(_11256_),
    .C1(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__o211a_1 _21132_ (.A1(_11254_),
    .A2(_11257_),
    .B1(_11009_),
    .C1(_11050_),
    .X(_11260_));
 sky130_fd_sc_hd__o21ai_1 _21133_ (.A1(_11254_),
    .A2(_11257_),
    .B1(_11177_),
    .Y(_11261_));
 sky130_fd_sc_hd__nand3_2 _21134_ (.A(_11256_),
    .B(_11258_),
    .C(_11177_),
    .Y(_11262_));
 sky130_fd_sc_hd__o22ai_4 _21135_ (.A1(_11008_),
    .A2(_11049_),
    .B1(_11254_),
    .B2(_11257_),
    .Y(_11263_));
 sky130_fd_sc_hd__o211ai_4 _21136_ (.A1(_11173_),
    .A2(_11175_),
    .B1(_11262_),
    .C1(_11263_),
    .Y(_11264_));
 sky130_fd_sc_hd__nand3_1 _21137_ (.A(_11174_),
    .B(_11176_),
    .C(_11259_),
    .Y(_11265_));
 sky130_fd_sc_hd__nand4_2 _21138_ (.A(_11174_),
    .B(_11176_),
    .C(_11259_),
    .D(_11261_),
    .Y(_11267_));
 sky130_fd_sc_hd__o22a_1 _21139_ (.A1(_10971_),
    .A2(_10963_),
    .B1(_11062_),
    .B2(_11060_),
    .X(_11268_));
 sky130_fd_sc_hd__nand2_1 _21140_ (.A(_10968_),
    .B(_11063_),
    .Y(_11269_));
 sky130_fd_sc_hd__o22ai_2 _21141_ (.A1(_10963_),
    .A2(_10971_),
    .B1(_11060_),
    .B2(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__o211a_1 _21142_ (.A1(_11260_),
    .A2(_11265_),
    .B1(_11264_),
    .C1(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__o211ai_1 _21143_ (.A1(_11260_),
    .A2(_11265_),
    .B1(_11264_),
    .C1(_11270_),
    .Y(_11272_));
 sky130_fd_sc_hd__a21oi_1 _21144_ (.A1(_11264_),
    .A2(_11267_),
    .B1(_11270_),
    .Y(_11273_));
 sky130_fd_sc_hd__o2bb2ai_2 _21145_ (.A1_N(_11264_),
    .A2_N(_11267_),
    .B1(_11268_),
    .B2(_10969_),
    .Y(_11274_));
 sky130_fd_sc_hd__o211a_1 _21146_ (.A1(_11056_),
    .A2(_11104_),
    .B1(_11272_),
    .C1(_11274_),
    .X(_11275_));
 sky130_fd_sc_hd__o211ai_1 _21147_ (.A1(_11056_),
    .A2(_11104_),
    .B1(_11272_),
    .C1(_11274_),
    .Y(_11276_));
 sky130_fd_sc_hd__o22a_1 _21148_ (.A1(_11052_),
    .A2(_11103_),
    .B1(_11271_),
    .B2(_11273_),
    .X(_00001_));
 sky130_fd_sc_hd__o22ai_1 _21149_ (.A1(_11052_),
    .A2(_11103_),
    .B1(_11271_),
    .B2(_11273_),
    .Y(_00002_));
 sky130_fd_sc_hd__a21oi_1 _21150_ (.A1(_11276_),
    .A2(_00002_),
    .B1(_11102_),
    .Y(_00003_));
 sky130_fd_sc_hd__o21bai_1 _21151_ (.A1(_11275_),
    .A2(_00001_),
    .B1_N(_11102_),
    .Y(_00004_));
 sky130_fd_sc_hd__nand3_1 _21152_ (.A(_11102_),
    .B(_11276_),
    .C(_00002_),
    .Y(_00005_));
 sky130_fd_sc_hd__o32a_1 _21153_ (.A1(_02229_),
    .A2(_02240_),
    .A3(_10687_),
    .B1(_11010_),
    .B2(_11039_),
    .X(_00006_));
 sky130_fd_sc_hd__a22oi_2 _21154_ (.A1(_11042_),
    .A2(_11045_),
    .B1(_00004_),
    .B2(_00005_),
    .Y(_00007_));
 sky130_fd_sc_hd__o211a_1 _21155_ (.A1(_11040_),
    .A2(_00006_),
    .B1(_00005_),
    .C1(_00004_),
    .X(_00008_));
 sky130_fd_sc_hd__a211o_1 _21156_ (.A1(_11082_),
    .A2(_11100_),
    .B1(_00007_),
    .C1(_00008_),
    .X(_00009_));
 sky130_fd_sc_hd__o211ai_2 _21157_ (.A1(_00007_),
    .A2(_00008_),
    .B1(_11082_),
    .C1(_11100_),
    .Y(_00010_));
 sky130_fd_sc_hd__nand2_2 _21158_ (.A(_00009_),
    .B(_00010_),
    .Y(_00012_));
 sky130_fd_sc_hd__o22ai_1 _21159_ (.A1(_10104_),
    .A2(_10364_),
    .B1(_10363_),
    .B2(_09836_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand4_1 _21160_ (.A(_10875_),
    .B(_10876_),
    .C(_11093_),
    .D(_11095_),
    .Y(_00014_));
 sky130_fd_sc_hd__nor2_1 _21161_ (.A(_10878_),
    .B(_00014_),
    .Y(_00015_));
 sky130_fd_sc_hd__a31oi_1 _21162_ (.A1(_11093_),
    .A2(_10871_),
    .A3(_10874_),
    .B1(_11094_),
    .Y(_00016_));
 sky130_fd_sc_hd__o21ai_2 _21163_ (.A1(_00014_),
    .A2(_10880_),
    .B1(_00016_),
    .Y(_00017_));
 sky130_fd_sc_hd__a21oi_1 _21164_ (.A1(_00015_),
    .A2(_00013_),
    .B1(_00017_),
    .Y(_00018_));
 sky130_fd_sc_hd__a21o_2 _21165_ (.A1(_00015_),
    .A2(_00013_),
    .B1(_00017_),
    .X(_00019_));
 sky130_fd_sc_hd__and4_2 _21166_ (.A(_09234_),
    .B(_09530_),
    .C(_10362_),
    .D(_00015_),
    .X(_00020_));
 sky130_fd_sc_hd__a41o_1 _21167_ (.A1(_09234_),
    .A2(_09530_),
    .A3(_10362_),
    .A4(_00015_),
    .B1(_00019_),
    .X(_00021_));
 sky130_fd_sc_hd__o211ai_4 _21168_ (.A1(_09238_),
    .A2(_07989_),
    .B1(_00018_),
    .C1(_09239_),
    .Y(_00023_));
 sky130_fd_sc_hd__o22ai_4 _21169_ (.A1(_00019_),
    .A2(_00020_),
    .B1(_00023_),
    .B2(_09243_),
    .Y(_00024_));
 sky130_fd_sc_hd__xor2_1 _21170_ (.A(_00012_),
    .B(_00024_),
    .X(net107));
 sky130_fd_sc_hd__and3_1 _21171_ (.A(_11009_),
    .B(_11050_),
    .C(_11258_),
    .X(_00025_));
 sky130_fd_sc_hd__o21ai_1 _21172_ (.A1(_11177_),
    .A2(_11254_),
    .B1(_11258_),
    .Y(_00026_));
 sky130_fd_sc_hd__o21a_1 _21173_ (.A1(_11177_),
    .A2(_11254_),
    .B1(_11258_),
    .X(_00027_));
 sky130_fd_sc_hd__o211ai_4 _21174_ (.A1(_11170_),
    .A2(_11172_),
    .B1(_11262_),
    .C1(_11263_),
    .Y(_00028_));
 sky130_fd_sc_hd__o21ai_1 _21175_ (.A1(_09386_),
    .A2(_10752_),
    .B1(_11169_),
    .Y(_00029_));
 sky130_fd_sc_hd__nand2_1 _21176_ (.A(_11125_),
    .B(_11158_),
    .Y(_00030_));
 sky130_fd_sc_hd__and2_1 _21177_ (.A(net45),
    .B(net22),
    .X(_00031_));
 sky130_fd_sc_hd__a22oi_1 _21178_ (.A1(net43),
    .A2(net24),
    .B1(net25),
    .B2(net42),
    .Y(_00033_));
 sky130_fd_sc_hd__a22o_1 _21179_ (.A1(net43),
    .A2(net24),
    .B1(net25),
    .B2(net42),
    .X(_00034_));
 sky130_fd_sc_hd__and3_1 _21180_ (.A(net42),
    .B(net43),
    .C(net25),
    .X(_00035_));
 sky130_fd_sc_hd__nand3_4 _21181_ (.A(net42),
    .B(net43),
    .C(net25),
    .Y(_00036_));
 sky130_fd_sc_hd__and4_1 _21182_ (.A(net42),
    .B(net43),
    .C(net24),
    .D(net25),
    .X(_00037_));
 sky130_fd_sc_hd__nand4_1 _21183_ (.A(net42),
    .B(net43),
    .C(net24),
    .D(net25),
    .Y(_00038_));
 sky130_fd_sc_hd__o22ai_2 _21184_ (.A1(_02054_),
    .A2(_02196_),
    .B1(_00033_),
    .B2(_00037_),
    .Y(_00039_));
 sky130_fd_sc_hd__nand3_2 _21185_ (.A(_00034_),
    .B(_00038_),
    .C(_00031_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _21186_ (.A(_00039_),
    .B(_00040_),
    .Y(_00041_));
 sky130_fd_sc_hd__o31a_1 _21187_ (.A1(_02054_),
    .A2(_02185_),
    .A3(_11136_),
    .B1(_11139_),
    .X(_00042_));
 sky130_fd_sc_hd__a31o_1 _21188_ (.A1(_11137_),
    .A2(net21),
    .A3(net45),
    .B1(_11138_),
    .X(_00044_));
 sky130_fd_sc_hd__and3_1 _21189_ (.A(_00039_),
    .B(_00040_),
    .C(_00044_),
    .X(_00045_));
 sky130_fd_sc_hd__nand3_1 _21190_ (.A(_00039_),
    .B(_00040_),
    .C(_00044_),
    .Y(_00046_));
 sky130_fd_sc_hd__nand2_2 _21191_ (.A(_00041_),
    .B(_00042_),
    .Y(_00047_));
 sky130_fd_sc_hd__inv_2 _21192_ (.A(_00047_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2_1 _21193_ (.A(net48),
    .B(net19),
    .Y(_00049_));
 sky130_fd_sc_hd__nand4_1 _21194_ (.A(net46),
    .B(net47),
    .C(net20),
    .D(net21),
    .Y(_00050_));
 sky130_fd_sc_hd__a22oi_1 _21195_ (.A1(net47),
    .A2(net20),
    .B1(net21),
    .B2(net46),
    .Y(_00051_));
 sky130_fd_sc_hd__a22o_1 _21196_ (.A1(net47),
    .A2(net20),
    .B1(net21),
    .B2(net46),
    .X(_00052_));
 sky130_fd_sc_hd__and4_1 _21197_ (.A(_00052_),
    .B(net19),
    .C(net48),
    .D(_00050_),
    .X(_00053_));
 sky130_fd_sc_hd__o2bb2a_1 _21198_ (.A1_N(_00050_),
    .A2_N(_00052_),
    .B1(_02109_),
    .B2(_02142_),
    .X(_00055_));
 sky130_fd_sc_hd__nor2_1 _21199_ (.A(_00053_),
    .B(_00055_),
    .Y(_00056_));
 sky130_fd_sc_hd__o2bb2ai_1 _21200_ (.A1_N(_00046_),
    .A2_N(_00047_),
    .B1(_00053_),
    .B2(_00055_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand3_1 _21201_ (.A(_00056_),
    .B(_00047_),
    .C(_00046_),
    .Y(_00058_));
 sky130_fd_sc_hd__o211ai_1 _21202_ (.A1(_11111_),
    .A2(_10928_),
    .B1(_10804_),
    .C1(_11119_),
    .Y(_00059_));
 sky130_fd_sc_hd__o211ai_1 _21203_ (.A1(net41),
    .A2(_10803_),
    .B1(_10929_),
    .C1(_11118_),
    .Y(_00060_));
 sky130_fd_sc_hd__nand3_1 _21204_ (.A(_11121_),
    .B(_00059_),
    .C(_00060_),
    .Y(_00061_));
 sky130_fd_sc_hd__a21o_1 _21205_ (.A1(_00057_),
    .A2(_00058_),
    .B1(_00061_),
    .X(_00062_));
 sky130_fd_sc_hd__nand3_2 _21206_ (.A(_00057_),
    .B(_00058_),
    .C(_00061_),
    .Y(_00063_));
 sky130_fd_sc_hd__a21oi_1 _21207_ (.A1(_00062_),
    .A2(_00063_),
    .B1(_10894_),
    .Y(_00064_));
 sky130_fd_sc_hd__a21o_1 _21208_ (.A1(_00062_),
    .A2(_00063_),
    .B1(_10894_),
    .X(_00066_));
 sky130_fd_sc_hd__o211a_1 _21209_ (.A1(_10481_),
    .A2(_10748_),
    .B1(_00062_),
    .C1(_00063_),
    .X(_00067_));
 sky130_fd_sc_hd__o211ai_1 _21210_ (.A1(_10481_),
    .A2(_10748_),
    .B1(_00062_),
    .C1(_00063_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand3b_2 _21211_ (.A_N(_00030_),
    .B(_00066_),
    .C(_00068_),
    .Y(_00069_));
 sky130_fd_sc_hd__o21ai_2 _21212_ (.A1(_00064_),
    .A2(_00067_),
    .B1(_00030_),
    .Y(_00070_));
 sky130_fd_sc_hd__o211a_1 _21213_ (.A1(_10885_),
    .A2(_10887_),
    .B1(_00069_),
    .C1(_00070_),
    .X(_00071_));
 sky130_fd_sc_hd__a21oi_4 _21214_ (.A1(_00069_),
    .A2(_00070_),
    .B1(_10890_),
    .Y(_00072_));
 sky130_fd_sc_hd__nor2_1 _21215_ (.A(_00071_),
    .B(_00072_),
    .Y(_00073_));
 sky130_fd_sc_hd__o221ai_4 _21216_ (.A1(_09386_),
    .A2(_10752_),
    .B1(_00071_),
    .B2(_00072_),
    .C1(_11169_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_2 _21217_ (.A(_00073_),
    .B(_00029_),
    .Y(_00075_));
 sky130_fd_sc_hd__nand2_1 _21218_ (.A(_00074_),
    .B(_00075_),
    .Y(_00077_));
 sky130_fd_sc_hd__a21o_1 _21219_ (.A1(_11217_),
    .A2(_11249_),
    .B1(_11218_),
    .X(_00078_));
 sky130_fd_sc_hd__o21ai_2 _21220_ (.A1(_11106_),
    .A2(_11160_),
    .B1(_11162_),
    .Y(_00079_));
 sky130_fd_sc_hd__o2bb2ai_1 _21221_ (.A1_N(_11224_),
    .A2_N(_11236_),
    .B1(_11237_),
    .B2(_11234_),
    .Y(_00080_));
 sky130_fd_sc_hd__and4_1 _21222_ (.A(_02021_),
    .B(net11),
    .C(net56),
    .D(net57),
    .X(_00081_));
 sky130_fd_sc_hd__or4_1 _21223_ (.A(net10),
    .B(_02032_),
    .C(_02229_),
    .D(_02240_),
    .X(_00082_));
 sky130_fd_sc_hd__o22a_1 _21224_ (.A1(net10),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02032_),
    .X(_00083_));
 sky130_fd_sc_hd__nor2_1 _21225_ (.A(_00081_),
    .B(_00083_),
    .Y(_00084_));
 sky130_fd_sc_hd__a21boi_1 _21226_ (.A1(_11230_),
    .A2(_11226_),
    .B1_N(_11228_),
    .Y(_00085_));
 sky130_fd_sc_hd__and2_1 _21227_ (.A(net13),
    .B(net54),
    .X(_00086_));
 sky130_fd_sc_hd__nand2_1 _21228_ (.A(net15),
    .B(net53),
    .Y(_00088_));
 sky130_fd_sc_hd__nand4_1 _21229_ (.A(net14),
    .B(net15),
    .C(net52),
    .D(net53),
    .Y(_00089_));
 sky130_fd_sc_hd__a22o_1 _21230_ (.A1(net15),
    .A2(net52),
    .B1(net53),
    .B2(net14),
    .X(_00090_));
 sky130_fd_sc_hd__a2bb2oi_1 _21231_ (.A1_N(_02043_),
    .A2_N(_02207_),
    .B1(_00089_),
    .B2(_00090_),
    .Y(_00091_));
 sky130_fd_sc_hd__o211a_1 _21232_ (.A1(_11229_),
    .A2(_00088_),
    .B1(_00086_),
    .C1(_00090_),
    .X(_00092_));
 sky130_fd_sc_hd__o21a_1 _21233_ (.A1(_00091_),
    .A2(_00092_),
    .B1(_00085_),
    .X(_00093_));
 sky130_fd_sc_hd__o21ai_1 _21234_ (.A1(_00091_),
    .A2(_00092_),
    .B1(_00085_),
    .Y(_00094_));
 sky130_fd_sc_hd__a211oi_1 _21235_ (.A1(_11228_),
    .A2(_11235_),
    .B1(_00091_),
    .C1(_00092_),
    .Y(_00095_));
 sky130_fd_sc_hd__a211o_1 _21236_ (.A1(_11228_),
    .A2(_11235_),
    .B1(_00091_),
    .C1(_00092_),
    .X(_00096_));
 sky130_fd_sc_hd__nand3_1 _21237_ (.A(_00096_),
    .B(_00084_),
    .C(_00094_),
    .Y(_00097_));
 sky130_fd_sc_hd__o22ai_1 _21238_ (.A1(_00081_),
    .A2(_00083_),
    .B1(_00093_),
    .B2(_00095_),
    .Y(_00099_));
 sky130_fd_sc_hd__o21ai_1 _21239_ (.A1(_00093_),
    .A2(_00095_),
    .B1(_00084_),
    .Y(_00100_));
 sky130_fd_sc_hd__o211ai_1 _21240_ (.A1(_00081_),
    .A2(_00083_),
    .B1(_00094_),
    .C1(_00096_),
    .Y(_00101_));
 sky130_fd_sc_hd__nand3b_2 _21241_ (.A_N(_00080_),
    .B(_00100_),
    .C(_00101_),
    .Y(_00102_));
 sky130_fd_sc_hd__nand3_2 _21242_ (.A(_00080_),
    .B(_00097_),
    .C(_00099_),
    .Y(_00103_));
 sky130_fd_sc_hd__a21o_1 _21243_ (.A1(_00102_),
    .A2(_00103_),
    .B1(_11220_),
    .X(_00104_));
 sky130_fd_sc_hd__nand3_2 _21244_ (.A(_00102_),
    .B(_00103_),
    .C(_11220_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand3_1 _21245_ (.A(_11221_),
    .B(_00102_),
    .C(_00103_),
    .Y(_00106_));
 sky130_fd_sc_hd__a21o_1 _21246_ (.A1(_00102_),
    .A2(_00103_),
    .B1(_11221_),
    .X(_00107_));
 sky130_fd_sc_hd__o22a_1 _21247_ (.A1(_11202_),
    .A2(_11207_),
    .B1(_11210_),
    .B2(_11205_),
    .X(_00108_));
 sky130_fd_sc_hd__o22ai_4 _21248_ (.A1(_11202_),
    .A2(_11207_),
    .B1(_11210_),
    .B2(_11205_),
    .Y(_00110_));
 sky130_fd_sc_hd__o21ai_1 _21249_ (.A1(_11195_),
    .A2(_11201_),
    .B1(_11193_),
    .Y(_00111_));
 sky130_fd_sc_hd__a31o_1 _21250_ (.A1(_11185_),
    .A2(net51),
    .A3(net15),
    .B1(_11184_),
    .X(_00112_));
 sky130_fd_sc_hd__o21ai_2 _21251_ (.A1(_11127_),
    .A2(_11129_),
    .B1(_11128_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_1 _21252_ (.A(net49),
    .B(net18),
    .Y(_00114_));
 sky130_fd_sc_hd__a22o_1 _21253_ (.A1(net49),
    .A2(net18),
    .B1(net50),
    .B2(net17),
    .X(_00115_));
 sky130_fd_sc_hd__nand4_1 _21254_ (.A(net17),
    .B(net49),
    .C(net18),
    .D(net50),
    .Y(_00116_));
 sky130_fd_sc_hd__nand3_1 _21255_ (.A(_00114_),
    .B(net50),
    .C(net17),
    .Y(_00117_));
 sky130_fd_sc_hd__nand3_1 _21256_ (.A(_11182_),
    .B(net18),
    .C(net49),
    .Y(_00118_));
 sky130_fd_sc_hd__o211ai_2 _21257_ (.A1(_02098_),
    .A2(_02152_),
    .B1(_00117_),
    .C1(_00118_),
    .Y(_00119_));
 sky130_fd_sc_hd__and4_2 _21258_ (.A(_00115_),
    .B(_00116_),
    .C(net16),
    .D(net51),
    .X(_00121_));
 sky130_fd_sc_hd__nand4_2 _21259_ (.A(_00115_),
    .B(_00116_),
    .C(net16),
    .D(net51),
    .Y(_00122_));
 sky130_fd_sc_hd__a21oi_1 _21260_ (.A1(_00119_),
    .A2(_00122_),
    .B1(_00113_),
    .Y(_00123_));
 sky130_fd_sc_hd__a21o_1 _21261_ (.A1(_00119_),
    .A2(_00122_),
    .B1(_00113_),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_1 _21262_ (.A(_00113_),
    .B(_00119_),
    .Y(_00125_));
 sky130_fd_sc_hd__and3_1 _21263_ (.A(_00113_),
    .B(_00119_),
    .C(_00122_),
    .X(_00126_));
 sky130_fd_sc_hd__nand3_1 _21264_ (.A(_00113_),
    .B(_00119_),
    .C(_00122_),
    .Y(_00127_));
 sky130_fd_sc_hd__o221a_1 _21265_ (.A1(_11184_),
    .A2(_11188_),
    .B1(_00121_),
    .B2(_00125_),
    .C1(_00124_),
    .X(_00128_));
 sky130_fd_sc_hd__o221ai_4 _21266_ (.A1(_11184_),
    .A2(_11188_),
    .B1(_00121_),
    .B2(_00125_),
    .C1(_00124_),
    .Y(_00129_));
 sky130_fd_sc_hd__o21bai_1 _21267_ (.A1(_00123_),
    .A2(_00126_),
    .B1_N(_00112_),
    .Y(_00130_));
 sky130_fd_sc_hd__o22ai_1 _21268_ (.A1(_11184_),
    .A2(_11188_),
    .B1(_00123_),
    .B2(_00126_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand3b_1 _21269_ (.A_N(_00112_),
    .B(_00124_),
    .C(_00127_),
    .Y(_00133_));
 sky130_fd_sc_hd__o211ai_4 _21270_ (.A1(_11148_),
    .A2(_11150_),
    .B1(_00129_),
    .C1(_00130_),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_2 _21271_ (.A(_00134_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand3_2 _21272_ (.A(_00132_),
    .B(_00133_),
    .C(_11151_),
    .Y(_00136_));
 sky130_fd_sc_hd__a21oi_1 _21273_ (.A1(_00134_),
    .A2(_00136_),
    .B1(_00111_),
    .Y(_00137_));
 sky130_fd_sc_hd__a21o_1 _21274_ (.A1(_00134_),
    .A2(_00136_),
    .B1(_00111_),
    .X(_00138_));
 sky130_fd_sc_hd__o211a_1 _21275_ (.A1(_11194_),
    .A2(_11202_),
    .B1(_00134_),
    .C1(_00136_),
    .X(_00139_));
 sky130_fd_sc_hd__o211ai_4 _21276_ (.A1(_11194_),
    .A2(_11202_),
    .B1(_00134_),
    .C1(_00136_),
    .Y(_00140_));
 sky130_fd_sc_hd__a21oi_1 _21277_ (.A1(_00138_),
    .A2(_00140_),
    .B1(_00110_),
    .Y(_00141_));
 sky130_fd_sc_hd__o21ai_4 _21278_ (.A1(_00137_),
    .A2(_00139_),
    .B1(_00108_),
    .Y(_00143_));
 sky130_fd_sc_hd__o211a_1 _21279_ (.A1(_11208_),
    .A2(_11213_),
    .B1(_00138_),
    .C1(_00140_),
    .X(_00144_));
 sky130_fd_sc_hd__o211ai_1 _21280_ (.A1(_11208_),
    .A2(_11213_),
    .B1(_00138_),
    .C1(_00140_),
    .Y(_00145_));
 sky130_fd_sc_hd__a32oi_4 _21281_ (.A1(_00110_),
    .A2(_00138_),
    .A3(_00140_),
    .B1(_00107_),
    .B2(_00106_),
    .Y(_00146_));
 sky130_fd_sc_hd__and4_1 _21282_ (.A(_00104_),
    .B(_00105_),
    .C(_00143_),
    .D(_00145_),
    .X(_00147_));
 sky130_fd_sc_hd__nand2_1 _21283_ (.A(_00146_),
    .B(_00143_),
    .Y(_00148_));
 sky130_fd_sc_hd__a22oi_2 _21284_ (.A1(_00104_),
    .A2(_00105_),
    .B1(_00143_),
    .B2(_00145_),
    .Y(_00149_));
 sky130_fd_sc_hd__o2bb2ai_2 _21285_ (.A1_N(_00104_),
    .A2_N(_00105_),
    .B1(_00141_),
    .B2(_00144_),
    .Y(_00150_));
 sky130_fd_sc_hd__a221oi_2 _21286_ (.A1(_00146_),
    .A2(_00143_),
    .B1(_11164_),
    .B2(_11162_),
    .C1(_00149_),
    .Y(_00151_));
 sky130_fd_sc_hd__a221o_1 _21287_ (.A1(_00146_),
    .A2(_00143_),
    .B1(_11164_),
    .B2(_11162_),
    .C1(_00149_),
    .X(_00152_));
 sky130_fd_sc_hd__a21oi_2 _21288_ (.A1(_00148_),
    .A2(_00150_),
    .B1(_00079_),
    .Y(_00154_));
 sky130_fd_sc_hd__a21o_1 _21289_ (.A1(_00148_),
    .A2(_00150_),
    .B1(_00079_),
    .X(_00155_));
 sky130_fd_sc_hd__nand3_2 _21290_ (.A(_00078_),
    .B(_00152_),
    .C(_00155_),
    .Y(_00156_));
 sky130_fd_sc_hd__o21bai_4 _21291_ (.A1(_00151_),
    .A2(_00154_),
    .B1_N(_00078_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand2_1 _21292_ (.A(_00156_),
    .B(_00157_),
    .Y(_00158_));
 sky130_fd_sc_hd__a22oi_2 _21293_ (.A1(_00074_),
    .A2(_00075_),
    .B1(_00156_),
    .B2(_00157_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand2_1 _21294_ (.A(_00077_),
    .B(_00158_),
    .Y(_00160_));
 sky130_fd_sc_hd__nand4_4 _21295_ (.A(_00074_),
    .B(_00075_),
    .C(_00156_),
    .D(_00157_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand3_2 _21296_ (.A(_11174_),
    .B(_00028_),
    .C(_00161_),
    .Y(_00162_));
 sky130_fd_sc_hd__a21oi_1 _21297_ (.A1(_00077_),
    .A2(_00158_),
    .B1(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__a21o_1 _21298_ (.A1(_00077_),
    .A2(_00158_),
    .B1(_00162_),
    .X(_00165_));
 sky130_fd_sc_hd__a22oi_4 _21299_ (.A1(_11174_),
    .A2(_00028_),
    .B1(_00160_),
    .B2(_00161_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand3b_1 _21300_ (.A_N(_00166_),
    .B(_00026_),
    .C(_00165_),
    .Y(_00167_));
 sky130_fd_sc_hd__o22ai_1 _21301_ (.A1(_11254_),
    .A2(_00025_),
    .B1(_00163_),
    .B2(_00166_),
    .Y(_00168_));
 sky130_fd_sc_hd__a221oi_2 _21302_ (.A1(_11174_),
    .A2(_00028_),
    .B1(_00160_),
    .B2(_00161_),
    .C1(_00026_),
    .Y(_00169_));
 sky130_fd_sc_hd__o22ai_4 _21303_ (.A1(_00159_),
    .A2(_00162_),
    .B1(_00027_),
    .B2(_00166_),
    .Y(_00170_));
 sky130_fd_sc_hd__a21oi_1 _21304_ (.A1(_11274_),
    .A2(_11105_),
    .B1(_11271_),
    .Y(_00171_));
 sky130_fd_sc_hd__a32o_1 _21305_ (.A1(_11264_),
    .A2(_11267_),
    .A3(_11270_),
    .B1(_11274_),
    .B2(_11105_),
    .X(_00172_));
 sky130_fd_sc_hd__o221ai_4 _21306_ (.A1(_00027_),
    .A2(_00165_),
    .B1(_00169_),
    .B2(_00170_),
    .C1(_00171_),
    .Y(_00173_));
 sky130_fd_sc_hd__nand3_1 _21307_ (.A(_00167_),
    .B(_00168_),
    .C(_00172_),
    .Y(_00174_));
 sky130_fd_sc_hd__o41a_1 _21308_ (.A1(net8),
    .A2(_01999_),
    .A3(_02229_),
    .A4(_02240_),
    .B1(_11246_),
    .X(_00176_));
 sky130_fd_sc_hd__a21oi_1 _21309_ (.A1(_11013_),
    .A2(_11246_),
    .B1(_11245_),
    .Y(_00177_));
 sky130_fd_sc_hd__a21boi_2 _21310_ (.A1(_00173_),
    .A2(_00177_),
    .B1_N(_00174_),
    .Y(_00178_));
 sky130_fd_sc_hd__o2bb2ai_1 _21311_ (.A1_N(_00173_),
    .A2_N(_00174_),
    .B1(_00176_),
    .B2(_11245_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand3_1 _21312_ (.A(_00173_),
    .B(_00174_),
    .C(_00177_),
    .Y(_00180_));
 sky130_fd_sc_hd__a31oi_1 _21313_ (.A1(_11042_),
    .A2(_11045_),
    .A3(_00005_),
    .B1(_00003_),
    .Y(_00181_));
 sky130_fd_sc_hd__a21oi_1 _21314_ (.A1(_00179_),
    .A2(_00180_),
    .B1(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand3_1 _21315_ (.A(_00181_),
    .B(_00180_),
    .C(_00179_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2b_1 _21316_ (.A_N(_00182_),
    .B(_00183_),
    .Y(_00184_));
 sky130_fd_sc_hd__o21ai_1 _21317_ (.A1(_00012_),
    .A2(_00024_),
    .B1(_00010_),
    .Y(_00185_));
 sky130_fd_sc_hd__xnor2_1 _21318_ (.A(_00184_),
    .B(_00185_),
    .Y(net108));
 sky130_fd_sc_hd__o211ai_1 _21319_ (.A1(_00029_),
    .A2(_00073_),
    .B1(_00156_),
    .C1(_00157_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _21320_ (.A(_00075_),
    .B(_00186_),
    .Y(_00187_));
 sky130_fd_sc_hd__and4_2 _21321_ (.A(_10119_),
    .B(_10470_),
    .C(_10928_),
    .D(_11111_),
    .X(_00188_));
 sky130_fd_sc_hd__o2111ai_4 _21322_ (.A1(_02010_),
    .A2(_02251_),
    .B1(_10119_),
    .C1(_10928_),
    .D1(_10470_),
    .Y(_00189_));
 sky130_fd_sc_hd__and3_2 _21323_ (.A(_10799_),
    .B(_10803_),
    .C(_11110_),
    .X(_00190_));
 sky130_fd_sc_hd__nand4_4 _21324_ (.A(_10799_),
    .B(_10803_),
    .C(net41),
    .D(net25),
    .Y(_00191_));
 sky130_fd_sc_hd__o31a_2 _21325_ (.A1(_11110_),
    .A2(_10929_),
    .A3(_10799_),
    .B1(_00191_),
    .X(_00192_));
 sky130_fd_sc_hd__o21ai_2 _21326_ (.A1(_10804_),
    .A2(_11117_),
    .B1(_00189_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _21327_ (.A(net48),
    .B(net20),
    .Y(_00194_));
 sky130_fd_sc_hd__nand4_2 _21328_ (.A(net46),
    .B(net47),
    .C(net21),
    .D(net22),
    .Y(_00196_));
 sky130_fd_sc_hd__a22oi_2 _21329_ (.A1(net47),
    .A2(net21),
    .B1(net22),
    .B2(net46),
    .Y(_00197_));
 sky130_fd_sc_hd__a22o_1 _21330_ (.A1(net47),
    .A2(net21),
    .B1(net22),
    .B2(net46),
    .X(_00198_));
 sky130_fd_sc_hd__nor3b_1 _21331_ (.A(_00197_),
    .B(_00194_),
    .C_N(_00196_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand4_1 _21332_ (.A(_00198_),
    .B(net20),
    .C(net48),
    .D(_00196_),
    .Y(_00200_));
 sky130_fd_sc_hd__a22oi_2 _21333_ (.A1(net48),
    .A2(net20),
    .B1(_00196_),
    .B2(_00198_),
    .Y(_00201_));
 sky130_fd_sc_hd__a22o_1 _21334_ (.A1(net48),
    .A2(net20),
    .B1(_00196_),
    .B2(_00198_),
    .X(_00202_));
 sky130_fd_sc_hd__nor2_1 _21335_ (.A(_00199_),
    .B(_00201_),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _21336_ (.A(_00200_),
    .B(_00202_),
    .Y(_00204_));
 sky130_fd_sc_hd__o21a_1 _21337_ (.A1(_02218_),
    .A2(_00036_),
    .B1(_00040_),
    .X(_00205_));
 sky130_fd_sc_hd__o21ai_1 _21338_ (.A1(_02218_),
    .A2(_00036_),
    .B1(_00040_),
    .Y(_00207_));
 sky130_fd_sc_hd__o21ai_2 _21339_ (.A1(net42),
    .A2(net43),
    .B1(net25),
    .Y(_00208_));
 sky130_fd_sc_hd__o21a_4 _21340_ (.A1(net42),
    .A2(net43),
    .B1(net25),
    .X(_00209_));
 sky130_fd_sc_hd__a22oi_1 _21341_ (.A1(net45),
    .A2(net24),
    .B1(_00036_),
    .B2(_00209_),
    .Y(_00210_));
 sky130_fd_sc_hd__o22ai_4 _21342_ (.A1(_02054_),
    .A2(_02218_),
    .B1(_00035_),
    .B2(_00208_),
    .Y(_00211_));
 sky130_fd_sc_hd__and4_1 _21343_ (.A(_00209_),
    .B(net24),
    .C(net45),
    .D(_00036_),
    .X(_00212_));
 sky130_fd_sc_hd__nand4_2 _21344_ (.A(_00209_),
    .B(net24),
    .C(net45),
    .D(_00036_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand3_1 _21345_ (.A(_00207_),
    .B(_00211_),
    .C(_00213_),
    .Y(_00214_));
 sky130_fd_sc_hd__a21oi_1 _21346_ (.A1(_00211_),
    .A2(_00213_),
    .B1(_00207_),
    .Y(_00215_));
 sky130_fd_sc_hd__o21ai_1 _21347_ (.A1(_00210_),
    .A2(_00212_),
    .B1(_00205_),
    .Y(_00216_));
 sky130_fd_sc_hd__a22o_1 _21348_ (.A1(_00038_),
    .A2(_00040_),
    .B1(_00211_),
    .B2(_00213_),
    .X(_00218_));
 sky130_fd_sc_hd__nand3_1 _21349_ (.A(_00205_),
    .B(_00211_),
    .C(_00213_),
    .Y(_00219_));
 sky130_fd_sc_hd__o211ai_2 _21350_ (.A1(_00199_),
    .A2(_00201_),
    .B1(_00218_),
    .C1(_00219_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand3_2 _21351_ (.A(_00216_),
    .B(_00203_),
    .C(_00214_),
    .Y(_00221_));
 sky130_fd_sc_hd__a21oi_1 _21352_ (.A1(_00220_),
    .A2(_00221_),
    .B1(_00192_),
    .Y(_00222_));
 sky130_fd_sc_hd__and3_1 _21353_ (.A(_00220_),
    .B(_00221_),
    .C(_00192_),
    .X(_00223_));
 sky130_fd_sc_hd__a21oi_1 _21354_ (.A1(_00220_),
    .A2(_00221_),
    .B1(_00193_),
    .Y(_00224_));
 sky130_fd_sc_hd__and3_1 _21355_ (.A(_00193_),
    .B(_00220_),
    .C(_00221_),
    .X(_00225_));
 sky130_fd_sc_hd__o21ai_2 _21356_ (.A1(_00224_),
    .A2(_00225_),
    .B1(_10894_),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _21357_ (.A(_00226_),
    .Y(_00227_));
 sky130_fd_sc_hd__o21ai_1 _21358_ (.A1(_00222_),
    .A2(_00223_),
    .B1(_10892_),
    .Y(_00229_));
 sky130_fd_sc_hd__o21ai_1 _21359_ (.A1(_10804_),
    .A2(_11117_),
    .B1(_00063_),
    .Y(_00230_));
 sky130_fd_sc_hd__a21o_1 _21360_ (.A1(_00226_),
    .A2(_00229_),
    .B1(_00230_),
    .X(_00231_));
 sky130_fd_sc_hd__and3_1 _21361_ (.A(_00226_),
    .B(_00229_),
    .C(_00230_),
    .X(_00232_));
 sky130_fd_sc_hd__nand3_2 _21362_ (.A(_00226_),
    .B(_00229_),
    .C(_00230_),
    .Y(_00233_));
 sky130_fd_sc_hd__a22o_1 _21363_ (.A1(_10886_),
    .A2(_10888_),
    .B1(_00231_),
    .B2(_00233_),
    .X(_00234_));
 sky130_fd_sc_hd__o2111ai_4 _21364_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .C1(_00231_),
    .D1(_00233_),
    .Y(_00235_));
 sky130_fd_sc_hd__o211ai_4 _21365_ (.A1(_10887_),
    .A2(_00072_),
    .B1(_00234_),
    .C1(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__a22o_1 _21366_ (.A1(_09385_),
    .A2(_10750_),
    .B1(_00234_),
    .B2(_00235_),
    .X(_00237_));
 sky130_fd_sc_hd__o21ai_1 _21367_ (.A1(_00072_),
    .A2(_00237_),
    .B1(_00236_),
    .Y(_00238_));
 sky130_fd_sc_hd__a31o_1 _21368_ (.A1(_00104_),
    .A2(_00105_),
    .A3(_00143_),
    .B1(_00144_),
    .X(_00240_));
 sky130_fd_sc_hd__a21o_1 _21369_ (.A1(_00030_),
    .A2(_00066_),
    .B1(_00067_),
    .X(_00241_));
 sky130_fd_sc_hd__a21o_1 _21370_ (.A1(_00084_),
    .A2(_00094_),
    .B1(_00095_),
    .X(_00242_));
 sky130_fd_sc_hd__and4_1 _21371_ (.A(_02032_),
    .B(net13),
    .C(net56),
    .D(net57),
    .X(_00243_));
 sky130_fd_sc_hd__or4_1 _21372_ (.A(net11),
    .B(_02043_),
    .C(_02229_),
    .D(_02240_),
    .X(_00244_));
 sky130_fd_sc_hd__o22a_1 _21373_ (.A1(net11),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02043_),
    .X(_00245_));
 sky130_fd_sc_hd__nor2_1 _21374_ (.A(_00243_),
    .B(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__o2bb2ai_1 _21375_ (.A1_N(_00086_),
    .A2_N(_00090_),
    .B1(_00088_),
    .B2(_11229_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand3_1 _21376_ (.A(net15),
    .B(net16),
    .C(net53),
    .Y(_00248_));
 sky130_fd_sc_hd__and4_1 _21377_ (.A(net15),
    .B(net16),
    .C(net52),
    .D(net53),
    .X(_00249_));
 sky130_fd_sc_hd__nand4_1 _21378_ (.A(net15),
    .B(net16),
    .C(net52),
    .D(net53),
    .Y(_00251_));
 sky130_fd_sc_hd__a22o_1 _21379_ (.A1(net16),
    .A2(net52),
    .B1(net53),
    .B2(net15),
    .X(_00252_));
 sky130_fd_sc_hd__a22oi_1 _21380_ (.A1(net14),
    .A2(net54),
    .B1(_00251_),
    .B2(_00252_),
    .Y(_00253_));
 sky130_fd_sc_hd__a22o_1 _21381_ (.A1(net14),
    .A2(net54),
    .B1(_00251_),
    .B2(_00252_),
    .X(_00254_));
 sky130_fd_sc_hd__o2111a_1 _21382_ (.A1(_02174_),
    .A2(_00248_),
    .B1(net54),
    .C1(net14),
    .D1(_00252_),
    .X(_00255_));
 sky130_fd_sc_hd__o2111ai_1 _21383_ (.A1(_02174_),
    .A2(_00248_),
    .B1(net54),
    .C1(net14),
    .D1(_00252_),
    .Y(_00256_));
 sky130_fd_sc_hd__o21bai_2 _21384_ (.A1(_00253_),
    .A2(_00255_),
    .B1_N(_00247_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand3_2 _21385_ (.A(_00247_),
    .B(_00254_),
    .C(_00256_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand3_1 _21386_ (.A(_00257_),
    .B(_00258_),
    .C(_00246_),
    .Y(_00259_));
 sky130_fd_sc_hd__a2bb2o_1 _21387_ (.A1_N(_00243_),
    .A2_N(_00245_),
    .B1(_00257_),
    .B2(_00258_),
    .X(_00260_));
 sky130_fd_sc_hd__a21bo_1 _21388_ (.A1(_00257_),
    .A2(_00258_),
    .B1_N(_00246_),
    .X(_00262_));
 sky130_fd_sc_hd__o211ai_1 _21389_ (.A1(_00243_),
    .A2(_00245_),
    .B1(_00257_),
    .C1(_00258_),
    .Y(_00263_));
 sky130_fd_sc_hd__a22o_1 _21390_ (.A1(_00096_),
    .A2(_00097_),
    .B1(_00262_),
    .B2(_00263_),
    .X(_00264_));
 sky130_fd_sc_hd__a21oi_2 _21391_ (.A1(_00259_),
    .A2(_00260_),
    .B1(_00242_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand4_1 _21392_ (.A(_00096_),
    .B(_00097_),
    .C(_00262_),
    .D(_00263_),
    .Y(_00266_));
 sky130_fd_sc_hd__nor2_1 _21393_ (.A(_00082_),
    .B(_00265_),
    .Y(_00267_));
 sky130_fd_sc_hd__a21oi_1 _21394_ (.A1(_00264_),
    .A2(_00266_),
    .B1(_00081_),
    .Y(_00268_));
 sky130_fd_sc_hd__and3_1 _21395_ (.A(_00082_),
    .B(_00264_),
    .C(_00266_),
    .X(_00269_));
 sky130_fd_sc_hd__a21oi_1 _21396_ (.A1(_00264_),
    .A2(_00266_),
    .B1(_00082_),
    .Y(_00270_));
 sky130_fd_sc_hd__a21oi_2 _21397_ (.A1(_00267_),
    .A2(_00264_),
    .B1(_00268_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _21398_ (.A(_00134_),
    .B(_00140_),
    .Y(_00273_));
 sky130_fd_sc_hd__o2bb2a_1 _21399_ (.A1_N(_00112_),
    .A2_N(_00124_),
    .B1(_00125_),
    .B2(_00121_),
    .X(_00274_));
 sky130_fd_sc_hd__o21ai_1 _21400_ (.A1(_00049_),
    .A2(_00051_),
    .B1(_00050_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _21401_ (.A(net49),
    .B(net19),
    .Y(_00276_));
 sky130_fd_sc_hd__a22oi_1 _21402_ (.A1(net18),
    .A2(net50),
    .B1(net19),
    .B2(net49),
    .Y(_00277_));
 sky130_fd_sc_hd__a22o_1 _21403_ (.A1(net18),
    .A2(net50),
    .B1(net19),
    .B2(net49),
    .X(_00278_));
 sky130_fd_sc_hd__nand2_1 _21404_ (.A(net50),
    .B(net19),
    .Y(_00279_));
 sky130_fd_sc_hd__and4_1 _21405_ (.A(net49),
    .B(net18),
    .C(net50),
    .D(net19),
    .X(_00280_));
 sky130_fd_sc_hd__o2111ai_4 _21406_ (.A1(_00114_),
    .A2(_00279_),
    .B1(net17),
    .C1(net51),
    .D1(_00278_),
    .Y(_00281_));
 sky130_fd_sc_hd__o2bb2ai_1 _21407_ (.A1_N(net17),
    .A2_N(net51),
    .B1(_00277_),
    .B2(_00280_),
    .Y(_00282_));
 sky130_fd_sc_hd__a21oi_2 _21408_ (.A1(_00281_),
    .A2(_00282_),
    .B1(_00275_),
    .Y(_00284_));
 sky130_fd_sc_hd__and3_1 _21409_ (.A(_00275_),
    .B(_00281_),
    .C(_00282_),
    .X(_00285_));
 sky130_fd_sc_hd__nand3_1 _21410_ (.A(_00275_),
    .B(_00281_),
    .C(_00282_),
    .Y(_00286_));
 sky130_fd_sc_hd__o31a_1 _21411_ (.A1(_02120_),
    .A2(_02131_),
    .A3(_11182_),
    .B1(_00122_),
    .X(_00287_));
 sky130_fd_sc_hd__a41o_1 _21412_ (.A1(net17),
    .A2(net49),
    .A3(net18),
    .A4(net50),
    .B1(_00121_),
    .X(_00288_));
 sky130_fd_sc_hd__o21ai_4 _21413_ (.A1(_00284_),
    .A2(_00285_),
    .B1(_00287_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand3b_2 _21414_ (.A_N(_00284_),
    .B(_00286_),
    .C(_00288_),
    .Y(_00290_));
 sky130_fd_sc_hd__a211oi_1 _21415_ (.A1(_00041_),
    .A2(_00042_),
    .B1(_00053_),
    .C1(_00055_),
    .Y(_00291_));
 sky130_fd_sc_hd__o22a_1 _21416_ (.A1(_00053_),
    .A2(_00055_),
    .B1(_00042_),
    .B2(_00041_),
    .X(_00292_));
 sky130_fd_sc_hd__a31o_1 _21417_ (.A1(_00039_),
    .A2(_00040_),
    .A3(_00044_),
    .B1(_00056_),
    .X(_00293_));
 sky130_fd_sc_hd__o211a_1 _21418_ (.A1(_00045_),
    .A2(_00291_),
    .B1(_00290_),
    .C1(_00289_),
    .X(_00295_));
 sky130_fd_sc_hd__o2111ai_4 _21419_ (.A1(_00045_),
    .A2(_00056_),
    .B1(_00289_),
    .C1(_00290_),
    .D1(_00047_),
    .Y(_00296_));
 sky130_fd_sc_hd__a22oi_2 _21420_ (.A1(_00289_),
    .A2(_00290_),
    .B1(_00293_),
    .B2(_00047_),
    .Y(_00297_));
 sky130_fd_sc_hd__o2bb2ai_1 _21421_ (.A1_N(_00289_),
    .A2_N(_00290_),
    .B1(_00292_),
    .B2(_00048_),
    .Y(_00298_));
 sky130_fd_sc_hd__o211a_1 _21422_ (.A1(_00126_),
    .A2(_00128_),
    .B1(_00296_),
    .C1(_00298_),
    .X(_00299_));
 sky130_fd_sc_hd__o211ai_2 _21423_ (.A1(_00126_),
    .A2(_00128_),
    .B1(_00296_),
    .C1(_00298_),
    .Y(_00300_));
 sky130_fd_sc_hd__a21boi_1 _21424_ (.A1(_00296_),
    .A2(_00298_),
    .B1_N(_00274_),
    .Y(_00301_));
 sky130_fd_sc_hd__o21ai_2 _21425_ (.A1(_00295_),
    .A2(_00297_),
    .B1(_00274_),
    .Y(_00302_));
 sky130_fd_sc_hd__o211a_2 _21426_ (.A1(_00135_),
    .A2(_00139_),
    .B1(_00300_),
    .C1(_00302_),
    .X(_00303_));
 sky130_fd_sc_hd__o211ai_1 _21427_ (.A1(_00135_),
    .A2(_00139_),
    .B1(_00300_),
    .C1(_00302_),
    .Y(_00304_));
 sky130_fd_sc_hd__a21oi_2 _21428_ (.A1(_00300_),
    .A2(_00302_),
    .B1(_00273_),
    .Y(_00306_));
 sky130_fd_sc_hd__o21bai_1 _21429_ (.A1(_00299_),
    .A2(_00301_),
    .B1_N(_00273_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _21430_ (.A(_00307_),
    .B(_00271_),
    .Y(_00308_));
 sky130_fd_sc_hd__o21bai_1 _21431_ (.A1(_00303_),
    .A2(_00306_),
    .B1_N(_00271_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand3b_1 _21432_ (.A_N(_00271_),
    .B(_00304_),
    .C(_00307_),
    .Y(_00310_));
 sky130_fd_sc_hd__o22ai_1 _21433_ (.A1(_00269_),
    .A2(_00270_),
    .B1(_00303_),
    .B2(_00306_),
    .Y(_00311_));
 sky130_fd_sc_hd__o211ai_4 _21434_ (.A1(_00303_),
    .A2(_00308_),
    .B1(_00241_),
    .C1(_00309_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand3b_2 _21435_ (.A_N(_00241_),
    .B(_00310_),
    .C(_00311_),
    .Y(_00313_));
 sky130_fd_sc_hd__o211a_1 _21436_ (.A1(_00144_),
    .A2(_00147_),
    .B1(_00312_),
    .C1(_00313_),
    .X(_00314_));
 sky130_fd_sc_hd__o211ai_2 _21437_ (.A1(_00144_),
    .A2(_00147_),
    .B1(_00312_),
    .C1(_00313_),
    .Y(_00315_));
 sky130_fd_sc_hd__a21oi_1 _21438_ (.A1(_00312_),
    .A2(_00313_),
    .B1(_00240_),
    .Y(_00317_));
 sky130_fd_sc_hd__a21o_1 _21439_ (.A1(_00312_),
    .A2(_00313_),
    .B1(_00240_),
    .X(_00318_));
 sky130_fd_sc_hd__o21ai_1 _21440_ (.A1(_00314_),
    .A2(_00317_),
    .B1(_00238_),
    .Y(_00319_));
 sky130_fd_sc_hd__o2111ai_4 _21441_ (.A1(_00237_),
    .A2(_00072_),
    .B1(_00236_),
    .C1(_00315_),
    .D1(_00318_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand3_2 _21442_ (.A(_00187_),
    .B(_00319_),
    .C(_00320_),
    .Y(_00321_));
 sky130_fd_sc_hd__a21o_2 _21443_ (.A1(_00319_),
    .A2(_00320_),
    .B1(_00187_),
    .X(_00322_));
 sky130_fd_sc_hd__and3_1 _21444_ (.A(_11219_),
    .B(_11251_),
    .C(_00152_),
    .X(_00323_));
 sky130_fd_sc_hd__a31o_1 _21445_ (.A1(_00079_),
    .A2(_00148_),
    .A3(_00150_),
    .B1(_00078_),
    .X(_00324_));
 sky130_fd_sc_hd__o21ai_2 _21446_ (.A1(_00154_),
    .A2(_00323_),
    .B1(_00321_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand4_2 _21447_ (.A(_00155_),
    .B(_00321_),
    .C(_00322_),
    .D(_00324_),
    .Y(_00326_));
 sky130_fd_sc_hd__o2bb2ai_1 _21448_ (.A1_N(_00321_),
    .A2_N(_00322_),
    .B1(_00323_),
    .B2(_00154_),
    .Y(_00328_));
 sky130_fd_sc_hd__a21oi_1 _21449_ (.A1(_00326_),
    .A2(_00328_),
    .B1(_00170_),
    .Y(_00329_));
 sky130_fd_sc_hd__a21o_1 _21450_ (.A1(_00326_),
    .A2(_00328_),
    .B1(_00170_),
    .X(_00330_));
 sky130_fd_sc_hd__nand3_2 _21451_ (.A(_00328_),
    .B(_00170_),
    .C(_00326_),
    .Y(_00331_));
 sky130_fd_sc_hd__a21bo_1 _21452_ (.A1(_11221_),
    .A2(_00103_),
    .B1_N(_00102_),
    .X(_00332_));
 sky130_fd_sc_hd__inv_2 _21453_ (.A(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__a21o_1 _21454_ (.A1(_00330_),
    .A2(_00331_),
    .B1(_00332_),
    .X(_00334_));
 sky130_fd_sc_hd__nand3_1 _21455_ (.A(_00330_),
    .B(_00331_),
    .C(_00332_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand3_1 _21456_ (.A(_00330_),
    .B(_00331_),
    .C(_00333_),
    .Y(_00336_));
 sky130_fd_sc_hd__a21o_1 _21457_ (.A1(_00330_),
    .A2(_00331_),
    .B1(_00333_),
    .X(_00337_));
 sky130_fd_sc_hd__nand3b_4 _21458_ (.A_N(_00178_),
    .B(_00336_),
    .C(_00337_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand3_2 _21459_ (.A(_00178_),
    .B(_00334_),
    .C(_00335_),
    .Y(_00340_));
 sky130_fd_sc_hd__o21a_1 _21460_ (.A1(_00182_),
    .A2(_00010_),
    .B1(_00183_),
    .X(_00341_));
 sky130_fd_sc_hd__o31a_1 _21461_ (.A1(_00012_),
    .A2(_00024_),
    .A3(_00184_),
    .B1(_00341_),
    .X(_00342_));
 sky130_fd_sc_hd__a21oi_1 _21462_ (.A1(_00339_),
    .A2(_00340_),
    .B1(_00342_),
    .Y(_00343_));
 sky130_fd_sc_hd__and3_1 _21463_ (.A(_00342_),
    .B(_00340_),
    .C(_00339_),
    .X(_00344_));
 sky130_fd_sc_hd__or2_1 _21464_ (.A(_00343_),
    .B(_00344_),
    .X(net110));
 sky130_fd_sc_hd__a31o_1 _21465_ (.A1(_00231_),
    .A2(_00233_),
    .A3(_10889_),
    .B1(_10887_),
    .X(_00345_));
 sky130_fd_sc_hd__a31o_1 _21466_ (.A1(_00189_),
    .A2(_00220_),
    .A3(_00221_),
    .B1(_00190_),
    .X(_00346_));
 sky130_fd_sc_hd__a22oi_2 _21467_ (.A1(net47),
    .A2(net22),
    .B1(net24),
    .B2(net46),
    .Y(_00347_));
 sky130_fd_sc_hd__a22o_1 _21468_ (.A1(net47),
    .A2(net22),
    .B1(net24),
    .B2(net46),
    .X(_00349_));
 sky130_fd_sc_hd__and4_1 _21469_ (.A(net46),
    .B(net47),
    .C(net22),
    .D(net24),
    .X(_00350_));
 sky130_fd_sc_hd__nand4_1 _21470_ (.A(net46),
    .B(net47),
    .C(net22),
    .D(net24),
    .Y(_00351_));
 sky130_fd_sc_hd__o211ai_2 _21471_ (.A1(_00347_),
    .A2(_00350_),
    .B1(net48),
    .C1(net21),
    .Y(_00352_));
 sky130_fd_sc_hd__o211ai_2 _21472_ (.A1(_02109_),
    .A2(_02185_),
    .B1(_00349_),
    .C1(_00351_),
    .Y(_00353_));
 sky130_fd_sc_hd__nand2_1 _21473_ (.A(_00352_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__o2111a_1 _21474_ (.A1(net42),
    .A2(net43),
    .B1(net45),
    .C1(net24),
    .D1(net25),
    .X(_00355_));
 sky130_fd_sc_hd__o31a_1 _21475_ (.A1(_02054_),
    .A2(_02218_),
    .A3(_00208_),
    .B1(_00036_),
    .X(_00356_));
 sky130_fd_sc_hd__nor2_2 _21476_ (.A(_02054_),
    .B(_02251_),
    .Y(_00357_));
 sky130_fd_sc_hd__o211ai_2 _21477_ (.A1(_02054_),
    .A2(_02251_),
    .B1(_00036_),
    .C1(_00209_),
    .Y(_00358_));
 sky130_fd_sc_hd__o21ai_1 _21478_ (.A1(_00035_),
    .A2(_00208_),
    .B1(_00357_),
    .Y(_00360_));
 sky130_fd_sc_hd__a22o_1 _21479_ (.A1(net45),
    .A2(net25),
    .B1(_00036_),
    .B2(_00209_),
    .X(_00361_));
 sky130_fd_sc_hd__nand4_1 _21480_ (.A(_00209_),
    .B(net25),
    .C(net45),
    .D(_00036_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand3_1 _21481_ (.A(_00356_),
    .B(_00361_),
    .C(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__o211ai_1 _21482_ (.A1(_00035_),
    .A2(_00355_),
    .B1(_00358_),
    .C1(_00360_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand3_2 _21483_ (.A(_00356_),
    .B(_00358_),
    .C(_00360_),
    .Y(_00365_));
 sky130_fd_sc_hd__and4_4 _21484_ (.A(net42),
    .B(net43),
    .C(net45),
    .D(net25),
    .X(_00366_));
 sky130_fd_sc_hd__nand4_4 _21485_ (.A(net42),
    .B(net43),
    .C(net45),
    .D(net25),
    .Y(_00367_));
 sky130_fd_sc_hd__o211ai_4 _21486_ (.A1(_02054_),
    .A2(_00036_),
    .B1(_00354_),
    .C1(_00365_),
    .Y(_00368_));
 sky130_fd_sc_hd__nand4_2 _21487_ (.A(_00352_),
    .B(_00353_),
    .C(_00363_),
    .D(_00364_),
    .Y(_00369_));
 sky130_fd_sc_hd__o211a_1 _21488_ (.A1(_00188_),
    .A2(_00190_),
    .B1(_00368_),
    .C1(_00369_),
    .X(_00371_));
 sky130_fd_sc_hd__a21oi_1 _21489_ (.A1(_00368_),
    .A2(_00369_),
    .B1(_00193_),
    .Y(_00372_));
 sky130_fd_sc_hd__a21o_1 _21490_ (.A1(_00368_),
    .A2(_00369_),
    .B1(_00193_),
    .X(_00373_));
 sky130_fd_sc_hd__o21ai_1 _21491_ (.A1(_00371_),
    .A2(_00372_),
    .B1(_10894_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand3b_2 _21492_ (.A_N(_00371_),
    .B(_00373_),
    .C(_10892_),
    .Y(_00375_));
 sky130_fd_sc_hd__inv_2 _21493_ (.A(_00375_),
    .Y(_00376_));
 sky130_fd_sc_hd__a21o_1 _21494_ (.A1(_00374_),
    .A2(_00375_),
    .B1(_00346_),
    .X(_00377_));
 sky130_fd_sc_hd__nand3_2 _21495_ (.A(_00346_),
    .B(_00374_),
    .C(_00375_),
    .Y(_00378_));
 sky130_fd_sc_hd__a22o_1 _21496_ (.A1(_10886_),
    .A2(_10888_),
    .B1(_00377_),
    .B2(_00378_),
    .X(_00379_));
 sky130_fd_sc_hd__o2111ai_2 _21497_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .C1(_00377_),
    .D1(_00378_),
    .Y(_00380_));
 sky130_fd_sc_hd__a21o_1 _21498_ (.A1(_00379_),
    .A2(_00380_),
    .B1(_00345_),
    .X(_00382_));
 sky130_fd_sc_hd__and3_1 _21499_ (.A(_00345_),
    .B(_00379_),
    .C(_00380_),
    .X(_00383_));
 sky130_fd_sc_hd__nand3_1 _21500_ (.A(_00345_),
    .B(_00379_),
    .C(_00380_),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_1 _21501_ (.A(_00382_),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__o31a_1 _21502_ (.A1(_10892_),
    .A2(_00222_),
    .A3(_00223_),
    .B1(_00233_),
    .X(_00386_));
 sky130_fd_sc_hd__o21ai_1 _21503_ (.A1(_00274_),
    .A2(_00297_),
    .B1(_00296_),
    .Y(_00387_));
 sky130_fd_sc_hd__o21ai_2 _21504_ (.A1(_00284_),
    .A2(_00287_),
    .B1(_00286_),
    .Y(_00388_));
 sky130_fd_sc_hd__o21ai_1 _21505_ (.A1(_00204_),
    .A2(_00215_),
    .B1(_00214_),
    .Y(_00389_));
 sky130_fd_sc_hd__a31o_1 _21506_ (.A1(_00278_),
    .A2(net51),
    .A3(net17),
    .B1(_00280_),
    .X(_00390_));
 sky130_fd_sc_hd__o21ai_2 _21507_ (.A1(_00194_),
    .A2(_00197_),
    .B1(_00196_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_2 _21508_ (.A(net49),
    .B(net20),
    .Y(_00393_));
 sky130_fd_sc_hd__a22o_1 _21509_ (.A1(net50),
    .A2(net19),
    .B1(net20),
    .B2(net49),
    .X(_00394_));
 sky130_fd_sc_hd__nand2_1 _21510_ (.A(net50),
    .B(net20),
    .Y(_00395_));
 sky130_fd_sc_hd__and4_1 _21511_ (.A(net49),
    .B(net50),
    .C(net19),
    .D(net20),
    .X(_00396_));
 sky130_fd_sc_hd__nand3_1 _21512_ (.A(_00393_),
    .B(net19),
    .C(net50),
    .Y(_00397_));
 sky130_fd_sc_hd__nand3_1 _21513_ (.A(_00279_),
    .B(net20),
    .C(net49),
    .Y(_00398_));
 sky130_fd_sc_hd__o2111a_1 _21514_ (.A1(_00276_),
    .A2(_00395_),
    .B1(net18),
    .C1(net51),
    .D1(_00394_),
    .X(_00399_));
 sky130_fd_sc_hd__o2111ai_4 _21515_ (.A1(_00276_),
    .A2(_00395_),
    .B1(net18),
    .C1(net51),
    .D1(_00394_),
    .Y(_00400_));
 sky130_fd_sc_hd__o211ai_2 _21516_ (.A1(_02131_),
    .A2(_02152_),
    .B1(_00397_),
    .C1(_00398_),
    .Y(_00401_));
 sky130_fd_sc_hd__a21o_1 _21517_ (.A1(_00400_),
    .A2(_00401_),
    .B1(_00391_),
    .X(_00402_));
 sky130_fd_sc_hd__nand2_1 _21518_ (.A(_00391_),
    .B(_00401_),
    .Y(_00404_));
 sky130_fd_sc_hd__and3_1 _21519_ (.A(_00391_),
    .B(_00400_),
    .C(_00401_),
    .X(_00405_));
 sky130_fd_sc_hd__nand3_1 _21520_ (.A(_00391_),
    .B(_00400_),
    .C(_00401_),
    .Y(_00406_));
 sky130_fd_sc_hd__o211a_2 _21521_ (.A1(_00404_),
    .A2(_00399_),
    .B1(_00390_),
    .C1(_00402_),
    .X(_00407_));
 sky130_fd_sc_hd__o211ai_1 _21522_ (.A1(_00404_),
    .A2(_00399_),
    .B1(_00390_),
    .C1(_00402_),
    .Y(_00408_));
 sky130_fd_sc_hd__a21oi_2 _21523_ (.A1(_00402_),
    .A2(_00406_),
    .B1(_00390_),
    .Y(_00409_));
 sky130_fd_sc_hd__a21o_1 _21524_ (.A1(_00402_),
    .A2(_00406_),
    .B1(_00390_),
    .X(_00410_));
 sky130_fd_sc_hd__o21bai_2 _21525_ (.A1(_00407_),
    .A2(_00409_),
    .B1_N(_00389_),
    .Y(_00411_));
 sky130_fd_sc_hd__a32o_1 _21526_ (.A1(_00390_),
    .A2(_00402_),
    .A3(_00406_),
    .B1(_00221_),
    .B2(_00214_),
    .X(_00412_));
 sky130_fd_sc_hd__nand3_1 _21527_ (.A(_00389_),
    .B(_00408_),
    .C(_00410_),
    .Y(_00413_));
 sky130_fd_sc_hd__a21o_1 _21528_ (.A1(_00411_),
    .A2(_00413_),
    .B1(_00388_),
    .X(_00415_));
 sky130_fd_sc_hd__o211ai_4 _21529_ (.A1(_00409_),
    .A2(_00412_),
    .B1(_00411_),
    .C1(_00388_),
    .Y(_00416_));
 sky130_fd_sc_hd__a21o_1 _21530_ (.A1(_00415_),
    .A2(_00416_),
    .B1(_00387_),
    .X(_00417_));
 sky130_fd_sc_hd__and3_1 _21531_ (.A(_00387_),
    .B(_00415_),
    .C(_00416_),
    .X(_00418_));
 sky130_fd_sc_hd__o211ai_4 _21532_ (.A1(_00295_),
    .A2(_00299_),
    .B1(_00415_),
    .C1(_00416_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _21533_ (.A(_00258_),
    .B(_00259_),
    .Y(_00420_));
 sky130_fd_sc_hd__and4_2 _21534_ (.A(_02043_),
    .B(net14),
    .C(net56),
    .D(net57),
    .X(_00421_));
 sky130_fd_sc_hd__o22a_1 _21535_ (.A1(net13),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02065_),
    .X(_00422_));
 sky130_fd_sc_hd__nor2_1 _21536_ (.A(_00421_),
    .B(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__a31o_1 _21537_ (.A1(_00252_),
    .A2(net54),
    .A3(net14),
    .B1(_00249_),
    .X(_00424_));
 sky130_fd_sc_hd__and4_1 _21538_ (.A(net16),
    .B(net17),
    .C(net52),
    .D(net53),
    .X(_00426_));
 sky130_fd_sc_hd__nand4_1 _21539_ (.A(net16),
    .B(net17),
    .C(net52),
    .D(net53),
    .Y(_00427_));
 sky130_fd_sc_hd__a22o_1 _21540_ (.A1(net17),
    .A2(net52),
    .B1(net53),
    .B2(net16),
    .X(_00428_));
 sky130_fd_sc_hd__a22o_1 _21541_ (.A1(net15),
    .A2(net54),
    .B1(_00427_),
    .B2(_00428_),
    .X(_00429_));
 sky130_fd_sc_hd__nand4_2 _21542_ (.A(_00428_),
    .B(net54),
    .C(net15),
    .D(_00427_),
    .Y(_00430_));
 sky130_fd_sc_hd__a21oi_1 _21543_ (.A1(_00429_),
    .A2(_00430_),
    .B1(_00424_),
    .Y(_00431_));
 sky130_fd_sc_hd__a21o_1 _21544_ (.A1(_00429_),
    .A2(_00430_),
    .B1(_00424_),
    .X(_00432_));
 sky130_fd_sc_hd__and3_1 _21545_ (.A(_00424_),
    .B(_00429_),
    .C(_00430_),
    .X(_00433_));
 sky130_fd_sc_hd__o211ai_2 _21546_ (.A1(_00249_),
    .A2(_00255_),
    .B1(_00429_),
    .C1(_00430_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand3_2 _21547_ (.A(_00434_),
    .B(_00423_),
    .C(_00432_),
    .Y(_00435_));
 sky130_fd_sc_hd__o22ai_2 _21548_ (.A1(_00421_),
    .A2(_00422_),
    .B1(_00431_),
    .B2(_00433_),
    .Y(_00437_));
 sky130_fd_sc_hd__a21o_1 _21549_ (.A1(_00435_),
    .A2(_00437_),
    .B1(_00420_),
    .X(_00438_));
 sky130_fd_sc_hd__nand3_1 _21550_ (.A(_00420_),
    .B(_00435_),
    .C(_00437_),
    .Y(_00439_));
 sky130_fd_sc_hd__a21oi_1 _21551_ (.A1(_00438_),
    .A2(_00439_),
    .B1(_00243_),
    .Y(_00440_));
 sky130_fd_sc_hd__and2_1 _21552_ (.A(_00438_),
    .B(_00243_),
    .X(_00441_));
 sky130_fd_sc_hd__and3_1 _21553_ (.A(_00438_),
    .B(_00439_),
    .C(_00243_),
    .X(_00442_));
 sky130_fd_sc_hd__and3_1 _21554_ (.A(_00244_),
    .B(_00438_),
    .C(_00439_),
    .X(_00443_));
 sky130_fd_sc_hd__a21oi_2 _21555_ (.A1(_00438_),
    .A2(_00439_),
    .B1(_00244_),
    .Y(_00444_));
 sky130_fd_sc_hd__o2bb2ai_1 _21556_ (.A1_N(_00417_),
    .A2_N(_00419_),
    .B1(_00440_),
    .B2(_00442_),
    .Y(_00445_));
 sky130_fd_sc_hd__o21ai_2 _21557_ (.A1(_00443_),
    .A2(_00444_),
    .B1(_00417_),
    .Y(_00446_));
 sky130_fd_sc_hd__o2bb2ai_1 _21558_ (.A1_N(_00417_),
    .A2_N(_00419_),
    .B1(_00443_),
    .B2(_00444_),
    .Y(_00448_));
 sky130_fd_sc_hd__o211ai_1 _21559_ (.A1(_00440_),
    .A2(_00442_),
    .B1(_00417_),
    .C1(_00419_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand3_1 _21560_ (.A(_00448_),
    .B(_00449_),
    .C(_00386_),
    .Y(_00450_));
 sky130_fd_sc_hd__o221ai_4 _21561_ (.A1(_00227_),
    .A2(_00232_),
    .B1(_00418_),
    .B2(_00446_),
    .C1(_00445_),
    .Y(_00451_));
 sky130_fd_sc_hd__nor2_1 _21562_ (.A(_00271_),
    .B(_00303_),
    .Y(_00452_));
 sky130_fd_sc_hd__o31a_1 _21563_ (.A1(_00269_),
    .A2(_00270_),
    .A3(_00303_),
    .B1(_00307_),
    .X(_00453_));
 sky130_fd_sc_hd__o2bb2ai_2 _21564_ (.A1_N(_00450_),
    .A2_N(_00451_),
    .B1(_00452_),
    .B2(_00306_),
    .Y(_00454_));
 sky130_fd_sc_hd__nand3_2 _21565_ (.A(_00450_),
    .B(_00451_),
    .C(_00453_),
    .Y(_00455_));
 sky130_fd_sc_hd__a21oi_1 _21566_ (.A1(_00454_),
    .A2(_00455_),
    .B1(_00385_),
    .Y(_00456_));
 sky130_fd_sc_hd__a21o_1 _21567_ (.A1(_00454_),
    .A2(_00455_),
    .B1(_00385_),
    .X(_00457_));
 sky130_fd_sc_hd__and3_1 _21568_ (.A(_00385_),
    .B(_00454_),
    .C(_00455_),
    .X(_00459_));
 sky130_fd_sc_hd__nand3_1 _21569_ (.A(_00385_),
    .B(_00454_),
    .C(_00455_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand4_2 _21570_ (.A(_00236_),
    .B(_00320_),
    .C(_00457_),
    .D(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__o2bb2ai_4 _21571_ (.A1_N(_00236_),
    .A2_N(_00320_),
    .B1(_00456_),
    .B2(_00459_),
    .Y(_00462_));
 sky130_fd_sc_hd__a21bo_1 _21572_ (.A1(_00240_),
    .A2(_00313_),
    .B1_N(_00312_),
    .X(_00463_));
 sky130_fd_sc_hd__a21oi_1 _21573_ (.A1(_00461_),
    .A2(_00462_),
    .B1(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__a21o_1 _21574_ (.A1(_00461_),
    .A2(_00462_),
    .B1(_00463_),
    .X(_00465_));
 sky130_fd_sc_hd__and3_1 _21575_ (.A(_00461_),
    .B(_00462_),
    .C(_00463_),
    .X(_00466_));
 sky130_fd_sc_hd__nand3_2 _21576_ (.A(_00461_),
    .B(_00462_),
    .C(_00463_),
    .Y(_00467_));
 sky130_fd_sc_hd__o211a_1 _21577_ (.A1(_00464_),
    .A2(_00466_),
    .B1(_00321_),
    .C1(_00326_),
    .X(_00468_));
 sky130_fd_sc_hd__o2bb2ai_2 _21578_ (.A1_N(_00322_),
    .A2_N(_00325_),
    .B1(_00464_),
    .B2(_00466_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand4_4 _21579_ (.A(_00322_),
    .B(_00325_),
    .C(_00465_),
    .D(_00467_),
    .Y(_00471_));
 sky130_fd_sc_hd__o41a_1 _21580_ (.A1(net10),
    .A2(_02032_),
    .A3(_02229_),
    .A4(_02240_),
    .B1(_00264_),
    .X(_00472_));
 sky130_fd_sc_hd__a31o_1 _21581_ (.A1(_00242_),
    .A2(_00259_),
    .A3(_00260_),
    .B1(_00267_),
    .X(_00473_));
 sky130_fd_sc_hd__o2bb2ai_2 _21582_ (.A1_N(_00470_),
    .A2_N(_00471_),
    .B1(_00472_),
    .B2(_00265_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand3_2 _21583_ (.A(_00470_),
    .B(_00471_),
    .C(_00473_),
    .Y(_00475_));
 sky130_fd_sc_hd__o21ai_2 _21584_ (.A1(_00329_),
    .A2(_00332_),
    .B1(_00331_),
    .Y(_00476_));
 sky130_fd_sc_hd__a21oi_2 _21585_ (.A1(_00474_),
    .A2(_00475_),
    .B1(_00476_),
    .Y(_00477_));
 sky130_fd_sc_hd__a21o_1 _21586_ (.A1(_00474_),
    .A2(_00475_),
    .B1(_00476_),
    .X(_00478_));
 sky130_fd_sc_hd__nand3_4 _21587_ (.A(_00476_),
    .B(_00475_),
    .C(_00474_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _21588_ (.A(_00478_),
    .B(_00479_),
    .Y(_00481_));
 sky130_fd_sc_hd__a32oi_2 _21589_ (.A1(_00178_),
    .A2(_00334_),
    .A3(_00335_),
    .B1(_00342_),
    .B2(_00339_),
    .Y(_00482_));
 sky130_fd_sc_hd__xnor2_1 _21590_ (.A(_00481_),
    .B(_00482_),
    .Y(net111));
 sky130_fd_sc_hd__o21a_1 _21591_ (.A1(_00265_),
    .A2(_00472_),
    .B1(_00471_),
    .X(_00483_));
 sky130_fd_sc_hd__nand2_1 _21592_ (.A(_00471_),
    .B(_00475_),
    .Y(_00484_));
 sky130_fd_sc_hd__o31a_1 _21593_ (.A1(_00265_),
    .A2(_00468_),
    .A3(_00472_),
    .B1(_00471_),
    .X(_00485_));
 sky130_fd_sc_hd__a31oi_1 _21594_ (.A1(_10886_),
    .A2(_00377_),
    .A3(_00378_),
    .B1(_10887_),
    .Y(_00486_));
 sky130_fd_sc_hd__a31o_1 _21595_ (.A1(_10886_),
    .A2(_00377_),
    .A3(_00378_),
    .B1(_10887_),
    .X(_00487_));
 sky130_fd_sc_hd__a31o_1 _21596_ (.A1(_00189_),
    .A2(_00368_),
    .A3(_00369_),
    .B1(_00190_),
    .X(_00488_));
 sky130_fd_sc_hd__o311a_2 _21597_ (.A1(net42),
    .A2(net43),
    .A3(net45),
    .B1(net25),
    .C1(_00367_),
    .X(_00489_));
 sky130_fd_sc_hd__nand2_1 _21598_ (.A(net48),
    .B(net22),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_2 _21599_ (.A(net46),
    .B(net25),
    .Y(_00492_));
 sky130_fd_sc_hd__and3_2 _21600_ (.A(net46),
    .B(net47),
    .C(net25),
    .X(_00493_));
 sky130_fd_sc_hd__nand3_4 _21601_ (.A(net46),
    .B(net47),
    .C(net25),
    .Y(_00494_));
 sky130_fd_sc_hd__nand4_1 _21602_ (.A(net46),
    .B(net47),
    .C(net24),
    .D(net25),
    .Y(_00495_));
 sky130_fd_sc_hd__a22oi_1 _21603_ (.A1(net47),
    .A2(net24),
    .B1(net25),
    .B2(net46),
    .Y(_00496_));
 sky130_fd_sc_hd__a22o_1 _21604_ (.A1(net47),
    .A2(net24),
    .B1(net25),
    .B2(net46),
    .X(_00497_));
 sky130_fd_sc_hd__o2111ai_4 _21605_ (.A1(_02218_),
    .A2(_00494_),
    .B1(net48),
    .C1(net22),
    .D1(_00497_),
    .Y(_00498_));
 sky130_fd_sc_hd__o2bb2ai_2 _21606_ (.A1_N(_00495_),
    .A2_N(_00497_),
    .B1(_02109_),
    .B2(_02196_),
    .Y(_00499_));
 sky130_fd_sc_hd__a21oi_1 _21607_ (.A1(_00498_),
    .A2(_00499_),
    .B1(_00489_),
    .Y(_00500_));
 sky130_fd_sc_hd__a21o_1 _21608_ (.A1(_00498_),
    .A2(_00499_),
    .B1(_00489_),
    .X(_00502_));
 sky130_fd_sc_hd__and3_1 _21609_ (.A(_00499_),
    .B(_00489_),
    .C(_00498_),
    .X(_00503_));
 sky130_fd_sc_hd__o2111ai_4 _21610_ (.A1(_00209_),
    .A2(_00357_),
    .B1(_00367_),
    .C1(_00498_),
    .D1(_00499_),
    .Y(_00504_));
 sky130_fd_sc_hd__and3_1 _21611_ (.A(_00192_),
    .B(_00502_),
    .C(_00504_),
    .X(_00505_));
 sky130_fd_sc_hd__o21ai_2 _21612_ (.A1(_00500_),
    .A2(_00503_),
    .B1(_00192_),
    .Y(_00506_));
 sky130_fd_sc_hd__o211ai_4 _21613_ (.A1(_00188_),
    .A2(_00190_),
    .B1(_00502_),
    .C1(_00504_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _21614_ (.A(_00506_),
    .B(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand4_2 _21615_ (.A(_10482_),
    .B(_10749_),
    .C(_00506_),
    .D(_00507_),
    .Y(_00509_));
 sky130_fd_sc_hd__a21oi_2 _21616_ (.A1(_00506_),
    .A2(_00507_),
    .B1(_10892_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _21617_ (.A(_10894_),
    .B(_00508_),
    .Y(_00511_));
 sky130_fd_sc_hd__a21o_1 _21618_ (.A1(_00509_),
    .A2(_00511_),
    .B1(_00488_),
    .X(_00513_));
 sky130_fd_sc_hd__nand3_4 _21619_ (.A(_00488_),
    .B(_00509_),
    .C(_00511_),
    .Y(_00514_));
 sky130_fd_sc_hd__inv_2 _21620_ (.A(_00514_),
    .Y(_00515_));
 sky130_fd_sc_hd__a21oi_1 _21621_ (.A1(_00513_),
    .A2(_00514_),
    .B1(_10889_),
    .Y(_00516_));
 sky130_fd_sc_hd__a22o_1 _21622_ (.A1(_10886_),
    .A2(_10888_),
    .B1(_00513_),
    .B2(_00514_),
    .X(_00517_));
 sky130_fd_sc_hd__o2111a_1 _21623_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .C1(_00513_),
    .D1(_00514_),
    .X(_00518_));
 sky130_fd_sc_hd__o2111ai_4 _21624_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .C1(_00513_),
    .D1(_00514_),
    .Y(_00519_));
 sky130_fd_sc_hd__and3_1 _21625_ (.A(_00487_),
    .B(_00517_),
    .C(_00519_),
    .X(_00520_));
 sky130_fd_sc_hd__nand3_1 _21626_ (.A(_00487_),
    .B(_00517_),
    .C(_00519_),
    .Y(_00521_));
 sky130_fd_sc_hd__o21ai_1 _21627_ (.A1(_00516_),
    .A2(_00518_),
    .B1(_00486_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_1 _21628_ (.A(_00521_),
    .B(_00522_),
    .Y(_00524_));
 sky130_fd_sc_hd__o2bb2a_1 _21629_ (.A1_N(_00388_),
    .A2_N(_00411_),
    .B1(_00412_),
    .B2(_00409_),
    .X(_00525_));
 sky130_fd_sc_hd__a2bb2o_1 _21630_ (.A1_N(_00412_),
    .A2_N(_00409_),
    .B1(_00388_),
    .B2(_00411_),
    .X(_00526_));
 sky130_fd_sc_hd__a31o_1 _21631_ (.A1(_00391_),
    .A2(_00400_),
    .A3(_00401_),
    .B1(_00407_),
    .X(_00527_));
 sky130_fd_sc_hd__a22o_1 _21632_ (.A1(net45),
    .A2(_00035_),
    .B1(_00365_),
    .B2(_00354_),
    .X(_00528_));
 sky130_fd_sc_hd__a31o_1 _21633_ (.A1(_00394_),
    .A2(net51),
    .A3(net18),
    .B1(_00396_),
    .X(_00529_));
 sky130_fd_sc_hd__nand2_2 _21634_ (.A(net50),
    .B(net21),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _21635_ (.A(net49),
    .B(net21),
    .Y(_00531_));
 sky130_fd_sc_hd__a22o_1 _21636_ (.A1(net50),
    .A2(net20),
    .B1(net21),
    .B2(net49),
    .X(_00532_));
 sky130_fd_sc_hd__nand3_1 _21637_ (.A(_00531_),
    .B(net20),
    .C(net50),
    .Y(_00533_));
 sky130_fd_sc_hd__nand3_1 _21638_ (.A(_00395_),
    .B(net21),
    .C(net49),
    .Y(_00535_));
 sky130_fd_sc_hd__o2111ai_4 _21639_ (.A1(_00393_),
    .A2(_00530_),
    .B1(net19),
    .C1(net51),
    .D1(_00532_),
    .Y(_00536_));
 sky130_fd_sc_hd__o211ai_2 _21640_ (.A1(_02142_),
    .A2(_02152_),
    .B1(_00533_),
    .C1(_00535_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _21641_ (.A(_00536_),
    .B(_00537_),
    .Y(_00538_));
 sky130_fd_sc_hd__o31a_1 _21642_ (.A1(_02109_),
    .A2(_02185_),
    .A3(_00347_),
    .B1(_00351_),
    .X(_00539_));
 sky130_fd_sc_hd__a31o_1 _21643_ (.A1(_00349_),
    .A2(net21),
    .A3(net48),
    .B1(_00350_),
    .X(_00540_));
 sky130_fd_sc_hd__nand3_2 _21644_ (.A(_00536_),
    .B(_00537_),
    .C(_00540_),
    .Y(_00541_));
 sky130_fd_sc_hd__inv_2 _21645_ (.A(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_2 _21646_ (.A(_00538_),
    .B(_00539_),
    .Y(_00543_));
 sky130_fd_sc_hd__a21oi_2 _21647_ (.A1(_00541_),
    .A2(_00543_),
    .B1(_00529_),
    .Y(_00544_));
 sky130_fd_sc_hd__a21o_1 _21648_ (.A1(_00541_),
    .A2(_00543_),
    .B1(_00529_),
    .X(_00546_));
 sky130_fd_sc_hd__o211a_2 _21649_ (.A1(_00396_),
    .A2(_00399_),
    .B1(_00541_),
    .C1(_00543_),
    .X(_00547_));
 sky130_fd_sc_hd__o211ai_2 _21650_ (.A1(_00396_),
    .A2(_00399_),
    .B1(_00541_),
    .C1(_00543_),
    .Y(_00548_));
 sky130_fd_sc_hd__o21bai_4 _21651_ (.A1(_00544_),
    .A2(_00547_),
    .B1_N(_00528_),
    .Y(_00549_));
 sky130_fd_sc_hd__a21oi_1 _21652_ (.A1(_00367_),
    .A2(_00368_),
    .B1(_00544_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _21653_ (.A(_00528_),
    .B(_00546_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand3_1 _21654_ (.A(_00528_),
    .B(_00546_),
    .C(_00548_),
    .Y(_00552_));
 sky130_fd_sc_hd__a21oi_1 _21655_ (.A1(_00549_),
    .A2(_00552_),
    .B1(_00527_),
    .Y(_00553_));
 sky130_fd_sc_hd__a21o_1 _21656_ (.A1(_00549_),
    .A2(_00552_),
    .B1(_00527_),
    .X(_00554_));
 sky130_fd_sc_hd__o221a_1 _21657_ (.A1(_00405_),
    .A2(_00407_),
    .B1(_00547_),
    .B2(_00551_),
    .C1(_00549_),
    .X(_00555_));
 sky130_fd_sc_hd__o221ai_4 _21658_ (.A1(_00405_),
    .A2(_00407_),
    .B1(_00547_),
    .B2(_00551_),
    .C1(_00549_),
    .Y(_00557_));
 sky130_fd_sc_hd__o21ai_2 _21659_ (.A1(_00553_),
    .A2(_00555_),
    .B1(_00525_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand3_4 _21660_ (.A(_00526_),
    .B(_00554_),
    .C(_00557_),
    .Y(_00559_));
 sky130_fd_sc_hd__a21o_1 _21661_ (.A1(_00432_),
    .A2(_00423_),
    .B1(_00433_),
    .X(_00560_));
 sky130_fd_sc_hd__nand2_1 _21662_ (.A(net15),
    .B(net56),
    .Y(_00561_));
 sky130_fd_sc_hd__and4_1 _21663_ (.A(_02065_),
    .B(net15),
    .C(net56),
    .D(net57),
    .X(_00562_));
 sky130_fd_sc_hd__or4_2 _21664_ (.A(net14),
    .B(_02076_),
    .C(_02229_),
    .D(_02240_),
    .X(_00563_));
 sky130_fd_sc_hd__o22a_1 _21665_ (.A1(net14),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02076_),
    .X(_00564_));
 sky130_fd_sc_hd__nor2_1 _21666_ (.A(_00562_),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__a31o_1 _21667_ (.A1(_00428_),
    .A2(net54),
    .A3(net15),
    .B1(_00426_),
    .X(_00566_));
 sky130_fd_sc_hd__nand4_2 _21668_ (.A(net17),
    .B(net18),
    .C(net52),
    .D(net53),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _21669_ (.A(net18),
    .B(net52),
    .Y(_00569_));
 sky130_fd_sc_hd__a22oi_1 _21670_ (.A1(net18),
    .A2(net52),
    .B1(net53),
    .B2(net17),
    .Y(_00570_));
 sky130_fd_sc_hd__a22o_1 _21671_ (.A1(net18),
    .A2(net52),
    .B1(net53),
    .B2(net17),
    .X(_00571_));
 sky130_fd_sc_hd__a22o_1 _21672_ (.A1(net16),
    .A2(net54),
    .B1(_00568_),
    .B2(_00571_),
    .X(_00572_));
 sky130_fd_sc_hd__nand4_2 _21673_ (.A(_00571_),
    .B(net54),
    .C(net16),
    .D(_00568_),
    .Y(_00573_));
 sky130_fd_sc_hd__a21o_1 _21674_ (.A1(_00572_),
    .A2(_00573_),
    .B1(_00566_),
    .X(_00574_));
 sky130_fd_sc_hd__nand3_4 _21675_ (.A(_00566_),
    .B(_00572_),
    .C(_00573_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand3_2 _21676_ (.A(_00574_),
    .B(_00575_),
    .C(_00565_),
    .Y(_00576_));
 sky130_fd_sc_hd__a2bb2o_1 _21677_ (.A1_N(_00562_),
    .A2_N(_00564_),
    .B1(_00574_),
    .B2(_00575_),
    .X(_00577_));
 sky130_fd_sc_hd__a21bo_1 _21678_ (.A1(_00574_),
    .A2(_00575_),
    .B1_N(_00565_),
    .X(_00579_));
 sky130_fd_sc_hd__o211ai_1 _21679_ (.A1(_00562_),
    .A2(_00564_),
    .B1(_00574_),
    .C1(_00575_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand4_2 _21680_ (.A(_00434_),
    .B(_00435_),
    .C(_00579_),
    .D(_00580_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand3_1 _21681_ (.A(_00560_),
    .B(_00576_),
    .C(_00577_),
    .Y(_00582_));
 sky130_fd_sc_hd__a21oi_1 _21682_ (.A1(_00581_),
    .A2(_00582_),
    .B1(_00421_),
    .Y(_00583_));
 sky130_fd_sc_hd__and3_1 _21683_ (.A(_00581_),
    .B(_00582_),
    .C(_00421_),
    .X(_00584_));
 sky130_fd_sc_hd__and3b_1 _21684_ (.A_N(_00421_),
    .B(_00581_),
    .C(_00582_),
    .X(_00585_));
 sky130_fd_sc_hd__a21boi_1 _21685_ (.A1(_00581_),
    .A2(_00582_),
    .B1_N(_00421_),
    .Y(_00586_));
 sky130_fd_sc_hd__o2bb2ai_2 _21686_ (.A1_N(_00558_),
    .A2_N(_00559_),
    .B1(_00583_),
    .B2(_00584_),
    .Y(_00587_));
 sky130_fd_sc_hd__o211ai_4 _21687_ (.A1(_00585_),
    .A2(_00586_),
    .B1(_00558_),
    .C1(_00559_),
    .Y(_00588_));
 sky130_fd_sc_hd__and2b_1 _21688_ (.A_N(_00346_),
    .B(_00374_),
    .X(_00590_));
 sky130_fd_sc_hd__nor2_1 _21689_ (.A(_00376_),
    .B(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__o2bb2a_1 _21690_ (.A1_N(_00587_),
    .A2_N(_00588_),
    .B1(_00590_),
    .B2(_00376_),
    .X(_00592_));
 sky130_fd_sc_hd__o2bb2ai_2 _21691_ (.A1_N(_00587_),
    .A2_N(_00588_),
    .B1(_00590_),
    .B2(_00376_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand3_2 _21692_ (.A(_00587_),
    .B(_00588_),
    .C(_00591_),
    .Y(_00594_));
 sky130_fd_sc_hd__o31a_1 _21693_ (.A1(_00418_),
    .A2(_00443_),
    .A3(_00444_),
    .B1(_00417_),
    .X(_00595_));
 sky130_fd_sc_hd__a21o_1 _21694_ (.A1(_00593_),
    .A2(_00594_),
    .B1(_00595_),
    .X(_00596_));
 sky130_fd_sc_hd__nand4_1 _21695_ (.A(_00419_),
    .B(_00446_),
    .C(_00593_),
    .D(_00594_),
    .Y(_00597_));
 sky130_fd_sc_hd__a22o_1 _21696_ (.A1(_00419_),
    .A2(_00446_),
    .B1(_00593_),
    .B2(_00594_),
    .X(_00598_));
 sky130_fd_sc_hd__nand3_2 _21697_ (.A(_00524_),
    .B(_00597_),
    .C(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__a31oi_4 _21698_ (.A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .B1(_00524_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_2 _21699_ (.A(_00601_),
    .B(_00596_),
    .Y(_00602_));
 sky130_fd_sc_hd__a31o_1 _21700_ (.A1(_00382_),
    .A2(_00454_),
    .A3(_00455_),
    .B1(_00383_),
    .X(_00603_));
 sky130_fd_sc_hd__a21oi_1 _21701_ (.A1(_00599_),
    .A2(_00602_),
    .B1(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__a21o_1 _21702_ (.A1(_00599_),
    .A2(_00602_),
    .B1(_00603_),
    .X(_00605_));
 sky130_fd_sc_hd__nand3_2 _21703_ (.A(_00603_),
    .B(_00602_),
    .C(_00599_),
    .Y(_00606_));
 sky130_fd_sc_hd__and2_1 _21704_ (.A(_00451_),
    .B(_00455_),
    .X(_00607_));
 sky130_fd_sc_hd__inv_2 _21705_ (.A(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__a22o_1 _21706_ (.A1(_00451_),
    .A2(_00455_),
    .B1(_00605_),
    .B2(_00606_),
    .X(_00609_));
 sky130_fd_sc_hd__nand4_1 _21707_ (.A(_00451_),
    .B(_00455_),
    .C(_00605_),
    .D(_00606_),
    .Y(_00610_));
 sky130_fd_sc_hd__a21o_1 _21708_ (.A1(_00605_),
    .A2(_00606_),
    .B1(_00608_),
    .X(_00612_));
 sky130_fd_sc_hd__nand3_1 _21709_ (.A(_00605_),
    .B(_00606_),
    .C(_00608_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _21710_ (.A(_00462_),
    .B(_00467_),
    .Y(_00614_));
 sky130_fd_sc_hd__and2_1 _21711_ (.A(_00462_),
    .B(_00467_),
    .X(_00615_));
 sky130_fd_sc_hd__and3_1 _21712_ (.A(_00609_),
    .B(_00610_),
    .C(_00615_),
    .X(_00616_));
 sky130_fd_sc_hd__nand4_2 _21713_ (.A(_00462_),
    .B(_00467_),
    .C(_00609_),
    .D(_00610_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand3_1 _21714_ (.A(_00614_),
    .B(_00613_),
    .C(_00612_),
    .Y(_00618_));
 sky130_fd_sc_hd__a31o_1 _21715_ (.A1(_00420_),
    .A2(_00435_),
    .A3(_00437_),
    .B1(_00441_),
    .X(_00619_));
 sky130_fd_sc_hd__and3_1 _21716_ (.A(_00617_),
    .B(_00618_),
    .C(_00619_),
    .X(_00620_));
 sky130_fd_sc_hd__nand3_1 _21717_ (.A(_00617_),
    .B(_00618_),
    .C(_00619_),
    .Y(_00621_));
 sky130_fd_sc_hd__a21oi_1 _21718_ (.A1(_00617_),
    .A2(_00618_),
    .B1(_00619_),
    .Y(_00623_));
 sky130_fd_sc_hd__a21o_1 _21719_ (.A1(_00617_),
    .A2(_00618_),
    .B1(_00619_),
    .X(_00624_));
 sky130_fd_sc_hd__nand2_1 _21720_ (.A(_00621_),
    .B(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand3_2 _21721_ (.A(_00484_),
    .B(_00621_),
    .C(_00624_),
    .Y(_00626_));
 sky130_fd_sc_hd__o22ai_1 _21722_ (.A1(_00468_),
    .A2(_00483_),
    .B1(_00620_),
    .B2(_00623_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand4_4 _21723_ (.A(_00339_),
    .B(_00340_),
    .C(_00478_),
    .D(_00479_),
    .Y(_00628_));
 sky130_fd_sc_hd__o221a_2 _21724_ (.A1(_00477_),
    .A2(_00339_),
    .B1(_00341_),
    .B2(_00628_),
    .C1(_00479_),
    .X(_00629_));
 sky130_fd_sc_hd__o221ai_4 _21725_ (.A1(_00477_),
    .A2(_00339_),
    .B1(_00341_),
    .B2(_00628_),
    .C1(_00479_),
    .Y(_00630_));
 sky130_fd_sc_hd__nor3_2 _21726_ (.A(_00012_),
    .B(_00184_),
    .C(_00628_),
    .Y(_00631_));
 sky130_fd_sc_hd__o211ai_4 _21727_ (.A1(_00023_),
    .A2(_09243_),
    .B1(_00631_),
    .C1(_00021_),
    .Y(_00632_));
 sky130_fd_sc_hd__a22oi_4 _21728_ (.A1(_00485_),
    .A2(_00625_),
    .B1(_00632_),
    .B2(_00629_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _21729_ (.A(_00626_),
    .B(_00627_),
    .Y(_00635_));
 sky130_fd_sc_hd__a32oi_4 _21730_ (.A1(_00629_),
    .A2(_00632_),
    .A3(_00635_),
    .B1(_00634_),
    .B2(_00626_),
    .Y(net112));
 sky130_fd_sc_hd__o21a_1 _21731_ (.A1(_00607_),
    .A2(_00604_),
    .B1(_00606_),
    .X(_00636_));
 sky130_fd_sc_hd__a32o_1 _21732_ (.A1(_00599_),
    .A2(_00602_),
    .A3(_00603_),
    .B1(_00605_),
    .B2(_00608_),
    .X(_00637_));
 sky130_fd_sc_hd__a21oi_1 _21733_ (.A1(_00601_),
    .A2(_00596_),
    .B1(_00520_),
    .Y(_00638_));
 sky130_fd_sc_hd__o31a_1 _21734_ (.A1(_08007_),
    .A2(_08962_),
    .A3(_10752_),
    .B1(_00519_),
    .X(_00639_));
 sky130_fd_sc_hd__a31o_1 _21735_ (.A1(_10799_),
    .A2(_10803_),
    .A3(_11110_),
    .B1(_00505_),
    .X(_00640_));
 sky130_fd_sc_hd__nand2_1 _21736_ (.A(net48),
    .B(net24),
    .Y(_00641_));
 sky130_fd_sc_hd__o21a_2 _21737_ (.A1(net46),
    .A2(net47),
    .B1(net25),
    .X(_00642_));
 sky130_fd_sc_hd__o21ai_4 _21738_ (.A1(net46),
    .A2(net47),
    .B1(net25),
    .Y(_00644_));
 sky130_fd_sc_hd__nor3_1 _21739_ (.A(_00641_),
    .B(_00644_),
    .C(_00493_),
    .Y(_00645_));
 sky130_fd_sc_hd__o2111ai_4 _21740_ (.A1(_02087_),
    .A2(_00492_),
    .B1(_00642_),
    .C1(net48),
    .D1(net24),
    .Y(_00646_));
 sky130_fd_sc_hd__o22a_1 _21741_ (.A1(_02109_),
    .A2(_02218_),
    .B1(_00644_),
    .B2(_00493_),
    .X(_00647_));
 sky130_fd_sc_hd__a22o_1 _21742_ (.A1(net48),
    .A2(net24),
    .B1(_00642_),
    .B2(_00494_),
    .X(_00648_));
 sky130_fd_sc_hd__and3_1 _21743_ (.A(_00648_),
    .B(_00489_),
    .C(_00646_),
    .X(_00649_));
 sky130_fd_sc_hd__o2111ai_2 _21744_ (.A1(_00209_),
    .A2(_00357_),
    .B1(_00367_),
    .C1(_00646_),
    .D1(_00648_),
    .Y(_00650_));
 sky130_fd_sc_hd__o21bai_1 _21745_ (.A1(_00645_),
    .A2(_00647_),
    .B1_N(_00489_),
    .Y(_00651_));
 sky130_fd_sc_hd__nand4_2 _21746_ (.A(_00189_),
    .B(_00191_),
    .C(_00650_),
    .D(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__a22o_1 _21747_ (.A1(_00189_),
    .A2(_00191_),
    .B1(_00650_),
    .B2(_00651_),
    .X(_00653_));
 sky130_fd_sc_hd__nand2_1 _21748_ (.A(_00652_),
    .B(_00653_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand2_1 _21749_ (.A(_00655_),
    .B(_10892_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand3_2 _21750_ (.A(_10894_),
    .B(_00652_),
    .C(_00653_),
    .Y(_00657_));
 sky130_fd_sc_hd__a21oi_2 _21751_ (.A1(_00656_),
    .A2(_00657_),
    .B1(_00640_),
    .Y(_00658_));
 sky130_fd_sc_hd__a21o_1 _21752_ (.A1(_00656_),
    .A2(_00657_),
    .B1(_00640_),
    .X(_00659_));
 sky130_fd_sc_hd__and3_1 _21753_ (.A(_00640_),
    .B(_00656_),
    .C(_00657_),
    .X(_00660_));
 sky130_fd_sc_hd__o211ai_2 _21754_ (.A1(_00190_),
    .A2(_00505_),
    .B1(_00656_),
    .C1(_00657_),
    .Y(_00661_));
 sky130_fd_sc_hd__o22ai_4 _21755_ (.A1(_10885_),
    .A2(_10887_),
    .B1(_00658_),
    .B2(_00660_),
    .Y(_00662_));
 sky130_fd_sc_hd__o2111ai_4 _21756_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .C1(_00659_),
    .D1(_00661_),
    .Y(_00663_));
 sky130_fd_sc_hd__nand2_1 _21757_ (.A(_00662_),
    .B(_00663_),
    .Y(_00664_));
 sky130_fd_sc_hd__a21o_1 _21758_ (.A1(_10888_),
    .A2(_00519_),
    .B1(_00664_),
    .X(_00666_));
 sky130_fd_sc_hd__a22oi_4 _21759_ (.A1(_10888_),
    .A2(_00519_),
    .B1(_00662_),
    .B2(_00663_),
    .Y(_00667_));
 sky130_fd_sc_hd__and4_1 _21760_ (.A(_10888_),
    .B(_00519_),
    .C(_00662_),
    .D(_00663_),
    .X(_00668_));
 sky130_fd_sc_hd__nor2_1 _21761_ (.A(_00667_),
    .B(_00668_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand2_1 _21762_ (.A(_00559_),
    .B(_00588_),
    .Y(_00670_));
 sky130_fd_sc_hd__a21oi_1 _21763_ (.A1(_00488_),
    .A2(_00509_),
    .B1(_00510_),
    .Y(_00671_));
 sky130_fd_sc_hd__a22oi_2 _21764_ (.A1(_00548_),
    .A2(_00550_),
    .B1(_00549_),
    .B2(_00527_),
    .Y(_00672_));
 sky130_fd_sc_hd__o2bb2ai_1 _21765_ (.A1_N(_00527_),
    .A2_N(_00549_),
    .B1(_00551_),
    .B2(_00547_),
    .Y(_00673_));
 sky130_fd_sc_hd__a32oi_1 _21766_ (.A1(_00536_),
    .A2(_00537_),
    .A3(_00540_),
    .B1(_00543_),
    .B2(_00529_),
    .Y(_00674_));
 sky130_fd_sc_hd__o21a_1 _21767_ (.A1(_02054_),
    .A2(_00036_),
    .B1(_00504_),
    .X(_00675_));
 sky130_fd_sc_hd__o31a_1 _21768_ (.A1(_02120_),
    .A2(_02163_),
    .A3(_00530_),
    .B1(_00536_),
    .X(_00677_));
 sky130_fd_sc_hd__o21ai_1 _21769_ (.A1(_00393_),
    .A2(_00530_),
    .B1(_00536_),
    .Y(_00678_));
 sky130_fd_sc_hd__o21ai_1 _21770_ (.A1(_00491_),
    .A2(_00496_),
    .B1(_00495_),
    .Y(_00679_));
 sky130_fd_sc_hd__nand2_1 _21771_ (.A(net50),
    .B(net22),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _21772_ (.A(net49),
    .B(net22),
    .Y(_00681_));
 sky130_fd_sc_hd__nand4_1 _21773_ (.A(net49),
    .B(net50),
    .C(net21),
    .D(net22),
    .Y(_00682_));
 sky130_fd_sc_hd__a22o_1 _21774_ (.A1(net50),
    .A2(net21),
    .B1(net22),
    .B2(net49),
    .X(_00683_));
 sky130_fd_sc_hd__nand3_1 _21775_ (.A(_00681_),
    .B(net21),
    .C(net50),
    .Y(_00684_));
 sky130_fd_sc_hd__nand3_1 _21776_ (.A(_00530_),
    .B(net22),
    .C(net49),
    .Y(_00685_));
 sky130_fd_sc_hd__o211ai_2 _21777_ (.A1(_02152_),
    .A2(_02163_),
    .B1(_00684_),
    .C1(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand4_2 _21778_ (.A(_00683_),
    .B(net20),
    .C(net51),
    .D(_00682_),
    .Y(_00688_));
 sky130_fd_sc_hd__a21oi_1 _21779_ (.A1(_00686_),
    .A2(_00688_),
    .B1(_00679_),
    .Y(_00689_));
 sky130_fd_sc_hd__a21o_1 _21780_ (.A1(_00686_),
    .A2(_00688_),
    .B1(_00679_),
    .X(_00690_));
 sky130_fd_sc_hd__and3_1 _21781_ (.A(_00679_),
    .B(_00686_),
    .C(_00688_),
    .X(_00691_));
 sky130_fd_sc_hd__nand3_1 _21782_ (.A(_00679_),
    .B(_00686_),
    .C(_00688_),
    .Y(_00692_));
 sky130_fd_sc_hd__o21ai_1 _21783_ (.A1(_00689_),
    .A2(_00691_),
    .B1(_00677_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _21784_ (.A(_00678_),
    .B(_00690_),
    .Y(_00694_));
 sky130_fd_sc_hd__o2111ai_1 _21785_ (.A1(_00393_),
    .A2(_00530_),
    .B1(_00536_),
    .C1(_00690_),
    .D1(_00692_),
    .Y(_00695_));
 sky130_fd_sc_hd__o21ai_1 _21786_ (.A1(_00689_),
    .A2(_00691_),
    .B1(_00678_),
    .Y(_00696_));
 sky130_fd_sc_hd__o221ai_4 _21787_ (.A1(_00366_),
    .A2(_00503_),
    .B1(_00691_),
    .B2(_00694_),
    .C1(_00693_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand3_2 _21788_ (.A(_00696_),
    .B(_00675_),
    .C(_00695_),
    .Y(_00699_));
 sky130_fd_sc_hd__a21boi_1 _21789_ (.A1(_00697_),
    .A2(_00699_),
    .B1_N(_00674_),
    .Y(_00700_));
 sky130_fd_sc_hd__a21bo_1 _21790_ (.A1(_00697_),
    .A2(_00699_),
    .B1_N(_00674_),
    .X(_00701_));
 sky130_fd_sc_hd__o211a_1 _21791_ (.A1(_00542_),
    .A2(_00547_),
    .B1(_00697_),
    .C1(_00699_),
    .X(_00702_));
 sky130_fd_sc_hd__o211ai_2 _21792_ (.A1(_00542_),
    .A2(_00547_),
    .B1(_00697_),
    .C1(_00699_),
    .Y(_00703_));
 sky130_fd_sc_hd__o21ai_2 _21793_ (.A1(_00700_),
    .A2(_00702_),
    .B1(_00672_),
    .Y(_00704_));
 sky130_fd_sc_hd__inv_2 _21794_ (.A(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__and3_1 _21795_ (.A(_00673_),
    .B(_00701_),
    .C(_00703_),
    .X(_00706_));
 sky130_fd_sc_hd__nand3_1 _21796_ (.A(_00673_),
    .B(_00701_),
    .C(_00703_),
    .Y(_00707_));
 sky130_fd_sc_hd__and2_1 _21797_ (.A(_00575_),
    .B(_00576_),
    .X(_00708_));
 sky130_fd_sc_hd__and4_1 _21798_ (.A(_02076_),
    .B(net16),
    .C(net56),
    .D(net57),
    .X(_00710_));
 sky130_fd_sc_hd__or4_2 _21799_ (.A(net15),
    .B(_02098_),
    .C(_02229_),
    .D(_02240_),
    .X(_00711_));
 sky130_fd_sc_hd__o22a_1 _21800_ (.A1(net15),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02098_),
    .X(_00712_));
 sky130_fd_sc_hd__nor2_1 _21801_ (.A(_00710_),
    .B(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__o31ai_1 _21802_ (.A1(_02098_),
    .A2(_02207_),
    .A3(_00570_),
    .B1(_00568_),
    .Y(_00714_));
 sky130_fd_sc_hd__and2_1 _21803_ (.A(net17),
    .B(net54),
    .X(_00715_));
 sky130_fd_sc_hd__nand2_1 _21804_ (.A(net19),
    .B(net53),
    .Y(_00716_));
 sky130_fd_sc_hd__nand4_1 _21805_ (.A(net18),
    .B(net19),
    .C(net52),
    .D(net53),
    .Y(_00717_));
 sky130_fd_sc_hd__a22o_1 _21806_ (.A1(net19),
    .A2(net52),
    .B1(net53),
    .B2(net18),
    .X(_00718_));
 sky130_fd_sc_hd__a22oi_2 _21807_ (.A1(net17),
    .A2(net54),
    .B1(_00717_),
    .B2(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__a22o_1 _21808_ (.A1(net17),
    .A2(net54),
    .B1(_00717_),
    .B2(_00718_),
    .X(_00721_));
 sky130_fd_sc_hd__and3_1 _21809_ (.A(_00718_),
    .B(_00715_),
    .C(_00717_),
    .X(_00722_));
 sky130_fd_sc_hd__o2111ai_1 _21810_ (.A1(_00569_),
    .A2(_00716_),
    .B1(net17),
    .C1(net54),
    .D1(_00718_),
    .Y(_00723_));
 sky130_fd_sc_hd__o21bai_4 _21811_ (.A1(_00719_),
    .A2(_00722_),
    .B1_N(_00714_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand3_2 _21812_ (.A(_00714_),
    .B(_00721_),
    .C(_00723_),
    .Y(_00725_));
 sky130_fd_sc_hd__a21boi_1 _21813_ (.A1(_00724_),
    .A2(_00725_),
    .B1_N(_00713_),
    .Y(_00726_));
 sky130_fd_sc_hd__a21bo_1 _21814_ (.A1(_00724_),
    .A2(_00725_),
    .B1_N(_00713_),
    .X(_00727_));
 sky130_fd_sc_hd__o211a_1 _21815_ (.A1(_00710_),
    .A2(_00712_),
    .B1(_00724_),
    .C1(_00725_),
    .X(_00728_));
 sky130_fd_sc_hd__o211ai_2 _21816_ (.A1(_00710_),
    .A2(_00712_),
    .B1(_00724_),
    .C1(_00725_),
    .Y(_00729_));
 sky130_fd_sc_hd__o2bb2a_1 _21817_ (.A1_N(_00575_),
    .A2_N(_00576_),
    .B1(_00726_),
    .B2(_00728_),
    .X(_00730_));
 sky130_fd_sc_hd__o2bb2ai_2 _21818_ (.A1_N(_00575_),
    .A2_N(_00576_),
    .B1(_00726_),
    .B2(_00728_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand4_2 _21819_ (.A(_00575_),
    .B(_00576_),
    .C(_00727_),
    .D(_00729_),
    .Y(_00733_));
 sky130_fd_sc_hd__a21oi_1 _21820_ (.A1(_00732_),
    .A2(_00733_),
    .B1(_00562_),
    .Y(_00734_));
 sky130_fd_sc_hd__a31oi_2 _21821_ (.A1(_00727_),
    .A2(_00729_),
    .A3(_00708_),
    .B1(_00563_),
    .Y(_00735_));
 sky130_fd_sc_hd__a31o_1 _21822_ (.A1(_00727_),
    .A2(_00729_),
    .A3(_00708_),
    .B1(_00563_),
    .X(_00736_));
 sky130_fd_sc_hd__and3_1 _21823_ (.A(_00733_),
    .B(_00562_),
    .C(_00732_),
    .X(_00737_));
 sky130_fd_sc_hd__o311a_1 _21824_ (.A1(net14),
    .A2(_02240_),
    .A3(_00561_),
    .B1(_00732_),
    .C1(_00733_),
    .X(_00738_));
 sky130_fd_sc_hd__a21oi_2 _21825_ (.A1(_00732_),
    .A2(_00733_),
    .B1(_00563_),
    .Y(_00739_));
 sky130_fd_sc_hd__nor2_1 _21826_ (.A(_00738_),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__o2bb2ai_1 _21827_ (.A1_N(_00704_),
    .A2_N(_00707_),
    .B1(_00734_),
    .B2(_00737_),
    .Y(_00741_));
 sky130_fd_sc_hd__o21ai_1 _21828_ (.A1(_00738_),
    .A2(_00739_),
    .B1(_00704_),
    .Y(_00743_));
 sky130_fd_sc_hd__o2bb2ai_1 _21829_ (.A1_N(_00704_),
    .A2_N(_00707_),
    .B1(_00738_),
    .B2(_00739_),
    .Y(_00744_));
 sky130_fd_sc_hd__nand3_1 _21830_ (.A(_00704_),
    .B(_00707_),
    .C(_00740_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand3_2 _21831_ (.A(_00744_),
    .B(_00745_),
    .C(_00671_),
    .Y(_00746_));
 sky130_fd_sc_hd__inv_2 _21832_ (.A(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hd__o221ai_4 _21833_ (.A1(_00510_),
    .A2(_00515_),
    .B1(_00706_),
    .B2(_00743_),
    .C1(_00741_),
    .Y(_00748_));
 sky130_fd_sc_hd__a22o_1 _21834_ (.A1(_00559_),
    .A2(_00588_),
    .B1(_00746_),
    .B2(_00748_),
    .X(_00749_));
 sky130_fd_sc_hd__nand4_1 _21835_ (.A(_00559_),
    .B(_00588_),
    .C(_00746_),
    .D(_00748_),
    .Y(_00750_));
 sky130_fd_sc_hd__a21oi_1 _21836_ (.A1(_00746_),
    .A2(_00748_),
    .B1(_00670_),
    .Y(_00751_));
 sky130_fd_sc_hd__a21o_1 _21837_ (.A1(_00746_),
    .A2(_00748_),
    .B1(_00670_),
    .X(_00752_));
 sky130_fd_sc_hd__nand3_1 _21838_ (.A(_00670_),
    .B(_00746_),
    .C(_00748_),
    .Y(_00754_));
 sky130_fd_sc_hd__nand3_1 _21839_ (.A(_00669_),
    .B(_00749_),
    .C(_00750_),
    .Y(_00755_));
 sky130_fd_sc_hd__o21ai_2 _21840_ (.A1(_00667_),
    .A2(_00668_),
    .B1(_00754_),
    .Y(_00756_));
 sky130_fd_sc_hd__o211ai_2 _21841_ (.A1(_00667_),
    .A2(_00668_),
    .B1(_00752_),
    .C1(_00754_),
    .Y(_00757_));
 sky130_fd_sc_hd__o21ai_2 _21842_ (.A1(_00751_),
    .A2(_00756_),
    .B1(_00755_),
    .Y(_00758_));
 sky130_fd_sc_hd__a221oi_1 _21843_ (.A1(_00601_),
    .A2(_00596_),
    .B1(_00757_),
    .B2(_00755_),
    .C1(_00520_),
    .Y(_00759_));
 sky130_fd_sc_hd__a221o_1 _21844_ (.A1(_00601_),
    .A2(_00596_),
    .B1(_00757_),
    .B2(_00755_),
    .C1(_00520_),
    .X(_00760_));
 sky130_fd_sc_hd__a21oi_2 _21845_ (.A1(_00521_),
    .A2(_00602_),
    .B1(_00758_),
    .Y(_00761_));
 sky130_fd_sc_hd__a31o_1 _21846_ (.A1(_00419_),
    .A2(_00446_),
    .A3(_00594_),
    .B1(_00592_),
    .X(_00762_));
 sky130_fd_sc_hd__o21ai_1 _21847_ (.A1(_00759_),
    .A2(_00761_),
    .B1(_00762_),
    .Y(_00763_));
 sky130_fd_sc_hd__a21oi_1 _21848_ (.A1(_00638_),
    .A2(_00758_),
    .B1(_00762_),
    .Y(_00765_));
 sky130_fd_sc_hd__a31o_1 _21849_ (.A1(_00521_),
    .A2(_00602_),
    .A3(_00758_),
    .B1(_00762_),
    .X(_00766_));
 sky130_fd_sc_hd__o21ai_1 _21850_ (.A1(_00761_),
    .A2(_00766_),
    .B1(_00763_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand2_1 _21851_ (.A(_00767_),
    .B(_00636_),
    .Y(_00768_));
 sky130_fd_sc_hd__o211ai_2 _21852_ (.A1(_00761_),
    .A2(_00766_),
    .B1(_00763_),
    .C1(_00637_),
    .Y(_00769_));
 sky130_fd_sc_hd__a32o_1 _21853_ (.A1(_00560_),
    .A2(_00576_),
    .A3(_00577_),
    .B1(_00581_),
    .B2(_00421_),
    .X(_00770_));
 sky130_fd_sc_hd__a21o_1 _21854_ (.A1(_00768_),
    .A2(_00769_),
    .B1(_00770_),
    .X(_00771_));
 sky130_fd_sc_hd__nand3_2 _21855_ (.A(_00768_),
    .B(_00769_),
    .C(_00770_),
    .Y(_00772_));
 sky130_fd_sc_hd__a31oi_1 _21856_ (.A1(_00612_),
    .A2(_00614_),
    .A3(_00613_),
    .B1(_00619_),
    .Y(_00773_));
 sky130_fd_sc_hd__a31o_1 _21857_ (.A1(_00614_),
    .A2(_00613_),
    .A3(_00612_),
    .B1(_00619_),
    .X(_00774_));
 sky130_fd_sc_hd__o2bb2ai_2 _21858_ (.A1_N(_00771_),
    .A2_N(_00772_),
    .B1(_00773_),
    .B2(_00616_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand4_1 _21859_ (.A(_00617_),
    .B(_00771_),
    .C(_00772_),
    .D(_00774_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _21860_ (.A(_00776_),
    .B(_00777_),
    .Y(_00778_));
 sky130_fd_sc_hd__a31oi_1 _21861_ (.A1(_00484_),
    .A2(_00621_),
    .A3(_00624_),
    .B1(_00634_),
    .Y(_00779_));
 sky130_fd_sc_hd__xor2_1 _21862_ (.A(_00778_),
    .B(_00779_),
    .X(net113));
 sky130_fd_sc_hd__o21ai_1 _21863_ (.A1(_00758_),
    .A2(_00638_),
    .B1(_00762_),
    .Y(_00780_));
 sky130_fd_sc_hd__o311a_1 _21864_ (.A1(_00525_),
    .A2(_00553_),
    .A3(_00555_),
    .B1(_00588_),
    .C1(_00748_),
    .X(_00781_));
 sky130_fd_sc_hd__nand2_1 _21865_ (.A(_00748_),
    .B(_00754_),
    .Y(_00782_));
 sky130_fd_sc_hd__o22a_1 _21866_ (.A1(_00639_),
    .A2(_00664_),
    .B1(_00751_),
    .B2(_00756_),
    .X(_00783_));
 sky130_fd_sc_hd__o22ai_1 _21867_ (.A1(_00639_),
    .A2(_00664_),
    .B1(_00751_),
    .B2(_00756_),
    .Y(_00784_));
 sky130_fd_sc_hd__o31a_1 _21868_ (.A1(_10885_),
    .A2(_00658_),
    .A3(_00660_),
    .B1(_10888_),
    .X(_00786_));
 sky130_fd_sc_hd__o31a_1 _21869_ (.A1(_10798_),
    .A2(_10804_),
    .A3(_11111_),
    .B1(_00652_),
    .X(_00787_));
 sky130_fd_sc_hd__and2_1 _21870_ (.A(net48),
    .B(net25),
    .X(_00788_));
 sky130_fd_sc_hd__nand2_1 _21871_ (.A(net48),
    .B(net25),
    .Y(_00789_));
 sky130_fd_sc_hd__o211ai_4 _21872_ (.A1(_02087_),
    .A2(_00492_),
    .B1(_00642_),
    .C1(_00788_),
    .Y(_00790_));
 sky130_fd_sc_hd__o21ai_2 _21873_ (.A1(_00644_),
    .A2(_00493_),
    .B1(_00789_),
    .Y(_00791_));
 sky130_fd_sc_hd__and3_4 _21874_ (.A(_00791_),
    .B(_00489_),
    .C(_00790_),
    .X(_00792_));
 sky130_fd_sc_hd__o2111ai_4 _21875_ (.A1(_00209_),
    .A2(_00357_),
    .B1(_00367_),
    .C1(_00790_),
    .D1(_00791_),
    .Y(_00793_));
 sky130_fd_sc_hd__a21oi_1 _21876_ (.A1(_00790_),
    .A2(_00791_),
    .B1(_00489_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand3b_4 _21877_ (.A_N(_00794_),
    .B(_00192_),
    .C(_00793_),
    .Y(_00795_));
 sky130_fd_sc_hd__o21ai_2 _21878_ (.A1(_00792_),
    .A2(_00794_),
    .B1(_00193_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_4 _21879_ (.A(_00795_),
    .B(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__a21oi_4 _21880_ (.A1(_10482_),
    .A2(_10749_),
    .B1(_00798_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand3_4 _21881_ (.A(_10894_),
    .B(_00795_),
    .C(_00797_),
    .Y(_00800_));
 sky130_fd_sc_hd__nand2_4 _21882_ (.A(_10892_),
    .B(_00798_),
    .Y(_00801_));
 sky130_fd_sc_hd__inv_2 _21883_ (.A(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__a21bo_1 _21884_ (.A1(_00800_),
    .A2(_00801_),
    .B1_N(_00787_),
    .X(_00803_));
 sky130_fd_sc_hd__nand3b_2 _21885_ (.A_N(_00787_),
    .B(_00800_),
    .C(_00801_),
    .Y(_00804_));
 sky130_fd_sc_hd__a22o_1 _21886_ (.A1(_10886_),
    .A2(_10888_),
    .B1(_00803_),
    .B2(_00804_),
    .X(_00805_));
 sky130_fd_sc_hd__o2111ai_4 _21887_ (.A1(_09384_),
    .A2(_10750_),
    .B1(_10888_),
    .C1(_00803_),
    .D1(_00804_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand2_1 _21888_ (.A(_00805_),
    .B(_00806_),
    .Y(_00808_));
 sky130_fd_sc_hd__a21oi_1 _21889_ (.A1(_00805_),
    .A2(_00806_),
    .B1(_00786_),
    .Y(_00809_));
 sky130_fd_sc_hd__a21o_1 _21890_ (.A1(_00805_),
    .A2(_00806_),
    .B1(_00786_),
    .X(_00810_));
 sky130_fd_sc_hd__and3_1 _21891_ (.A(_00786_),
    .B(_00805_),
    .C(_00806_),
    .X(_00811_));
 sky130_fd_sc_hd__nand3_1 _21892_ (.A(_00786_),
    .B(_00805_),
    .C(_00806_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _21893_ (.A(_00810_),
    .B(_00812_),
    .Y(_00813_));
 sky130_fd_sc_hd__o21a_1 _21894_ (.A1(_10892_),
    .A2(_00655_),
    .B1(_00661_),
    .X(_00814_));
 sky130_fd_sc_hd__nand2_1 _21895_ (.A(_00697_),
    .B(_00703_),
    .Y(_00815_));
 sky130_fd_sc_hd__a31o_1 _21896_ (.A1(_00648_),
    .A2(_00489_),
    .A3(_00646_),
    .B1(_00366_),
    .X(_00816_));
 sky130_fd_sc_hd__o21ai_1 _21897_ (.A1(_00641_),
    .A2(_00644_),
    .B1(_00494_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_1 _21898_ (.A(net49),
    .B(net24),
    .Y(_00819_));
 sky130_fd_sc_hd__a22o_1 _21899_ (.A1(net50),
    .A2(net22),
    .B1(net24),
    .B2(net49),
    .X(_00820_));
 sky130_fd_sc_hd__nand2_1 _21900_ (.A(net50),
    .B(net24),
    .Y(_00821_));
 sky130_fd_sc_hd__nand4_4 _21901_ (.A(net49),
    .B(net50),
    .C(net22),
    .D(net24),
    .Y(_00822_));
 sky130_fd_sc_hd__nand3_1 _21902_ (.A(_00819_),
    .B(net22),
    .C(net50),
    .Y(_00823_));
 sky130_fd_sc_hd__nand3_1 _21903_ (.A(_00680_),
    .B(net24),
    .C(net49),
    .Y(_00824_));
 sky130_fd_sc_hd__and2_1 _21904_ (.A(net51),
    .B(net21),
    .X(_00825_));
 sky130_fd_sc_hd__o211ai_2 _21905_ (.A1(_02152_),
    .A2(_02185_),
    .B1(_00823_),
    .C1(_00824_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand3_4 _21906_ (.A(_00820_),
    .B(_00822_),
    .C(_00825_),
    .Y(_00827_));
 sky130_fd_sc_hd__a21oi_1 _21907_ (.A1(_00826_),
    .A2(_00827_),
    .B1(_00817_),
    .Y(_00828_));
 sky130_fd_sc_hd__a21o_1 _21908_ (.A1(_00826_),
    .A2(_00827_),
    .B1(_00817_),
    .X(_00830_));
 sky130_fd_sc_hd__and3_1 _21909_ (.A(_00817_),
    .B(_00826_),
    .C(_00827_),
    .X(_00831_));
 sky130_fd_sc_hd__o211ai_2 _21910_ (.A1(_00493_),
    .A2(_00645_),
    .B1(_00826_),
    .C1(_00827_),
    .Y(_00832_));
 sky130_fd_sc_hd__o21ai_2 _21911_ (.A1(_00530_),
    .A2(_00681_),
    .B1(_00688_),
    .Y(_00833_));
 sky130_fd_sc_hd__and3_1 _21912_ (.A(_00830_),
    .B(_00832_),
    .C(_00833_),
    .X(_00834_));
 sky130_fd_sc_hd__nand3_2 _21913_ (.A(_00830_),
    .B(_00832_),
    .C(_00833_),
    .Y(_00835_));
 sky130_fd_sc_hd__o21bai_2 _21914_ (.A1(_00828_),
    .A2(_00831_),
    .B1_N(_00833_),
    .Y(_00836_));
 sky130_fd_sc_hd__o21ai_1 _21915_ (.A1(_00366_),
    .A2(_00649_),
    .B1(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__o211a_1 _21916_ (.A1(_00366_),
    .A2(_00649_),
    .B1(_00835_),
    .C1(_00836_),
    .X(_00838_));
 sky130_fd_sc_hd__a21oi_2 _21917_ (.A1(_00835_),
    .A2(_00836_),
    .B1(_00816_),
    .Y(_00839_));
 sky130_fd_sc_hd__a21o_1 _21918_ (.A1(_00835_),
    .A2(_00836_),
    .B1(_00816_),
    .X(_00841_));
 sky130_fd_sc_hd__o21ai_2 _21919_ (.A1(_00677_),
    .A2(_00689_),
    .B1(_00692_),
    .Y(_00842_));
 sky130_fd_sc_hd__inv_2 _21920_ (.A(_00842_),
    .Y(_00843_));
 sky130_fd_sc_hd__o21ai_2 _21921_ (.A1(_00838_),
    .A2(_00839_),
    .B1(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__a31o_1 _21922_ (.A1(_00816_),
    .A2(_00835_),
    .A3(_00836_),
    .B1(_00843_),
    .X(_00845_));
 sky130_fd_sc_hd__o211ai_1 _21923_ (.A1(_00834_),
    .A2(_00837_),
    .B1(_00842_),
    .C1(_00841_),
    .Y(_00846_));
 sky130_fd_sc_hd__a21oi_1 _21924_ (.A1(_00844_),
    .A2(_00846_),
    .B1(_00815_),
    .Y(_00847_));
 sky130_fd_sc_hd__a21o_1 _21925_ (.A1(_00844_),
    .A2(_00846_),
    .B1(_00815_),
    .X(_00848_));
 sky130_fd_sc_hd__o211a_1 _21926_ (.A1(_00839_),
    .A2(_00845_),
    .B1(_00844_),
    .C1(_00815_),
    .X(_00849_));
 sky130_fd_sc_hd__o211ai_2 _21927_ (.A1(_00839_),
    .A2(_00845_),
    .B1(_00844_),
    .C1(_00815_),
    .Y(_00850_));
 sky130_fd_sc_hd__a21boi_1 _21928_ (.A1(_00724_),
    .A2(_00713_),
    .B1_N(_00725_),
    .Y(_00852_));
 sky130_fd_sc_hd__a21bo_1 _21929_ (.A1(_00713_),
    .A2(_00724_),
    .B1_N(_00725_),
    .X(_00853_));
 sky130_fd_sc_hd__and4_2 _21930_ (.A(_02098_),
    .B(net17),
    .C(net56),
    .D(net57),
    .X(_00854_));
 sky130_fd_sc_hd__nand4_1 _21931_ (.A(_02098_),
    .B(net17),
    .C(net56),
    .D(net57),
    .Y(_00855_));
 sky130_fd_sc_hd__o2bb2a_1 _21932_ (.A1_N(net17),
    .A2_N(net56),
    .B1(net16),
    .B2(_02240_),
    .X(_00856_));
 sky130_fd_sc_hd__nor2_1 _21933_ (.A(_00854_),
    .B(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__o2bb2ai_1 _21934_ (.A1_N(_00715_),
    .A2_N(_00718_),
    .B1(_00716_),
    .B2(_00569_),
    .Y(_00858_));
 sky130_fd_sc_hd__nand4_2 _21935_ (.A(net19),
    .B(net20),
    .C(net52),
    .D(net53),
    .Y(_00859_));
 sky130_fd_sc_hd__a22oi_1 _21936_ (.A1(net20),
    .A2(net52),
    .B1(net53),
    .B2(net19),
    .Y(_00860_));
 sky130_fd_sc_hd__a22o_1 _21937_ (.A1(net20),
    .A2(net52),
    .B1(net53),
    .B2(net19),
    .X(_00861_));
 sky130_fd_sc_hd__a22oi_1 _21938_ (.A1(net18),
    .A2(net54),
    .B1(_00859_),
    .B2(_00861_),
    .Y(_00863_));
 sky130_fd_sc_hd__a22o_1 _21939_ (.A1(net18),
    .A2(net54),
    .B1(_00859_),
    .B2(_00861_),
    .X(_00864_));
 sky130_fd_sc_hd__and4_1 _21940_ (.A(_00861_),
    .B(net54),
    .C(net18),
    .D(_00859_),
    .X(_00865_));
 sky130_fd_sc_hd__nand4_1 _21941_ (.A(_00861_),
    .B(net54),
    .C(net18),
    .D(_00859_),
    .Y(_00866_));
 sky130_fd_sc_hd__o21bai_2 _21942_ (.A1(_00863_),
    .A2(_00865_),
    .B1_N(_00858_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand3_2 _21943_ (.A(_00858_),
    .B(_00864_),
    .C(_00866_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand3_2 _21944_ (.A(_00867_),
    .B(_00868_),
    .C(_00857_),
    .Y(_00869_));
 sky130_fd_sc_hd__a2bb2o_1 _21945_ (.A1_N(_00854_),
    .A2_N(_00856_),
    .B1(_00867_),
    .B2(_00868_),
    .X(_00870_));
 sky130_fd_sc_hd__a21bo_1 _21946_ (.A1(_00867_),
    .A2(_00868_),
    .B1_N(_00857_),
    .X(_00871_));
 sky130_fd_sc_hd__o211ai_2 _21947_ (.A1(_00854_),
    .A2(_00856_),
    .B1(_00867_),
    .C1(_00868_),
    .Y(_00872_));
 sky130_fd_sc_hd__nand3_2 _21948_ (.A(_00853_),
    .B(_00869_),
    .C(_00870_),
    .Y(_00874_));
 sky130_fd_sc_hd__nand3_1 _21949_ (.A(_00871_),
    .B(_00872_),
    .C(_00852_),
    .Y(_00875_));
 sky130_fd_sc_hd__a21oi_1 _21950_ (.A1(_00874_),
    .A2(_00875_),
    .B1(_00710_),
    .Y(_00876_));
 sky130_fd_sc_hd__a31oi_2 _21951_ (.A1(_00871_),
    .A2(_00872_),
    .A3(_00852_),
    .B1(_00711_),
    .Y(_00877_));
 sky130_fd_sc_hd__a31o_1 _21952_ (.A1(_00871_),
    .A2(_00872_),
    .A3(_00852_),
    .B1(_00711_),
    .X(_00878_));
 sky130_fd_sc_hd__nand3_1 _21953_ (.A(_00711_),
    .B(_00874_),
    .C(_00875_),
    .Y(_00879_));
 sky130_fd_sc_hd__a21o_1 _21954_ (.A1(_00874_),
    .A2(_00875_),
    .B1(_00711_),
    .X(_00880_));
 sky130_fd_sc_hd__a21oi_2 _21955_ (.A1(_00874_),
    .A2(_00877_),
    .B1(_00876_),
    .Y(_00881_));
 sky130_fd_sc_hd__o21bai_1 _21956_ (.A1(_00847_),
    .A2(_00849_),
    .B1_N(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand3_1 _21957_ (.A(_00848_),
    .B(_00850_),
    .C(_00881_),
    .Y(_00883_));
 sky130_fd_sc_hd__o21ai_1 _21958_ (.A1(_00847_),
    .A2(_00849_),
    .B1(_00881_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand4_1 _21959_ (.A(_00848_),
    .B(_00850_),
    .C(_00879_),
    .D(_00880_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand3_2 _21960_ (.A(_00885_),
    .B(_00886_),
    .C(_00814_),
    .Y(_00887_));
 sky130_fd_sc_hd__nand3b_2 _21961_ (.A_N(_00814_),
    .B(_00882_),
    .C(_00883_),
    .Y(_00888_));
 sky130_fd_sc_hd__o32a_1 _21962_ (.A1(_00672_),
    .A2(_00700_),
    .A3(_00702_),
    .B1(_00734_),
    .B2(_00737_),
    .X(_00889_));
 sky130_fd_sc_hd__o31a_1 _21963_ (.A1(_00706_),
    .A2(_00738_),
    .A3(_00739_),
    .B1(_00704_),
    .X(_00890_));
 sky130_fd_sc_hd__o2bb2ai_2 _21964_ (.A1_N(_00887_),
    .A2_N(_00888_),
    .B1(_00889_),
    .B2(_00705_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand3_2 _21965_ (.A(_00890_),
    .B(_00888_),
    .C(_00887_),
    .Y(_00892_));
 sky130_fd_sc_hd__a21oi_2 _21966_ (.A1(_00891_),
    .A2(_00892_),
    .B1(_00813_),
    .Y(_00893_));
 sky130_fd_sc_hd__a32oi_2 _21967_ (.A1(_00890_),
    .A2(_00888_),
    .A3(_00887_),
    .B1(_00810_),
    .B2(_00812_),
    .Y(_00894_));
 sky130_fd_sc_hd__o211a_1 _21968_ (.A1(_00809_),
    .A2(_00811_),
    .B1(_00891_),
    .C1(_00892_),
    .X(_00896_));
 sky130_fd_sc_hd__o211ai_2 _21969_ (.A1(_00809_),
    .A2(_00811_),
    .B1(_00891_),
    .C1(_00892_),
    .Y(_00897_));
 sky130_fd_sc_hd__nand2_1 _21970_ (.A(_00784_),
    .B(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__a221oi_2 _21971_ (.A1(_00894_),
    .A2(_00891_),
    .B1(_00757_),
    .B2(_00666_),
    .C1(_00893_),
    .Y(_00899_));
 sky130_fd_sc_hd__o21a_1 _21972_ (.A1(_00893_),
    .A2(_00896_),
    .B1(_00783_),
    .X(_00900_));
 sky130_fd_sc_hd__o21ai_1 _21973_ (.A1(_00893_),
    .A2(_00896_),
    .B1(_00783_),
    .Y(_00901_));
 sky130_fd_sc_hd__o211a_1 _21974_ (.A1(_00893_),
    .A2(_00898_),
    .B1(_00782_),
    .C1(_00901_),
    .X(_00902_));
 sky130_fd_sc_hd__o211ai_2 _21975_ (.A1(_00893_),
    .A2(_00898_),
    .B1(_00901_),
    .C1(_00782_),
    .Y(_00903_));
 sky130_fd_sc_hd__o22a_1 _21976_ (.A1(_00747_),
    .A2(_00781_),
    .B1(_00899_),
    .B2(_00900_),
    .X(_00904_));
 sky130_fd_sc_hd__o22ai_2 _21977_ (.A1(_00747_),
    .A2(_00781_),
    .B1(_00899_),
    .B2(_00900_),
    .Y(_00905_));
 sky130_fd_sc_hd__o211a_1 _21978_ (.A1(_00761_),
    .A2(_00765_),
    .B1(_00903_),
    .C1(_00905_),
    .X(_00907_));
 sky130_fd_sc_hd__o211ai_2 _21979_ (.A1(_00761_),
    .A2(_00765_),
    .B1(_00903_),
    .C1(_00905_),
    .Y(_00908_));
 sky130_fd_sc_hd__a22oi_1 _21980_ (.A1(_00760_),
    .A2(_00780_),
    .B1(_00903_),
    .B2(_00905_),
    .Y(_00909_));
 sky130_fd_sc_hd__o2bb2ai_1 _21981_ (.A1_N(_00760_),
    .A2_N(_00780_),
    .B1(_00902_),
    .B2(_00904_),
    .Y(_00910_));
 sky130_fd_sc_hd__o211ai_2 _21982_ (.A1(_00730_),
    .A2(_00735_),
    .B1(_00908_),
    .C1(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__o31a_1 _21983_ (.A1(_00730_),
    .A2(_00735_),
    .A3(_00907_),
    .B1(_00910_),
    .X(_00912_));
 sky130_fd_sc_hd__o211ai_2 _21984_ (.A1(_00907_),
    .A2(_00909_),
    .B1(_00732_),
    .C1(_00736_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand2_1 _21985_ (.A(_00911_),
    .B(_00913_),
    .Y(_00914_));
 sky130_fd_sc_hd__o21ai_1 _21986_ (.A1(_00636_),
    .A2(_00767_),
    .B1(_00772_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand3_1 _21987_ (.A(_00914_),
    .B(_00772_),
    .C(_00769_),
    .Y(_00916_));
 sky130_fd_sc_hd__and3_1 _21988_ (.A(_00915_),
    .B(_00913_),
    .C(_00911_),
    .X(_00918_));
 sky130_fd_sc_hd__nand3_2 _21989_ (.A(_00915_),
    .B(_00913_),
    .C(_00911_),
    .Y(_00919_));
 sky130_fd_sc_hd__and2_1 _21990_ (.A(_00916_),
    .B(_00919_),
    .X(_00920_));
 sky130_fd_sc_hd__o21ai_1 _21991_ (.A1(_00485_),
    .A2(_00625_),
    .B1(_00777_),
    .Y(_00921_));
 sky130_fd_sc_hd__o21a_1 _21992_ (.A1(_00921_),
    .A2(_00634_),
    .B1(_00776_),
    .X(_00922_));
 sky130_fd_sc_hd__o2111ai_1 _21993_ (.A1(_00921_),
    .A2(_00634_),
    .B1(_00916_),
    .C1(_00919_),
    .D1(_00776_),
    .Y(_00923_));
 sky130_fd_sc_hd__xor2_1 _21994_ (.A(_00920_),
    .B(_00922_),
    .X(net114));
 sky130_fd_sc_hd__a31o_1 _21995_ (.A1(_10886_),
    .A2(_00803_),
    .A3(_00804_),
    .B1(_10887_),
    .X(_00924_));
 sky130_fd_sc_hd__o21ai_4 _21996_ (.A1(_10804_),
    .A2(_11117_),
    .B1(_00795_),
    .Y(_00925_));
 sky130_fd_sc_hd__a21oi_2 _21997_ (.A1(_00800_),
    .A2(_00801_),
    .B1(_00925_),
    .Y(_00926_));
 sky130_fd_sc_hd__a21o_1 _21998_ (.A1(_00800_),
    .A2(_00801_),
    .B1(_00925_),
    .X(_00928_));
 sky130_fd_sc_hd__a22oi_4 _21999_ (.A1(_00191_),
    .A2(_00795_),
    .B1(_10892_),
    .B2(_00798_),
    .Y(_00929_));
 sky130_fd_sc_hd__and3_2 _22000_ (.A(_00800_),
    .B(_00801_),
    .C(_00925_),
    .X(_00930_));
 sky130_fd_sc_hd__o21ai_4 _22001_ (.A1(_10892_),
    .A2(_00798_),
    .B1(_00929_),
    .Y(_00931_));
 sky130_fd_sc_hd__a21oi_2 _22002_ (.A1(_00800_),
    .A2(_00929_),
    .B1(_00926_),
    .Y(_00932_));
 sky130_fd_sc_hd__a21o_2 _22003_ (.A1(_00800_),
    .A2(_00929_),
    .B1(_00926_),
    .X(_00933_));
 sky130_fd_sc_hd__a22o_1 _22004_ (.A1(_10886_),
    .A2(_10888_),
    .B1(_00928_),
    .B2(_00931_),
    .X(_00934_));
 sky130_fd_sc_hd__a211o_1 _22005_ (.A1(_00800_),
    .A2(_00929_),
    .B1(_00926_),
    .C1(_10890_),
    .X(_00935_));
 sky130_fd_sc_hd__a21oi_1 _22006_ (.A1(_00934_),
    .A2(_00935_),
    .B1(_00924_),
    .Y(_00936_));
 sky130_fd_sc_hd__and3_1 _22007_ (.A(_00924_),
    .B(_00934_),
    .C(_00935_),
    .X(_00937_));
 sky130_fd_sc_hd__nand3_4 _22008_ (.A(_00924_),
    .B(_00934_),
    .C(_00935_),
    .Y(_00939_));
 sky130_fd_sc_hd__nor2_1 _22009_ (.A(_00936_),
    .B(_00937_),
    .Y(_00940_));
 sky130_fd_sc_hd__o22a_1 _22010_ (.A1(_00834_),
    .A2(_00837_),
    .B1(_00843_),
    .B2(_00839_),
    .X(_00941_));
 sky130_fd_sc_hd__o22ai_2 _22011_ (.A1(_00834_),
    .A2(_00837_),
    .B1(_00843_),
    .B2(_00839_),
    .Y(_00942_));
 sky130_fd_sc_hd__a21oi_2 _22012_ (.A1(_00830_),
    .A2(_00833_),
    .B1(_00831_),
    .Y(_00943_));
 sky130_fd_sc_hd__a21o_1 _22013_ (.A1(_00830_),
    .A2(_00833_),
    .B1(_00831_),
    .X(_00944_));
 sky130_fd_sc_hd__o21a_4 _22014_ (.A1(_02054_),
    .A2(_00036_),
    .B1(_00793_),
    .X(_00945_));
 sky130_fd_sc_hd__a31o_1 _22015_ (.A1(_00791_),
    .A2(_00489_),
    .A3(_00790_),
    .B1(_00366_),
    .X(_00946_));
 sky130_fd_sc_hd__o31a_1 _22016_ (.A1(_02120_),
    .A2(_02218_),
    .A3(_00680_),
    .B1(_00827_),
    .X(_00947_));
 sky130_fd_sc_hd__o21ai_1 _22017_ (.A1(_00680_),
    .A2(_00819_),
    .B1(_00827_),
    .Y(_00948_));
 sky130_fd_sc_hd__a21oi_2 _22018_ (.A1(_00642_),
    .A2(_00788_),
    .B1(_00493_),
    .Y(_00950_));
 sky130_fd_sc_hd__o21ai_4 _22019_ (.A1(_00644_),
    .A2(_00789_),
    .B1(_00494_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand2_1 _22020_ (.A(net49),
    .B(net25),
    .Y(_00952_));
 sky130_fd_sc_hd__nand4_4 _22021_ (.A(net49),
    .B(net50),
    .C(net24),
    .D(net25),
    .Y(_00953_));
 sky130_fd_sc_hd__a22o_1 _22022_ (.A1(net50),
    .A2(net24),
    .B1(net25),
    .B2(net49),
    .X(_00954_));
 sky130_fd_sc_hd__nand3_1 _22023_ (.A(_00952_),
    .B(net24),
    .C(net50),
    .Y(_00955_));
 sky130_fd_sc_hd__nand3_1 _22024_ (.A(_00821_),
    .B(net25),
    .C(net49),
    .Y(_00956_));
 sky130_fd_sc_hd__nand4_4 _22025_ (.A(_00954_),
    .B(net22),
    .C(net51),
    .D(_00953_),
    .Y(_00957_));
 sky130_fd_sc_hd__o211ai_4 _22026_ (.A1(_02152_),
    .A2(_02196_),
    .B1(_00955_),
    .C1(_00956_),
    .Y(_00958_));
 sky130_fd_sc_hd__a21oi_4 _22027_ (.A1(_00957_),
    .A2(_00958_),
    .B1(_00951_),
    .Y(_00959_));
 sky130_fd_sc_hd__a21o_1 _22028_ (.A1(_00957_),
    .A2(_00958_),
    .B1(_00951_),
    .X(_00961_));
 sky130_fd_sc_hd__and3_1 _22029_ (.A(_00951_),
    .B(_00957_),
    .C(_00958_),
    .X(_00962_));
 sky130_fd_sc_hd__nand3_1 _22030_ (.A(_00951_),
    .B(_00957_),
    .C(_00958_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand4_4 _22031_ (.A(_00822_),
    .B(_00827_),
    .C(_00961_),
    .D(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__o21ai_2 _22032_ (.A1(_00959_),
    .A2(_00962_),
    .B1(_00948_),
    .Y(_00965_));
 sky130_fd_sc_hd__a31o_1 _22033_ (.A1(_00951_),
    .A2(_00957_),
    .A3(_00958_),
    .B1(_00947_),
    .X(_00966_));
 sky130_fd_sc_hd__o21ai_2 _22034_ (.A1(_00959_),
    .A2(_00962_),
    .B1(_00947_),
    .Y(_00967_));
 sky130_fd_sc_hd__o221a_2 _22035_ (.A1(_00366_),
    .A2(_00792_),
    .B1(_00959_),
    .B2(_00966_),
    .C1(_00967_),
    .X(_00968_));
 sky130_fd_sc_hd__o221ai_4 _22036_ (.A1(_00366_),
    .A2(_00792_),
    .B1(_00959_),
    .B2(_00966_),
    .C1(_00967_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand3_1 _22037_ (.A(_00965_),
    .B(_00945_),
    .C(_00964_),
    .Y(_00970_));
 sky130_fd_sc_hd__a31oi_2 _22038_ (.A1(_00965_),
    .A2(_00945_),
    .A3(_00964_),
    .B1(_00943_),
    .Y(_00972_));
 sky130_fd_sc_hd__a31o_1 _22039_ (.A1(_00965_),
    .A2(_00945_),
    .A3(_00964_),
    .B1(_00943_),
    .X(_00973_));
 sky130_fd_sc_hd__o211a_1 _22040_ (.A1(_00831_),
    .A2(_00834_),
    .B1(_00969_),
    .C1(_00970_),
    .X(_00974_));
 sky130_fd_sc_hd__a21oi_1 _22041_ (.A1(_00969_),
    .A2(_00970_),
    .B1(_00944_),
    .Y(_00975_));
 sky130_fd_sc_hd__a21o_1 _22042_ (.A1(_00969_),
    .A2(_00970_),
    .B1(_00944_),
    .X(_00976_));
 sky130_fd_sc_hd__o21ai_2 _22043_ (.A1(_00974_),
    .A2(_00975_),
    .B1(_00941_),
    .Y(_00977_));
 sky130_fd_sc_hd__o211ai_4 _22044_ (.A1(_00968_),
    .A2(_00973_),
    .B1(_00976_),
    .C1(_00942_),
    .Y(_00978_));
 sky130_fd_sc_hd__and4b_2 _22045_ (.A_N(net17),
    .B(net18),
    .C(net56),
    .D(net57),
    .X(_00979_));
 sky130_fd_sc_hd__o22a_1 _22046_ (.A1(net17),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02131_),
    .X(_00980_));
 sky130_fd_sc_hd__nor2_1 _22047_ (.A(_00979_),
    .B(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__o31ai_1 _22048_ (.A1(_02131_),
    .A2(_02207_),
    .A3(_00860_),
    .B1(_00859_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_1 _22049_ (.A(net21),
    .B(net53),
    .Y(_00984_));
 sky130_fd_sc_hd__nand4_2 _22050_ (.A(net20),
    .B(net52),
    .C(net21),
    .D(net53),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _22051_ (.A(net52),
    .B(net21),
    .Y(_00986_));
 sky130_fd_sc_hd__a22oi_1 _22052_ (.A1(net52),
    .A2(net21),
    .B1(net53),
    .B2(net20),
    .Y(_00987_));
 sky130_fd_sc_hd__a22o_1 _22053_ (.A1(net52),
    .A2(net21),
    .B1(net53),
    .B2(net20),
    .X(_00988_));
 sky130_fd_sc_hd__o2bb2ai_1 _22054_ (.A1_N(_00985_),
    .A2_N(_00988_),
    .B1(_02142_),
    .B2(_02207_),
    .Y(_00989_));
 sky130_fd_sc_hd__and4_1 _22055_ (.A(_00988_),
    .B(net54),
    .C(net19),
    .D(_00985_),
    .X(_00990_));
 sky130_fd_sc_hd__nand4_1 _22056_ (.A(_00988_),
    .B(net54),
    .C(net19),
    .D(_00985_),
    .Y(_00991_));
 sky130_fd_sc_hd__a21o_1 _22057_ (.A1(_00989_),
    .A2(_00991_),
    .B1(_00983_),
    .X(_00992_));
 sky130_fd_sc_hd__nand2_1 _22058_ (.A(_00983_),
    .B(_00989_),
    .Y(_00994_));
 sky130_fd_sc_hd__o21ai_1 _22059_ (.A1(_00990_),
    .A2(_00994_),
    .B1(_00992_),
    .Y(_00995_));
 sky130_fd_sc_hd__nand2_1 _22060_ (.A(_00995_),
    .B(_00981_),
    .Y(_00996_));
 sky130_fd_sc_hd__o221ai_2 _22061_ (.A1(_00979_),
    .A2(_00980_),
    .B1(_00990_),
    .B2(_00994_),
    .C1(_00992_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand4_2 _22062_ (.A(_00868_),
    .B(_00869_),
    .C(_00996_),
    .D(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hd__a22o_1 _22063_ (.A1(_00868_),
    .A2(_00869_),
    .B1(_00996_),
    .B2(_00997_),
    .X(_00999_));
 sky130_fd_sc_hd__a21oi_1 _22064_ (.A1(_00998_),
    .A2(_00999_),
    .B1(_00854_),
    .Y(_01000_));
 sky130_fd_sc_hd__a21o_1 _22065_ (.A1(_00998_),
    .A2(_00999_),
    .B1(_00854_),
    .X(_01001_));
 sky130_fd_sc_hd__and3_1 _22066_ (.A(_00998_),
    .B(_00999_),
    .C(_00854_),
    .X(_01002_));
 sky130_fd_sc_hd__nand3_1 _22067_ (.A(_00998_),
    .B(_00999_),
    .C(_00854_),
    .Y(_01003_));
 sky130_fd_sc_hd__o2bb2ai_2 _22068_ (.A1_N(_00977_),
    .A2_N(_00978_),
    .B1(_01000_),
    .B2(_01002_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand4_4 _22069_ (.A(_00977_),
    .B(_00978_),
    .C(_01001_),
    .D(_01003_),
    .Y(_01006_));
 sky130_fd_sc_hd__o221a_1 _22070_ (.A1(_10804_),
    .A2(_11117_),
    .B1(_00798_),
    .B2(_10892_),
    .C1(_00652_),
    .X(_01007_));
 sky130_fd_sc_hd__o21ai_1 _22071_ (.A1(_00798_),
    .A2(_10892_),
    .B1(_00787_),
    .Y(_01008_));
 sky130_fd_sc_hd__o2bb2ai_2 _22072_ (.A1_N(_01005_),
    .A2_N(_01006_),
    .B1(_01007_),
    .B2(_00802_),
    .Y(_01009_));
 sky130_fd_sc_hd__nand4_4 _22073_ (.A(_00801_),
    .B(_01005_),
    .C(_01006_),
    .D(_01008_),
    .Y(_01010_));
 sky130_fd_sc_hd__and3_1 _22074_ (.A(_00850_),
    .B(_00879_),
    .C(_00880_),
    .X(_01011_));
 sky130_fd_sc_hd__a21o_1 _22075_ (.A1(_00848_),
    .A2(_00881_),
    .B1(_00849_),
    .X(_01012_));
 sky130_fd_sc_hd__o2bb2ai_2 _22076_ (.A1_N(_01009_),
    .A2_N(_01010_),
    .B1(_01011_),
    .B2(_00847_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _22077_ (.A(_01009_),
    .B(_01012_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand3_2 _22078_ (.A(_01009_),
    .B(_01010_),
    .C(_01012_),
    .Y(_01016_));
 sky130_fd_sc_hd__inv_2 _22079_ (.A(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__a2bb2o_1 _22080_ (.A1_N(_00936_),
    .A2_N(_00937_),
    .B1(_01013_),
    .B2(_01016_),
    .X(_01018_));
 sky130_fd_sc_hd__nand2_1 _22081_ (.A(_00940_),
    .B(_01013_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand3_4 _22082_ (.A(_00940_),
    .B(_01013_),
    .C(_01016_),
    .Y(_01020_));
 sky130_fd_sc_hd__o21ai_2 _22083_ (.A1(_00786_),
    .A2(_00808_),
    .B1(_00897_),
    .Y(_01021_));
 sky130_fd_sc_hd__a21oi_1 _22084_ (.A1(_01018_),
    .A2(_01020_),
    .B1(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__a21o_1 _22085_ (.A1(_01018_),
    .A2(_01020_),
    .B1(_01021_),
    .X(_01023_));
 sky130_fd_sc_hd__o211a_1 _22086_ (.A1(_01017_),
    .A2(_01019_),
    .B1(_01021_),
    .C1(_01018_),
    .X(_01024_));
 sky130_fd_sc_hd__o211ai_1 _22087_ (.A1(_01017_),
    .A2(_01019_),
    .B1(_01021_),
    .C1(_01018_),
    .Y(_01025_));
 sky130_fd_sc_hd__nand2_1 _22088_ (.A(_00888_),
    .B(_00892_),
    .Y(_01027_));
 sky130_fd_sc_hd__o21bai_1 _22089_ (.A1(_01022_),
    .A2(_01024_),
    .B1_N(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand3_1 _22090_ (.A(_01023_),
    .B(_01025_),
    .C(_01027_),
    .Y(_01029_));
 sky130_fd_sc_hd__a2bb2o_1 _22091_ (.A1_N(_00893_),
    .A2_N(_00898_),
    .B1(_00782_),
    .B2(_00901_),
    .X(_01030_));
 sky130_fd_sc_hd__a21oi_1 _22092_ (.A1(_01028_),
    .A2(_01029_),
    .B1(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__a21o_1 _22093_ (.A1(_01028_),
    .A2(_01029_),
    .B1(_01030_),
    .X(_01032_));
 sky130_fd_sc_hd__and3_1 _22094_ (.A(_01028_),
    .B(_01030_),
    .C(_01029_),
    .X(_01033_));
 sky130_fd_sc_hd__nand3_1 _22095_ (.A(_01028_),
    .B(_01029_),
    .C(_01030_),
    .Y(_01034_));
 sky130_fd_sc_hd__a31o_1 _22096_ (.A1(_00853_),
    .A2(_00869_),
    .A3(_00870_),
    .B1(_00877_),
    .X(_01035_));
 sky130_fd_sc_hd__nand3_1 _22097_ (.A(_01032_),
    .B(_01034_),
    .C(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__o211a_1 _22098_ (.A1(_01031_),
    .A2(_01033_),
    .B1(_00874_),
    .C1(_00878_),
    .X(_01038_));
 sky130_fd_sc_hd__o21bai_1 _22099_ (.A1(_01031_),
    .A2(_01033_),
    .B1_N(_01035_),
    .Y(_01039_));
 sky130_fd_sc_hd__a21o_1 _22100_ (.A1(_01036_),
    .A2(_01039_),
    .B1(_00912_),
    .X(_01040_));
 sky130_fd_sc_hd__a32o_1 _22101_ (.A1(_01032_),
    .A2(_01034_),
    .A3(_01035_),
    .B1(_00911_),
    .B2(_00908_),
    .X(_01041_));
 sky130_fd_sc_hd__o21ai_1 _22102_ (.A1(_01038_),
    .A2(_01041_),
    .B1(_01040_),
    .Y(_01042_));
 sky130_fd_sc_hd__and3_1 _22103_ (.A(_00919_),
    .B(_00923_),
    .C(_01042_),
    .X(_01043_));
 sky130_fd_sc_hd__a21oi_1 _22104_ (.A1(_00919_),
    .A2(_00923_),
    .B1(_01042_),
    .Y(_01044_));
 sky130_fd_sc_hd__nor2_1 _22105_ (.A(_01043_),
    .B(_01044_),
    .Y(net115));
 sky130_fd_sc_hd__and3_2 _22106_ (.A(_00928_),
    .B(_00931_),
    .C(_10887_),
    .X(_01045_));
 sky130_fd_sc_hd__nand4_4 _22107_ (.A(_00928_),
    .B(_00931_),
    .C(_09385_),
    .D(_10750_),
    .Y(_01046_));
 sky130_fd_sc_hd__o221a_2 _22108_ (.A1(_10746_),
    .A2(_10748_),
    .B1(_00926_),
    .B2(_00930_),
    .C1(_09383_),
    .X(_01048_));
 sky130_fd_sc_hd__o31a_2 _22109_ (.A1(_09384_),
    .A2(_10750_),
    .A3(_00932_),
    .B1(_01046_),
    .X(_01049_));
 sky130_fd_sc_hd__o21ai_2 _22110_ (.A1(_10886_),
    .A2(_00932_),
    .B1(_01046_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand2_1 _22111_ (.A(_00978_),
    .B(_01006_),
    .Y(_01051_));
 sky130_fd_sc_hd__a21oi_2 _22112_ (.A1(_00801_),
    .A2(_00925_),
    .B1(_00799_),
    .Y(_01052_));
 sky130_fd_sc_hd__a21o_2 _22113_ (.A1(_00801_),
    .A2(_00925_),
    .B1(_00799_),
    .X(_01053_));
 sky130_fd_sc_hd__o21ai_2 _22114_ (.A1(_00821_),
    .A2(_00952_),
    .B1(_00957_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _22115_ (.A(net51),
    .B(net24),
    .Y(_01055_));
 sky130_fd_sc_hd__o21ai_4 _22116_ (.A1(net49),
    .A2(net50),
    .B1(net25),
    .Y(_01056_));
 sky130_fd_sc_hd__o21a_2 _22117_ (.A1(net49),
    .A2(net50),
    .B1(net25),
    .X(_01057_));
 sky130_fd_sc_hd__and3_2 _22118_ (.A(net49),
    .B(net50),
    .C(net25),
    .X(_01059_));
 sky130_fd_sc_hd__nand3_4 _22119_ (.A(net49),
    .B(net50),
    .C(net25),
    .Y(_01060_));
 sky130_fd_sc_hd__o211ai_1 _22120_ (.A1(_02152_),
    .A2(_02218_),
    .B1(_01057_),
    .C1(_01060_),
    .Y(_01061_));
 sky130_fd_sc_hd__a21o_1 _22121_ (.A1(_01057_),
    .A2(_01060_),
    .B1(_01055_),
    .X(_01062_));
 sky130_fd_sc_hd__o22ai_1 _22122_ (.A1(_02152_),
    .A2(_02218_),
    .B1(_01056_),
    .B2(_01059_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand4_1 _22123_ (.A(_01057_),
    .B(_01060_),
    .C(net51),
    .D(net24),
    .Y(_01064_));
 sky130_fd_sc_hd__nand3_2 _22124_ (.A(_01062_),
    .B(_00950_),
    .C(_01061_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand3_2 _22125_ (.A(_00951_),
    .B(_01063_),
    .C(_01064_),
    .Y(_01066_));
 sky130_fd_sc_hd__inv_2 _22126_ (.A(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__and3_1 _22127_ (.A(_01054_),
    .B(_01065_),
    .C(_01066_),
    .X(_01068_));
 sky130_fd_sc_hd__nand3_1 _22128_ (.A(_01054_),
    .B(_01065_),
    .C(_01066_),
    .Y(_01070_));
 sky130_fd_sc_hd__a21o_1 _22129_ (.A1(_01065_),
    .A2(_01066_),
    .B1(_01054_),
    .X(_01071_));
 sky130_fd_sc_hd__a22oi_1 _22130_ (.A1(_00953_),
    .A2(_00957_),
    .B1(_01065_),
    .B2(_01066_),
    .Y(_01072_));
 sky130_fd_sc_hd__a22o_1 _22131_ (.A1(_00953_),
    .A2(_00957_),
    .B1(_01065_),
    .B2(_01066_),
    .X(_01073_));
 sky130_fd_sc_hd__nand4_1 _22132_ (.A(_00953_),
    .B(_00957_),
    .C(_01065_),
    .D(_01066_),
    .Y(_01074_));
 sky130_fd_sc_hd__o211ai_2 _22133_ (.A1(_00366_),
    .A2(_00792_),
    .B1(_01070_),
    .C1(_01071_),
    .Y(_01075_));
 sky130_fd_sc_hd__nor3b_1 _22134_ (.A(_00946_),
    .B(_01072_),
    .C_N(_01074_),
    .Y(_01076_));
 sky130_fd_sc_hd__nand3_1 _22135_ (.A(_01073_),
    .B(_01074_),
    .C(_00945_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand4_1 _22136_ (.A(_00367_),
    .B(_00793_),
    .C(_01070_),
    .D(_01071_),
    .Y(_01078_));
 sky130_fd_sc_hd__o211ai_1 _22137_ (.A1(_00366_),
    .A2(_00792_),
    .B1(_01073_),
    .C1(_01074_),
    .Y(_01079_));
 sky130_fd_sc_hd__a32o_1 _22138_ (.A1(_00951_),
    .A2(_00957_),
    .A3(_00958_),
    .B1(_00961_),
    .B2(_00948_),
    .X(_01081_));
 sky130_fd_sc_hd__o21a_1 _22139_ (.A1(_00947_),
    .A2(_00959_),
    .B1(_00963_),
    .X(_01082_));
 sky130_fd_sc_hd__nand3_2 _22140_ (.A(_01075_),
    .B(_01077_),
    .C(_01081_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand3_2 _22141_ (.A(_01078_),
    .B(_01079_),
    .C(_01082_),
    .Y(_01084_));
 sky130_fd_sc_hd__a32oi_2 _22142_ (.A1(_00945_),
    .A2(_00964_),
    .A3(_00965_),
    .B1(_00969_),
    .B2(_00943_),
    .Y(_01085_));
 sky130_fd_sc_hd__a21oi_1 _22143_ (.A1(_01083_),
    .A2(_01084_),
    .B1(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__a21o_1 _22144_ (.A1(_01083_),
    .A2(_01084_),
    .B1(_01085_),
    .X(_01087_));
 sky130_fd_sc_hd__o211a_1 _22145_ (.A1(_00968_),
    .A2(_00972_),
    .B1(_01083_),
    .C1(_01084_),
    .X(_01088_));
 sky130_fd_sc_hd__o211ai_2 _22146_ (.A1(_00968_),
    .A2(_00972_),
    .B1(_01083_),
    .C1(_01084_),
    .Y(_01089_));
 sky130_fd_sc_hd__a2bb2oi_1 _22147_ (.A1_N(_00990_),
    .A2_N(_00994_),
    .B1(_00981_),
    .B2(_00992_),
    .Y(_01090_));
 sky130_fd_sc_hd__nand2_1 _22148_ (.A(_02131_),
    .B(net57),
    .Y(_01092_));
 sky130_fd_sc_hd__and4_1 _22149_ (.A(_02131_),
    .B(net19),
    .C(net56),
    .D(net57),
    .X(_01093_));
 sky130_fd_sc_hd__o22a_1 _22150_ (.A1(net18),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02142_),
    .X(_01094_));
 sky130_fd_sc_hd__nor2_1 _22151_ (.A(_01093_),
    .B(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__o31ai_1 _22152_ (.A1(_02142_),
    .A2(_02207_),
    .A3(_00987_),
    .B1(_00985_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_2 _22153_ (.A(net53),
    .B(net22),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_1 _22154_ (.A(net52),
    .B(net22),
    .Y(_01098_));
 sky130_fd_sc_hd__a22oi_2 _22155_ (.A1(net21),
    .A2(net53),
    .B1(net22),
    .B2(net52),
    .Y(_01099_));
 sky130_fd_sc_hd__a22o_1 _22156_ (.A1(net21),
    .A2(net53),
    .B1(net22),
    .B2(net52),
    .X(_01100_));
 sky130_fd_sc_hd__nand3_1 _22157_ (.A(_01098_),
    .B(net53),
    .C(net21),
    .Y(_01101_));
 sky130_fd_sc_hd__nand3_1 _22158_ (.A(_00984_),
    .B(net22),
    .C(net52),
    .Y(_01103_));
 sky130_fd_sc_hd__o2111ai_2 _22159_ (.A1(_00986_),
    .A2(_01097_),
    .B1(net20),
    .C1(net54),
    .D1(_01100_),
    .Y(_01104_));
 sky130_fd_sc_hd__o211ai_2 _22160_ (.A1(_02163_),
    .A2(_02207_),
    .B1(_01101_),
    .C1(_01103_),
    .Y(_01105_));
 sky130_fd_sc_hd__a21o_1 _22161_ (.A1(_01104_),
    .A2(_01105_),
    .B1(_01096_),
    .X(_01106_));
 sky130_fd_sc_hd__and3_1 _22162_ (.A(_01096_),
    .B(_01104_),
    .C(_01105_),
    .X(_01107_));
 sky130_fd_sc_hd__nand3_1 _22163_ (.A(_01096_),
    .B(_01104_),
    .C(_01105_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand3_1 _22164_ (.A(_01106_),
    .B(_01108_),
    .C(_01095_),
    .Y(_01109_));
 sky130_fd_sc_hd__a21o_1 _22165_ (.A1(_01106_),
    .A2(_01108_),
    .B1(_01095_),
    .X(_01110_));
 sky130_fd_sc_hd__a21bo_1 _22166_ (.A1(_01106_),
    .A2(_01108_),
    .B1_N(_01095_),
    .X(_01111_));
 sky130_fd_sc_hd__o211ai_1 _22167_ (.A1(_01093_),
    .A2(_01094_),
    .B1(_01106_),
    .C1(_01108_),
    .Y(_01112_));
 sky130_fd_sc_hd__nand3b_4 _22168_ (.A_N(_01090_),
    .B(_01109_),
    .C(_01110_),
    .Y(_01114_));
 sky130_fd_sc_hd__nand3_1 _22169_ (.A(_01111_),
    .B(_01112_),
    .C(_01090_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand3_4 _22170_ (.A(_01114_),
    .B(_01115_),
    .C(_00979_),
    .Y(_01116_));
 sky130_fd_sc_hd__a21o_1 _22171_ (.A1(_01114_),
    .A2(_01115_),
    .B1(_00979_),
    .X(_01117_));
 sky130_fd_sc_hd__nand2_1 _22172_ (.A(_01116_),
    .B(_01117_),
    .Y(_01118_));
 sky130_fd_sc_hd__o21ai_2 _22173_ (.A1(_01086_),
    .A2(_01088_),
    .B1(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__and4_1 _22174_ (.A(_01087_),
    .B(_01089_),
    .C(_01116_),
    .D(_01117_),
    .X(_01120_));
 sky130_fd_sc_hd__nand4_2 _22175_ (.A(_01087_),
    .B(_01089_),
    .C(_01116_),
    .D(_01117_),
    .Y(_01121_));
 sky130_fd_sc_hd__a21oi_1 _22176_ (.A1(_01119_),
    .A2(_01121_),
    .B1(_01053_),
    .Y(_01122_));
 sky130_fd_sc_hd__a21o_1 _22177_ (.A1(_01119_),
    .A2(_01121_),
    .B1(_01053_),
    .X(_01123_));
 sky130_fd_sc_hd__o211a_1 _22178_ (.A1(_00799_),
    .A2(_00930_),
    .B1(_01119_),
    .C1(_01121_),
    .X(_01125_));
 sky130_fd_sc_hd__o211ai_1 _22179_ (.A1(_00799_),
    .A2(_00930_),
    .B1(_01119_),
    .C1(_01121_),
    .Y(_01126_));
 sky130_fd_sc_hd__nand3b_1 _22180_ (.A_N(_01051_),
    .B(_01123_),
    .C(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__o21ai_1 _22181_ (.A1(_01122_),
    .A2(_01125_),
    .B1(_01051_),
    .Y(_01128_));
 sky130_fd_sc_hd__o21bai_1 _22182_ (.A1(_01122_),
    .A2(_01125_),
    .B1_N(_01051_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand3_1 _22183_ (.A(_01051_),
    .B(_01123_),
    .C(_01126_),
    .Y(_01130_));
 sky130_fd_sc_hd__o211ai_1 _22184_ (.A1(_01045_),
    .A2(_01048_),
    .B1(_01127_),
    .C1(_01128_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand3_2 _22185_ (.A(_01129_),
    .B(_01130_),
    .C(_01049_),
    .Y(_01132_));
 sky130_fd_sc_hd__nand2_2 _22186_ (.A(_01131_),
    .B(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__o211ai_4 _22187_ (.A1(_01017_),
    .A2(_01019_),
    .B1(_01133_),
    .C1(_00939_),
    .Y(_01134_));
 sky130_fd_sc_hd__a21oi_2 _22188_ (.A1(_00939_),
    .A2(_01020_),
    .B1(_01133_),
    .Y(_01136_));
 sky130_fd_sc_hd__a21o_1 _22189_ (.A1(_00939_),
    .A2(_01020_),
    .B1(_01133_),
    .X(_01137_));
 sky130_fd_sc_hd__nand2_1 _22190_ (.A(_01010_),
    .B(_01014_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand3_1 _22191_ (.A(_01134_),
    .B(_01137_),
    .C(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__a21o_1 _22192_ (.A1(_01134_),
    .A2(_01137_),
    .B1(_01138_),
    .X(_01140_));
 sky130_fd_sc_hd__a31o_1 _22193_ (.A1(_01018_),
    .A2(_01020_),
    .A3(_01021_),
    .B1(_01027_),
    .X(_01141_));
 sky130_fd_sc_hd__a221o_1 _22194_ (.A1(_01027_),
    .A2(_01023_),
    .B1(_01140_),
    .B2(_01139_),
    .C1(_01024_),
    .X(_01142_));
 sky130_fd_sc_hd__nand4_2 _22195_ (.A(_01023_),
    .B(_01139_),
    .C(_01140_),
    .D(_01141_),
    .Y(_01143_));
 sky130_fd_sc_hd__a21boi_2 _22196_ (.A1(_00855_),
    .A2(_00999_),
    .B1_N(_00998_),
    .Y(_01144_));
 sky130_fd_sc_hd__a21oi_1 _22197_ (.A1(_01142_),
    .A2(_01143_),
    .B1(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand2_1 _22198_ (.A(_01142_),
    .B(_01144_),
    .Y(_01147_));
 sky130_fd_sc_hd__and3_1 _22199_ (.A(_01142_),
    .B(_01143_),
    .C(_01144_),
    .X(_01148_));
 sky130_fd_sc_hd__a21oi_1 _22200_ (.A1(_01032_),
    .A2(_01035_),
    .B1(_01033_),
    .Y(_01149_));
 sky130_fd_sc_hd__o21ai_1 _22201_ (.A1(_01145_),
    .A2(_01148_),
    .B1(_01149_),
    .Y(_01150_));
 sky130_fd_sc_hd__or2_1 _22202_ (.A(_01149_),
    .B(_01145_),
    .X(_01151_));
 sky130_fd_sc_hd__o21a_1 _22203_ (.A1(_01148_),
    .A2(_01151_),
    .B1(_01150_),
    .X(_01152_));
 sky130_fd_sc_hd__o2111a_1 _22204_ (.A1(_01041_),
    .A2(_01038_),
    .B1(_00919_),
    .C1(_00916_),
    .D1(_01040_),
    .X(_01153_));
 sky130_fd_sc_hd__o2111ai_1 _22205_ (.A1(_01041_),
    .A2(_01038_),
    .B1(_00919_),
    .C1(_00916_),
    .D1(_01040_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand4_1 _22206_ (.A(_00626_),
    .B(_00627_),
    .C(_00776_),
    .D(_00777_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _22207_ (.A(_01154_),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__and2_1 _22208_ (.A(_00631_),
    .B(_01156_),
    .X(_01158_));
 sky130_fd_sc_hd__o221ai_4 _22209_ (.A1(_00019_),
    .A2(_00020_),
    .B1(_00023_),
    .B2(_09243_),
    .C1(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__a32o_1 _22210_ (.A1(_00912_),
    .A2(_01036_),
    .A3(_01039_),
    .B1(_00918_),
    .B2(_01040_),
    .X(_01160_));
 sky130_fd_sc_hd__a31o_1 _22211_ (.A1(_01153_),
    .A2(_00921_),
    .A3(_00776_),
    .B1(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__a21oi_2 _22212_ (.A1(_00630_),
    .A2(_01156_),
    .B1(_01161_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2_1 _22213_ (.A(_01159_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__xor2_1 _22214_ (.A(_01152_),
    .B(_01163_),
    .X(net116));
 sky130_fd_sc_hd__a32oi_4 _22215_ (.A1(_00939_),
    .A2(_01020_),
    .A3(_01133_),
    .B1(_01010_),
    .B2(_01014_),
    .Y(_01164_));
 sky130_fd_sc_hd__a31o_1 _22216_ (.A1(_01129_),
    .A2(_01130_),
    .A3(_01049_),
    .B1(_01045_),
    .X(_01165_));
 sky130_fd_sc_hd__a31o_1 _22217_ (.A1(_01087_),
    .A2(_01116_),
    .A3(_01117_),
    .B1(_01088_),
    .X(_01166_));
 sky130_fd_sc_hd__a21boi_1 _22218_ (.A1(_01077_),
    .A2(_01081_),
    .B1_N(_01075_),
    .Y(_01168_));
 sky130_fd_sc_hd__o21ai_1 _22219_ (.A1(_01082_),
    .A2(_01076_),
    .B1(_01075_),
    .Y(_01169_));
 sky130_fd_sc_hd__a21o_1 _22220_ (.A1(_01054_),
    .A2(_01065_),
    .B1(_01067_),
    .X(_01170_));
 sky130_fd_sc_hd__nand2_1 _22221_ (.A(net51),
    .B(net25),
    .Y(_01171_));
 sky130_fd_sc_hd__o211ai_2 _22222_ (.A1(_02152_),
    .A2(_02251_),
    .B1(_01057_),
    .C1(_01060_),
    .Y(_01172_));
 sky130_fd_sc_hd__o21bai_1 _22223_ (.A1(_01056_),
    .A2(_01059_),
    .B1_N(_01171_),
    .Y(_01173_));
 sky130_fd_sc_hd__o22ai_2 _22224_ (.A1(_02152_),
    .A2(_02251_),
    .B1(_01056_),
    .B2(_01059_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand4_2 _22225_ (.A(_01057_),
    .B(_01060_),
    .C(net51),
    .D(net25),
    .Y(_01175_));
 sky130_fd_sc_hd__nand3_4 _22226_ (.A(_01173_),
    .B(_00950_),
    .C(_01172_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand3_4 _22227_ (.A(_00951_),
    .B(_01174_),
    .C(_01175_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_2 _22228_ (.A(_01176_),
    .B(_01177_),
    .Y(_01179_));
 sky130_fd_sc_hd__o21a_1 _22229_ (.A1(_02152_),
    .A2(_02218_),
    .B1(_01060_),
    .X(_01180_));
 sky130_fd_sc_hd__and3_1 _22230_ (.A(_01057_),
    .B(net24),
    .C(net51),
    .X(_01181_));
 sky130_fd_sc_hd__o211ai_4 _22231_ (.A1(_01059_),
    .A2(_01181_),
    .B1(_01177_),
    .C1(_01176_),
    .Y(_01182_));
 sky130_fd_sc_hd__o2bb2ai_1 _22232_ (.A1_N(_01176_),
    .A2_N(_01177_),
    .B1(_01180_),
    .B2(_01056_),
    .Y(_01183_));
 sky130_fd_sc_hd__o2bb2ai_1 _22233_ (.A1_N(_01176_),
    .A2_N(_01177_),
    .B1(_01181_),
    .B2(_01059_),
    .Y(_01184_));
 sky130_fd_sc_hd__o2111ai_1 _22234_ (.A1(_01055_),
    .A2(_01056_),
    .B1(_01060_),
    .C1(_01176_),
    .D1(_01177_),
    .Y(_01185_));
 sky130_fd_sc_hd__o211ai_4 _22235_ (.A1(_00366_),
    .A2(_00792_),
    .B1(_01182_),
    .C1(_01183_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand3_2 _22236_ (.A(_01184_),
    .B(_01185_),
    .C(_00945_),
    .Y(_01187_));
 sky130_fd_sc_hd__a21oi_1 _22237_ (.A1(_01186_),
    .A2(_01187_),
    .B1(_01170_),
    .Y(_01188_));
 sky130_fd_sc_hd__a21o_1 _22238_ (.A1(_01186_),
    .A2(_01187_),
    .B1(_01170_),
    .X(_01190_));
 sky130_fd_sc_hd__o211a_1 _22239_ (.A1(_01067_),
    .A2(_01068_),
    .B1(_01186_),
    .C1(_01187_),
    .X(_01191_));
 sky130_fd_sc_hd__o211ai_2 _22240_ (.A1(_01067_),
    .A2(_01068_),
    .B1(_01186_),
    .C1(_01187_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand3_2 _22241_ (.A(_01169_),
    .B(_01190_),
    .C(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__o221a_1 _22242_ (.A1(_01076_),
    .A2(_01082_),
    .B1(_01188_),
    .B2(_01191_),
    .C1(_01075_),
    .X(_01194_));
 sky130_fd_sc_hd__o21ai_2 _22243_ (.A1(_01188_),
    .A2(_01191_),
    .B1(_01168_),
    .Y(_01195_));
 sky130_fd_sc_hd__a21oi_1 _22244_ (.A1(_01106_),
    .A2(_01095_),
    .B1(_01107_),
    .Y(_01196_));
 sky130_fd_sc_hd__a21o_1 _22245_ (.A1(_01106_),
    .A2(_01095_),
    .B1(_01107_),
    .X(_01197_));
 sky130_fd_sc_hd__and4_1 _22246_ (.A(_02142_),
    .B(net20),
    .C(net56),
    .D(net57),
    .X(_01198_));
 sky130_fd_sc_hd__o22a_1 _22247_ (.A1(net19),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02163_),
    .X(_01199_));
 sky130_fd_sc_hd__nor2_1 _22248_ (.A(_01198_),
    .B(_01199_),
    .Y(_01201_));
 sky130_fd_sc_hd__o32ai_4 _22249_ (.A1(_02163_),
    .A2(_02207_),
    .A3(_01099_),
    .B1(_01097_),
    .B2(_00986_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _22250_ (.A(net53),
    .B(net24),
    .Y(_01203_));
 sky130_fd_sc_hd__nand2_1 _22251_ (.A(net52),
    .B(net24),
    .Y(_01204_));
 sky130_fd_sc_hd__and4_1 _22252_ (.A(net52),
    .B(net53),
    .C(net22),
    .D(net24),
    .X(_01205_));
 sky130_fd_sc_hd__a22o_1 _22253_ (.A1(net53),
    .A2(net22),
    .B1(net24),
    .B2(net52),
    .X(_01206_));
 sky130_fd_sc_hd__nand3_1 _22254_ (.A(_01204_),
    .B(net22),
    .C(net53),
    .Y(_01207_));
 sky130_fd_sc_hd__nand3_1 _22255_ (.A(_01097_),
    .B(net24),
    .C(net52),
    .Y(_01208_));
 sky130_fd_sc_hd__o2111ai_4 _22256_ (.A1(_01098_),
    .A2(_01203_),
    .B1(net21),
    .C1(net54),
    .D1(_01206_),
    .Y(_01209_));
 sky130_fd_sc_hd__o211ai_2 _22257_ (.A1(_02185_),
    .A2(_02207_),
    .B1(_01207_),
    .C1(_01208_),
    .Y(_01210_));
 sky130_fd_sc_hd__a21oi_1 _22258_ (.A1(_01209_),
    .A2(_01210_),
    .B1(_01202_),
    .Y(_01212_));
 sky130_fd_sc_hd__a21o_1 _22259_ (.A1(_01209_),
    .A2(_01210_),
    .B1(_01202_),
    .X(_01213_));
 sky130_fd_sc_hd__and3_1 _22260_ (.A(_01202_),
    .B(_01209_),
    .C(_01210_),
    .X(_01214_));
 sky130_fd_sc_hd__nand3_2 _22261_ (.A(_01202_),
    .B(_01209_),
    .C(_01210_),
    .Y(_01215_));
 sky130_fd_sc_hd__nand3_2 _22262_ (.A(_01213_),
    .B(_01215_),
    .C(_01201_),
    .Y(_01216_));
 sky130_fd_sc_hd__a21o_1 _22263_ (.A1(_01213_),
    .A2(_01215_),
    .B1(_01201_),
    .X(_01217_));
 sky130_fd_sc_hd__o21ai_1 _22264_ (.A1(_01212_),
    .A2(_01214_),
    .B1(_01201_),
    .Y(_01218_));
 sky130_fd_sc_hd__o211ai_1 _22265_ (.A1(_01198_),
    .A2(_01199_),
    .B1(_01213_),
    .C1(_01215_),
    .Y(_01219_));
 sky130_fd_sc_hd__nand3_4 _22266_ (.A(_01197_),
    .B(_01216_),
    .C(_01217_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand3_2 _22267_ (.A(_01218_),
    .B(_01219_),
    .C(_01196_),
    .Y(_01221_));
 sky130_fd_sc_hd__and3_1 _22268_ (.A(_01220_),
    .B(_01221_),
    .C(_01093_),
    .X(_01223_));
 sky130_fd_sc_hd__nand3_1 _22269_ (.A(_01220_),
    .B(_01221_),
    .C(_01093_),
    .Y(_01224_));
 sky130_fd_sc_hd__a21oi_1 _22270_ (.A1(_01220_),
    .A2(_01221_),
    .B1(_01093_),
    .Y(_01225_));
 sky130_fd_sc_hd__a21boi_2 _22271_ (.A1(_01220_),
    .A2(_01221_),
    .B1_N(_01093_),
    .Y(_01226_));
 sky130_fd_sc_hd__o311a_1 _22272_ (.A1(_02142_),
    .A2(_02229_),
    .A3(_01092_),
    .B1(_01220_),
    .C1(_01221_),
    .X(_01227_));
 sky130_fd_sc_hd__o2bb2ai_1 _22273_ (.A1_N(_01193_),
    .A2_N(_01195_),
    .B1(_01226_),
    .B2(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__o211ai_1 _22274_ (.A1(_01223_),
    .A2(_01225_),
    .B1(_01193_),
    .C1(_01195_),
    .Y(_01229_));
 sky130_fd_sc_hd__o2bb2ai_2 _22275_ (.A1_N(_01193_),
    .A2_N(_01195_),
    .B1(_01223_),
    .B2(_01225_),
    .Y(_01230_));
 sky130_fd_sc_hd__o21ai_2 _22276_ (.A1(_01226_),
    .A2(_01227_),
    .B1(_01193_),
    .Y(_01231_));
 sky130_fd_sc_hd__o211ai_1 _22277_ (.A1(_01226_),
    .A2(_01227_),
    .B1(_01193_),
    .C1(_01195_),
    .Y(_01232_));
 sky130_fd_sc_hd__a21oi_1 _22278_ (.A1(_01230_),
    .A2(_01232_),
    .B1(_01053_),
    .Y(_01234_));
 sky130_fd_sc_hd__nand4_2 _22279_ (.A(_00800_),
    .B(_00931_),
    .C(_01228_),
    .D(_01229_),
    .Y(_01235_));
 sky130_fd_sc_hd__o221a_1 _22280_ (.A1(_00799_),
    .A2(_00930_),
    .B1(_01194_),
    .B2(_01231_),
    .C1(_01230_),
    .X(_01236_));
 sky130_fd_sc_hd__o221ai_4 _22281_ (.A1(_00799_),
    .A2(_00930_),
    .B1(_01194_),
    .B2(_01231_),
    .C1(_01230_),
    .Y(_01237_));
 sky130_fd_sc_hd__a21oi_2 _22282_ (.A1(_01235_),
    .A2(_01237_),
    .B1(_01166_),
    .Y(_01238_));
 sky130_fd_sc_hd__o22ai_1 _22283_ (.A1(_01088_),
    .A2(_01120_),
    .B1(_01234_),
    .B2(_01236_),
    .Y(_01239_));
 sky130_fd_sc_hd__o2111ai_1 _22284_ (.A1(_01118_),
    .A2(_01086_),
    .B1(_01089_),
    .C1(_01235_),
    .D1(_01237_),
    .Y(_01240_));
 sky130_fd_sc_hd__a31o_1 _22285_ (.A1(_01166_),
    .A2(_01235_),
    .A3(_01237_),
    .B1(_01050_),
    .X(_01241_));
 sky130_fd_sc_hd__o211ai_2 _22286_ (.A1(_01045_),
    .A2(_01048_),
    .B1(_01239_),
    .C1(_01240_),
    .Y(_01242_));
 sky130_fd_sc_hd__o21ai_1 _22287_ (.A1(_01238_),
    .A2(_01241_),
    .B1(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__o211ai_4 _22288_ (.A1(_01238_),
    .A2(_01241_),
    .B1(_01242_),
    .C1(_01165_),
    .Y(_01245_));
 sky130_fd_sc_hd__o211ai_2 _22289_ (.A1(_10888_),
    .A2(_00933_),
    .B1(_01132_),
    .C1(_01243_),
    .Y(_01246_));
 sky130_fd_sc_hd__a21oi_1 _22290_ (.A1(_01051_),
    .A2(_01123_),
    .B1(_01125_),
    .Y(_01247_));
 sky130_fd_sc_hd__a21bo_1 _22291_ (.A1(_01245_),
    .A2(_01246_),
    .B1_N(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__a31o_1 _22292_ (.A1(_01046_),
    .A2(_01132_),
    .A3(_01243_),
    .B1(_01247_),
    .X(_01249_));
 sky130_fd_sc_hd__nand3b_2 _22293_ (.A_N(_01247_),
    .B(_01246_),
    .C(_01245_),
    .Y(_01250_));
 sky130_fd_sc_hd__a221oi_4 _22294_ (.A1(_01134_),
    .A2(_01138_),
    .B1(_01248_),
    .B2(_01250_),
    .C1(_01136_),
    .Y(_01251_));
 sky130_fd_sc_hd__o211ai_4 _22295_ (.A1(_01136_),
    .A2(_01164_),
    .B1(_01248_),
    .C1(_01250_),
    .Y(_01252_));
 sky130_fd_sc_hd__inv_2 _22296_ (.A(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hd__a211oi_1 _22297_ (.A1(_01114_),
    .A2(_01116_),
    .B1(_01251_),
    .C1(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__o211a_1 _22298_ (.A1(_01251_),
    .A2(_01253_),
    .B1(_01114_),
    .C1(_01116_),
    .X(_01256_));
 sky130_fd_sc_hd__o211a_1 _22299_ (.A1(_01254_),
    .A2(_01256_),
    .B1(_01143_),
    .C1(_01147_),
    .X(_01257_));
 sky130_fd_sc_hd__inv_2 _22300_ (.A(_01257_),
    .Y(_01258_));
 sky130_fd_sc_hd__a211oi_1 _22301_ (.A1(_01143_),
    .A2(_01147_),
    .B1(_01254_),
    .C1(_01256_),
    .Y(_01259_));
 sky130_fd_sc_hd__inv_2 _22302_ (.A(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__nor2_1 _22303_ (.A(_01257_),
    .B(_01259_),
    .Y(_01261_));
 sky130_fd_sc_hd__a2bb2o_1 _22304_ (.A1_N(_01148_),
    .A2_N(_01151_),
    .B1(_01152_),
    .B2(_01163_),
    .X(_01262_));
 sky130_fd_sc_hd__xor2_1 _22305_ (.A(_01261_),
    .B(_01262_),
    .X(net117));
 sky130_fd_sc_hd__a31oi_2 _22306_ (.A1(_01197_),
    .A2(_01216_),
    .A3(_01217_),
    .B1(_01223_),
    .Y(_01263_));
 sky130_fd_sc_hd__nand2_1 _22307_ (.A(_01177_),
    .B(_01182_),
    .Y(_01264_));
 sky130_fd_sc_hd__and3_1 _22308_ (.A(_01057_),
    .B(net25),
    .C(net51),
    .X(_01266_));
 sky130_fd_sc_hd__o31a_2 _22309_ (.A1(_02152_),
    .A2(_02251_),
    .A3(_01056_),
    .B1(_01060_),
    .X(_01267_));
 sky130_fd_sc_hd__o211ai_2 _22310_ (.A1(_01059_),
    .A2(_01266_),
    .B1(_01177_),
    .C1(_01176_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand2_1 _22311_ (.A(_01179_),
    .B(_01267_),
    .Y(_01269_));
 sky130_fd_sc_hd__o2bb2ai_2 _22312_ (.A1_N(_01176_),
    .A2_N(_01177_),
    .B1(_01266_),
    .B2(_01059_),
    .Y(_01270_));
 sky130_fd_sc_hd__o2111ai_4 _22313_ (.A1(_01171_),
    .A2(_01056_),
    .B1(_01060_),
    .C1(_01176_),
    .D1(_01177_),
    .Y(_01271_));
 sky130_fd_sc_hd__o211ai_2 _22314_ (.A1(_00366_),
    .A2(_00792_),
    .B1(_01268_),
    .C1(_01269_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand4_4 _22315_ (.A(_00367_),
    .B(_00793_),
    .C(_01270_),
    .D(_01271_),
    .Y(_01273_));
 sky130_fd_sc_hd__a21o_1 _22316_ (.A1(_01270_),
    .A2(_01271_),
    .B1(_00946_),
    .X(_01274_));
 sky130_fd_sc_hd__o211ai_1 _22317_ (.A1(_00366_),
    .A2(_00792_),
    .B1(_01270_),
    .C1(_01271_),
    .Y(_01275_));
 sky130_fd_sc_hd__nand3_1 _22318_ (.A(_01264_),
    .B(_01274_),
    .C(_01275_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand4_1 _22319_ (.A(_01177_),
    .B(_01182_),
    .C(_01272_),
    .D(_01273_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand4_2 _22320_ (.A(_01186_),
    .B(_01192_),
    .C(_01277_),
    .D(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__o21ai_2 _22321_ (.A1(_01267_),
    .A2(_01179_),
    .B1(_01177_),
    .Y(_01280_));
 sky130_fd_sc_hd__a31o_1 _22322_ (.A1(_00945_),
    .A2(_01270_),
    .A3(_01271_),
    .B1(_01264_),
    .X(_01281_));
 sky130_fd_sc_hd__a22oi_2 _22323_ (.A1(_01177_),
    .A2(_01268_),
    .B1(_01272_),
    .B2(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__a22o_2 _22324_ (.A1(_01177_),
    .A2(_01268_),
    .B1(_01272_),
    .B2(_01281_),
    .X(_01283_));
 sky130_fd_sc_hd__nand2_1 _22325_ (.A(net21),
    .B(net56),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2_1 _22326_ (.A(_02163_),
    .B(net57),
    .Y(_01285_));
 sky130_fd_sc_hd__and4_1 _22327_ (.A(_02163_),
    .B(net21),
    .C(net56),
    .D(net57),
    .X(_01286_));
 sky130_fd_sc_hd__o22a_1 _22328_ (.A1(net20),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02185_),
    .X(_01288_));
 sky130_fd_sc_hd__nor2_1 _22329_ (.A(_01286_),
    .B(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__or2_1 _22330_ (.A(_01286_),
    .B(_01288_),
    .X(_01290_));
 sky130_fd_sc_hd__a31o_1 _22331_ (.A1(_01206_),
    .A2(net54),
    .A3(net21),
    .B1(_01205_),
    .X(_01291_));
 sky130_fd_sc_hd__nand2_1 _22332_ (.A(net22),
    .B(net54),
    .Y(_01292_));
 sky130_fd_sc_hd__nand3_4 _22333_ (.A(net52),
    .B(net53),
    .C(net25),
    .Y(_01293_));
 sky130_fd_sc_hd__and4_1 _22334_ (.A(net52),
    .B(net53),
    .C(net24),
    .D(net25),
    .X(_01294_));
 sky130_fd_sc_hd__nand4_1 _22335_ (.A(net52),
    .B(net53),
    .C(net24),
    .D(net25),
    .Y(_01295_));
 sky130_fd_sc_hd__a22oi_2 _22336_ (.A1(net53),
    .A2(net24),
    .B1(net25),
    .B2(net52),
    .Y(_01296_));
 sky130_fd_sc_hd__nand4b_2 _22337_ (.A_N(_01296_),
    .B(net54),
    .C(net22),
    .D(_01295_),
    .Y(_01297_));
 sky130_fd_sc_hd__o22ai_2 _22338_ (.A1(_02196_),
    .A2(_02207_),
    .B1(_01294_),
    .B2(_01296_),
    .Y(_01299_));
 sky130_fd_sc_hd__a21oi_1 _22339_ (.A1(_01297_),
    .A2(_01299_),
    .B1(_01291_),
    .Y(_01300_));
 sky130_fd_sc_hd__a21o_1 _22340_ (.A1(_01297_),
    .A2(_01299_),
    .B1(_01291_),
    .X(_01301_));
 sky130_fd_sc_hd__and3_1 _22341_ (.A(_01291_),
    .B(_01297_),
    .C(_01299_),
    .X(_01302_));
 sky130_fd_sc_hd__nand3_1 _22342_ (.A(_01291_),
    .B(_01297_),
    .C(_01299_),
    .Y(_01303_));
 sky130_fd_sc_hd__a21oi_1 _22343_ (.A1(_01301_),
    .A2(_01303_),
    .B1(_01290_),
    .Y(_01304_));
 sky130_fd_sc_hd__o21ai_1 _22344_ (.A1(_01300_),
    .A2(_01302_),
    .B1(_01289_),
    .Y(_01305_));
 sky130_fd_sc_hd__o211a_1 _22345_ (.A1(_01286_),
    .A2(_01288_),
    .B1(_01301_),
    .C1(_01303_),
    .X(_01306_));
 sky130_fd_sc_hd__o211ai_1 _22346_ (.A1(_01286_),
    .A2(_01288_),
    .B1(_01301_),
    .C1(_01303_),
    .Y(_01307_));
 sky130_fd_sc_hd__o2bb2ai_1 _22347_ (.A1_N(_01215_),
    .A2_N(_01216_),
    .B1(_01304_),
    .B2(_01306_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand4_1 _22348_ (.A(_01215_),
    .B(_01216_),
    .C(_01305_),
    .D(_01307_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand3_2 _22349_ (.A(_01308_),
    .B(_01310_),
    .C(_01198_),
    .Y(_01311_));
 sky130_fd_sc_hd__a21o_1 _22350_ (.A1(_01308_),
    .A2(_01310_),
    .B1(_01198_),
    .X(_01312_));
 sky130_fd_sc_hd__a22o_1 _22351_ (.A1(_01279_),
    .A2(_01283_),
    .B1(_01311_),
    .B2(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__nand4_2 _22352_ (.A(_01279_),
    .B(_01283_),
    .C(_01311_),
    .D(_01312_),
    .Y(_01314_));
 sky130_fd_sc_hd__a21oi_1 _22353_ (.A1(_01313_),
    .A2(_01314_),
    .B1(_01053_),
    .Y(_01315_));
 sky130_fd_sc_hd__a21o_1 _22354_ (.A1(_01313_),
    .A2(_01314_),
    .B1(_01053_),
    .X(_01316_));
 sky130_fd_sc_hd__o211a_1 _22355_ (.A1(_00799_),
    .A2(_00930_),
    .B1(_01313_),
    .C1(_01314_),
    .X(_01317_));
 sky130_fd_sc_hd__o211ai_1 _22356_ (.A1(_00799_),
    .A2(_00930_),
    .B1(_01313_),
    .C1(_01314_),
    .Y(_01318_));
 sky130_fd_sc_hd__o21a_1 _22357_ (.A1(_01226_),
    .A2(_01227_),
    .B1(_01195_),
    .X(_01319_));
 sky130_fd_sc_hd__a31o_1 _22358_ (.A1(_01169_),
    .A2(_01190_),
    .A3(_01192_),
    .B1(_01319_),
    .X(_01321_));
 sky130_fd_sc_hd__o21ai_1 _22359_ (.A1(_01315_),
    .A2(_01317_),
    .B1(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hd__nand3b_1 _22360_ (.A_N(_01321_),
    .B(_01318_),
    .C(_01316_),
    .Y(_01323_));
 sky130_fd_sc_hd__o21bai_1 _22361_ (.A1(_01315_),
    .A2(_01317_),
    .B1_N(_01321_),
    .Y(_01324_));
 sky130_fd_sc_hd__nand3_1 _22362_ (.A(_01316_),
    .B(_01318_),
    .C(_01321_),
    .Y(_01325_));
 sky130_fd_sc_hd__o211ai_2 _22363_ (.A1(_01045_),
    .A2(_01048_),
    .B1(_01322_),
    .C1(_01323_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand3_2 _22364_ (.A(_01324_),
    .B(_01325_),
    .C(_01049_),
    .Y(_01327_));
 sky130_fd_sc_hd__o21ai_1 _22365_ (.A1(_01238_),
    .A2(_01241_),
    .B1(_01046_),
    .Y(_01328_));
 sky130_fd_sc_hd__a21oi_1 _22366_ (.A1(_01326_),
    .A2(_01327_),
    .B1(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__a21o_1 _22367_ (.A1(_01326_),
    .A2(_01327_),
    .B1(_01328_),
    .X(_01330_));
 sky130_fd_sc_hd__nand3_1 _22368_ (.A(_01326_),
    .B(_01327_),
    .C(_01328_),
    .Y(_01332_));
 sky130_fd_sc_hd__a31o_1 _22369_ (.A1(_01089_),
    .A2(_01121_),
    .A3(_01237_),
    .B1(_01234_),
    .X(_01333_));
 sky130_fd_sc_hd__a21boi_1 _22370_ (.A1(_01330_),
    .A2(_01332_),
    .B1_N(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__and3b_1 _22371_ (.A_N(_01333_),
    .B(_01332_),
    .C(_01330_),
    .X(_01335_));
 sky130_fd_sc_hd__a211oi_2 _22372_ (.A1(_01245_),
    .A2(_01249_),
    .B1(_01334_),
    .C1(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__o211a_1 _22373_ (.A1(_01334_),
    .A2(_01335_),
    .B1(_01245_),
    .C1(_01249_),
    .X(_01337_));
 sky130_fd_sc_hd__a21oi_1 _22374_ (.A1(_01220_),
    .A2(_01224_),
    .B1(_01337_),
    .Y(_01338_));
 sky130_fd_sc_hd__a21o_1 _22375_ (.A1(_01220_),
    .A2(_01224_),
    .B1(_01337_),
    .X(_01339_));
 sky130_fd_sc_hd__o21ai_1 _22376_ (.A1(_01336_),
    .A2(_01337_),
    .B1(_01263_),
    .Y(_01340_));
 sky130_fd_sc_hd__o21ai_1 _22377_ (.A1(_01336_),
    .A2(_01339_),
    .B1(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__a21o_1 _22378_ (.A1(_01114_),
    .A2(_01116_),
    .B1(_01251_),
    .X(_01343_));
 sky130_fd_sc_hd__nand3_1 _22379_ (.A(_01252_),
    .B(_01341_),
    .C(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__a311o_2 _22380_ (.A1(_01114_),
    .A2(_01116_),
    .A3(_01252_),
    .B1(_01251_),
    .C1(_01341_),
    .X(_01345_));
 sky130_fd_sc_hd__nand2_1 _22381_ (.A(_01344_),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__o21ai_1 _22382_ (.A1(_01148_),
    .A2(_01151_),
    .B1(_01260_),
    .Y(_01347_));
 sky130_fd_sc_hd__o31a_1 _22383_ (.A1(_01148_),
    .A2(_01257_),
    .A3(_01151_),
    .B1(_01260_),
    .X(_01348_));
 sky130_fd_sc_hd__o2111ai_2 _22384_ (.A1(_01151_),
    .A2(_01148_),
    .B1(_01150_),
    .C1(_01258_),
    .D1(_01260_),
    .Y(_01349_));
 sky130_fd_sc_hd__inv_2 _22385_ (.A(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__a22oi_2 _22386_ (.A1(_01258_),
    .A2(_01347_),
    .B1(_01163_),
    .B2(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__xor2_1 _22387_ (.A(_01346_),
    .B(_01351_),
    .X(net118));
 sky130_fd_sc_hd__and2_1 _22388_ (.A(_01308_),
    .B(_01311_),
    .X(_01353_));
 sky130_fd_sc_hd__inv_2 _22389_ (.A(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__o21ai_1 _22390_ (.A1(_01333_),
    .A2(_01329_),
    .B1(_01332_),
    .Y(_01355_));
 sky130_fd_sc_hd__a21o_1 _22391_ (.A1(_01316_),
    .A2(_01321_),
    .B1(_01317_),
    .X(_01356_));
 sky130_fd_sc_hd__a31o_1 _22392_ (.A1(_01279_),
    .A2(_01311_),
    .A3(_01312_),
    .B1(_01282_),
    .X(_01357_));
 sky130_fd_sc_hd__o21ai_1 _22393_ (.A1(_01292_),
    .A2(_01296_),
    .B1(_01295_),
    .Y(_01358_));
 sky130_fd_sc_hd__nand2_1 _22394_ (.A(net54),
    .B(net24),
    .Y(_01359_));
 sky130_fd_sc_hd__o21a_2 _22395_ (.A1(net52),
    .A2(net53),
    .B1(net25),
    .X(_01360_));
 sky130_fd_sc_hd__o2bb2ai_1 _22396_ (.A1_N(_01293_),
    .A2_N(_01360_),
    .B1(_02207_),
    .B2(_02218_),
    .Y(_01361_));
 sky130_fd_sc_hd__nand4_1 _22397_ (.A(_01360_),
    .B(net24),
    .C(net54),
    .D(_01293_),
    .Y(_01362_));
 sky130_fd_sc_hd__a21o_1 _22398_ (.A1(_01293_),
    .A2(_01360_),
    .B1(_01359_),
    .X(_01364_));
 sky130_fd_sc_hd__o211ai_2 _22399_ (.A1(_02207_),
    .A2(_02218_),
    .B1(_01293_),
    .C1(_01360_),
    .Y(_01365_));
 sky130_fd_sc_hd__nand3b_4 _22400_ (.A_N(_01358_),
    .B(_01364_),
    .C(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__and3_1 _22401_ (.A(_01358_),
    .B(_01361_),
    .C(_01362_),
    .X(_01367_));
 sky130_fd_sc_hd__nand3_2 _22402_ (.A(_01358_),
    .B(_01361_),
    .C(_01362_),
    .Y(_01368_));
 sky130_fd_sc_hd__nand2_1 _22403_ (.A(net22),
    .B(net56),
    .Y(_01369_));
 sky130_fd_sc_hd__nand2_1 _22404_ (.A(_02185_),
    .B(net57),
    .Y(_01370_));
 sky130_fd_sc_hd__and4_1 _22405_ (.A(_02185_),
    .B(net22),
    .C(net56),
    .D(net57),
    .X(_01371_));
 sky130_fd_sc_hd__o22a_1 _22406_ (.A1(net21),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02196_),
    .X(_01372_));
 sky130_fd_sc_hd__nor2_2 _22407_ (.A(_01371_),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__a21oi_1 _22408_ (.A1(_01366_),
    .A2(_01368_),
    .B1(_01373_),
    .Y(_01375_));
 sky130_fd_sc_hd__and3_1 _22409_ (.A(_01366_),
    .B(_01368_),
    .C(_01373_),
    .X(_01376_));
 sky130_fd_sc_hd__nand3_2 _22410_ (.A(_01366_),
    .B(_01368_),
    .C(_01373_),
    .Y(_01377_));
 sky130_fd_sc_hd__a21oi_1 _22411_ (.A1(_01301_),
    .A2(_01289_),
    .B1(_01302_),
    .Y(_01378_));
 sky130_fd_sc_hd__o21ai_1 _22412_ (.A1(_01290_),
    .A2(_01300_),
    .B1(_01303_),
    .Y(_01379_));
 sky130_fd_sc_hd__o21ai_1 _22413_ (.A1(_01375_),
    .A2(_01376_),
    .B1(_01378_),
    .Y(_01380_));
 sky130_fd_sc_hd__nand3b_2 _22414_ (.A_N(_01375_),
    .B(_01377_),
    .C(_01379_),
    .Y(_01381_));
 sky130_fd_sc_hd__o2bb2ai_2 _22415_ (.A1_N(_01380_),
    .A2_N(_01381_),
    .B1(_01284_),
    .B2(_01285_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand3_2 _22416_ (.A(_01381_),
    .B(_01286_),
    .C(_01380_),
    .Y(_01383_));
 sky130_fd_sc_hd__nand4_4 _22417_ (.A(_00945_),
    .B(_01177_),
    .C(_01179_),
    .D(_01267_),
    .Y(_01384_));
 sky130_fd_sc_hd__inv_2 _22418_ (.A(_01384_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand4_4 _22419_ (.A(_01283_),
    .B(_01382_),
    .C(_01383_),
    .D(_01384_),
    .Y(_01387_));
 sky130_fd_sc_hd__o2bb2ai_2 _22420_ (.A1_N(_01382_),
    .A2_N(_01383_),
    .B1(_01386_),
    .B2(_01282_),
    .Y(_01388_));
 sky130_fd_sc_hd__a21oi_1 _22421_ (.A1(_01387_),
    .A2(_01388_),
    .B1(_01053_),
    .Y(_01389_));
 sky130_fd_sc_hd__a21o_1 _22422_ (.A1(_01387_),
    .A2(_01388_),
    .B1(_01053_),
    .X(_01390_));
 sky130_fd_sc_hd__and3_1 _22423_ (.A(_01053_),
    .B(_01387_),
    .C(_01388_),
    .X(_01391_));
 sky130_fd_sc_hd__o211ai_2 _22424_ (.A1(_00799_),
    .A2(_00929_),
    .B1(_01387_),
    .C1(_01388_),
    .Y(_01392_));
 sky130_fd_sc_hd__a22o_1 _22425_ (.A1(_01283_),
    .A2(_01314_),
    .B1(_01390_),
    .B2(_01392_),
    .X(_01393_));
 sky130_fd_sc_hd__nand4_1 _22426_ (.A(_01283_),
    .B(_01314_),
    .C(_01390_),
    .D(_01392_),
    .Y(_01394_));
 sky130_fd_sc_hd__o21bai_1 _22427_ (.A1(_01389_),
    .A2(_01391_),
    .B1_N(_01357_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _22428_ (.A(_01357_),
    .B(_01390_),
    .Y(_01397_));
 sky130_fd_sc_hd__o211ai_1 _22429_ (.A1(_01045_),
    .A2(_01048_),
    .B1(_01393_),
    .C1(_01394_),
    .Y(_01398_));
 sky130_fd_sc_hd__o211ai_2 _22430_ (.A1(_01391_),
    .A2(_01397_),
    .B1(_01395_),
    .C1(_01049_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2_1 _22431_ (.A(_01398_),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__a21oi_1 _22432_ (.A1(_01046_),
    .A2(_01327_),
    .B1(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__o311a_1 _22433_ (.A1(_09386_),
    .A2(_10752_),
    .A3(_00933_),
    .B1(_01327_),
    .C1(_01400_),
    .X(_01402_));
 sky130_fd_sc_hd__o211ai_2 _22434_ (.A1(_10888_),
    .A2(_00933_),
    .B1(_01327_),
    .C1(_01400_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand3b_1 _22435_ (.A_N(_01401_),
    .B(_01403_),
    .C(_01356_),
    .Y(_01404_));
 sky130_fd_sc_hd__o21bai_1 _22436_ (.A1(_01401_),
    .A2(_01402_),
    .B1_N(_01356_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand3_1 _22437_ (.A(_01404_),
    .B(_01405_),
    .C(_01355_),
    .Y(_01406_));
 sky130_fd_sc_hd__a21o_1 _22438_ (.A1(_01404_),
    .A2(_01405_),
    .B1(_01355_),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_1 _22439_ (.A(_01354_),
    .B(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__and3_1 _22440_ (.A(_01354_),
    .B(_01406_),
    .C(_01408_),
    .X(_01410_));
 sky130_fd_sc_hd__a31o_1 _22441_ (.A1(_01355_),
    .A2(_01404_),
    .A3(_01405_),
    .B1(_01409_),
    .X(_01411_));
 sky130_fd_sc_hd__a21oi_1 _22442_ (.A1(_01406_),
    .A2(_01408_),
    .B1(_01354_),
    .Y(_01412_));
 sky130_fd_sc_hd__inv_2 _22443_ (.A(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__o21ba_1 _22444_ (.A1(_01263_),
    .A2(_01337_),
    .B1_N(_01336_),
    .X(_01414_));
 sky130_fd_sc_hd__o21a_1 _22445_ (.A1(_01410_),
    .A2(_01412_),
    .B1(_01414_),
    .X(_01415_));
 sky130_fd_sc_hd__o211ai_2 _22446_ (.A1(_01336_),
    .A2(_01338_),
    .B1(_01411_),
    .C1(_01413_),
    .Y(_01416_));
 sky130_fd_sc_hd__nand2b_1 _22447_ (.A_N(_01415_),
    .B(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__a21boi_1 _22448_ (.A1(_01351_),
    .A2(_01345_),
    .B1_N(_01344_),
    .Y(_01419_));
 sky130_fd_sc_hd__xnor2_1 _22449_ (.A(_01417_),
    .B(_01419_),
    .Y(net119));
 sky130_fd_sc_hd__nand2_1 _22450_ (.A(_01381_),
    .B(_01383_),
    .Y(_01420_));
 sky130_fd_sc_hd__a21o_1 _22451_ (.A1(_01403_),
    .A2(_01356_),
    .B1(_01401_),
    .X(_01421_));
 sky130_fd_sc_hd__a211o_4 _22452_ (.A1(_00367_),
    .A2(_00793_),
    .B1(_01177_),
    .C1(_01267_),
    .X(_01422_));
 sky130_fd_sc_hd__inv_2 _22453_ (.A(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _22454_ (.A(_01387_),
    .B(_01422_),
    .Y(_01424_));
 sky130_fd_sc_hd__o32a_1 _22455_ (.A1(_00945_),
    .A2(_01267_),
    .A3(_01177_),
    .B1(_01280_),
    .B2(_01273_),
    .X(_01425_));
 sky130_fd_sc_hd__nand2_1 _22456_ (.A(_01384_),
    .B(_01422_),
    .Y(_01426_));
 sky130_fd_sc_hd__and4_1 _22457_ (.A(_02196_),
    .B(net24),
    .C(net56),
    .D(net57),
    .X(_01427_));
 sky130_fd_sc_hd__o22a_1 _22458_ (.A1(net22),
    .A2(_02240_),
    .B1(_02229_),
    .B2(_02218_),
    .X(_01429_));
 sky130_fd_sc_hd__a22o_1 _22459_ (.A1(net24),
    .A2(net56),
    .B1(_02196_),
    .B2(net57),
    .X(_01430_));
 sky130_fd_sc_hd__nor2_1 _22460_ (.A(_02207_),
    .B(_02251_),
    .Y(_01431_));
 sky130_fd_sc_hd__nand3_1 _22461_ (.A(_01293_),
    .B(net24),
    .C(net54),
    .Y(_01432_));
 sky130_fd_sc_hd__o31a_2 _22462_ (.A1(net52),
    .A2(net53),
    .A3(net54),
    .B1(net25),
    .X(_01433_));
 sky130_fd_sc_hd__o2111ai_4 _22463_ (.A1(net52),
    .A2(net53),
    .B1(net54),
    .C1(net25),
    .D1(_01432_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand4b_4 _22464_ (.A_N(_01427_),
    .B(_01430_),
    .C(_01433_),
    .D(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__a2bb2o_1 _22465_ (.A1_N(_01427_),
    .A2_N(_01429_),
    .B1(_01433_),
    .B2(_01434_),
    .X(_01436_));
 sky130_fd_sc_hd__nand2_1 _22466_ (.A(_01435_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__a221oi_4 _22467_ (.A1(_01373_),
    .A2(_01366_),
    .B1(_01436_),
    .B2(_01435_),
    .C1(_01367_),
    .Y(_01438_));
 sky130_fd_sc_hd__a221o_1 _22468_ (.A1(_01373_),
    .A2(_01366_),
    .B1(_01436_),
    .B2(_01435_),
    .C1(_01367_),
    .X(_01440_));
 sky130_fd_sc_hd__a21oi_2 _22469_ (.A1(_01368_),
    .A2(_01377_),
    .B1(_01437_),
    .Y(_01441_));
 sky130_fd_sc_hd__a21o_1 _22470_ (.A1(_01368_),
    .A2(_01377_),
    .B1(_01437_),
    .X(_01442_));
 sky130_fd_sc_hd__nand3_2 _22471_ (.A(_01442_),
    .B(_01371_),
    .C(_01440_),
    .Y(_01443_));
 sky130_fd_sc_hd__o22ai_4 _22472_ (.A1(_01369_),
    .A2(_01370_),
    .B1(_01438_),
    .B2(_01441_),
    .Y(_01444_));
 sky130_fd_sc_hd__o21ai_1 _22473_ (.A1(_01438_),
    .A2(_01441_),
    .B1(_01371_),
    .Y(_01445_));
 sky130_fd_sc_hd__o211ai_1 _22474_ (.A1(_01369_),
    .A2(_01370_),
    .B1(_01440_),
    .C1(_01442_),
    .Y(_01446_));
 sky130_fd_sc_hd__o2111ai_4 _22475_ (.A1(_01273_),
    .A2(_01280_),
    .B1(_01422_),
    .C1(_01443_),
    .D1(_01444_),
    .Y(_01447_));
 sky130_fd_sc_hd__o211ai_2 _22476_ (.A1(_01386_),
    .A2(_01423_),
    .B1(_01445_),
    .C1(_01446_),
    .Y(_01448_));
 sky130_fd_sc_hd__a21o_1 _22477_ (.A1(_01447_),
    .A2(_01448_),
    .B1(_01053_),
    .X(_01449_));
 sky130_fd_sc_hd__o211ai_4 _22478_ (.A1(_00799_),
    .A2(_00929_),
    .B1(_01447_),
    .C1(_01448_),
    .Y(_01451_));
 sky130_fd_sc_hd__nand3_1 _22479_ (.A(_01424_),
    .B(_01449_),
    .C(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__a21o_1 _22480_ (.A1(_01449_),
    .A2(_01451_),
    .B1(_01424_),
    .X(_01453_));
 sky130_fd_sc_hd__a22o_1 _22481_ (.A1(_01387_),
    .A2(_01422_),
    .B1(_01449_),
    .B2(_01451_),
    .X(_01454_));
 sky130_fd_sc_hd__nand4_1 _22482_ (.A(_01387_),
    .B(_01422_),
    .C(_01449_),
    .D(_01451_),
    .Y(_01455_));
 sky130_fd_sc_hd__o2111ai_2 _22483_ (.A1(_10886_),
    .A2(_00932_),
    .B1(_01046_),
    .C1(_01452_),
    .D1(_01453_),
    .Y(_01456_));
 sky130_fd_sc_hd__o211ai_1 _22484_ (.A1(_01045_),
    .A2(_01048_),
    .B1(_01454_),
    .C1(_01455_),
    .Y(_01457_));
 sky130_fd_sc_hd__nand2_1 _22485_ (.A(_01456_),
    .B(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__a21oi_1 _22486_ (.A1(_01046_),
    .A2(_01399_),
    .B1(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__o211ai_1 _22487_ (.A1(_10888_),
    .A2(_00933_),
    .B1(_01399_),
    .C1(_01458_),
    .Y(_01460_));
 sky130_fd_sc_hd__inv_2 _22488_ (.A(_01460_),
    .Y(_01462_));
 sky130_fd_sc_hd__o211ai_1 _22489_ (.A1(_01459_),
    .A2(_01462_),
    .B1(_01392_),
    .C1(_01397_),
    .Y(_01463_));
 sky130_fd_sc_hd__a211o_1 _22490_ (.A1(_01392_),
    .A2(_01397_),
    .B1(_01459_),
    .C1(_01462_),
    .X(_01464_));
 sky130_fd_sc_hd__a221o_1 _22491_ (.A1(_01403_),
    .A2(_01356_),
    .B1(_01464_),
    .B2(_01463_),
    .C1(_01401_),
    .X(_01465_));
 sky130_fd_sc_hd__nand3_1 _22492_ (.A(_01421_),
    .B(_01463_),
    .C(_01464_),
    .Y(_01466_));
 sky130_fd_sc_hd__and3_1 _22493_ (.A(_01420_),
    .B(_01465_),
    .C(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__a21oi_1 _22494_ (.A1(_01465_),
    .A2(_01466_),
    .B1(_01420_),
    .Y(_01468_));
 sky130_fd_sc_hd__a211o_1 _22495_ (.A1(_01406_),
    .A2(_01409_),
    .B1(_01467_),
    .C1(_01468_),
    .X(_01469_));
 sky130_fd_sc_hd__inv_2 _22496_ (.A(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__o211a_1 _22497_ (.A1(_01467_),
    .A2(_01468_),
    .B1(_01406_),
    .C1(_01409_),
    .X(_01471_));
 sky130_fd_sc_hd__inv_2 _22498_ (.A(_01471_),
    .Y(_01473_));
 sky130_fd_sc_hd__nand3b_1 _22499_ (.A_N(_01417_),
    .B(_01345_),
    .C(_01344_),
    .Y(_01474_));
 sky130_fd_sc_hd__or2_1 _22500_ (.A(_01349_),
    .B(_01474_),
    .X(_01475_));
 sky130_fd_sc_hd__a21oi_1 _22501_ (.A1(_01159_),
    .A2(_01162_),
    .B1(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__o221ai_4 _22502_ (.A1(_01415_),
    .A2(_01345_),
    .B1(_01348_),
    .B2(_01474_),
    .C1(_01416_),
    .Y(_01477_));
 sky130_fd_sc_hd__nor2_1 _22503_ (.A(_01477_),
    .B(_01476_),
    .Y(_01478_));
 sky130_fd_sc_hd__o21a_1 _22504_ (.A1(_01477_),
    .A2(_01476_),
    .B1(_01473_),
    .X(_01479_));
 sky130_fd_sc_hd__nand2_1 _22505_ (.A(_01469_),
    .B(_01473_),
    .Y(_01480_));
 sky130_fd_sc_hd__a22oi_1 _22506_ (.A1(_01478_),
    .A2(_01480_),
    .B1(_01479_),
    .B2(_01469_),
    .Y(net121));
 sky130_fd_sc_hd__o31a_1 _22507_ (.A1(_01369_),
    .A2(_01370_),
    .A3(_01438_),
    .B1(_01442_),
    .X(_01481_));
 sky130_fd_sc_hd__inv_2 _22508_ (.A(_01481_),
    .Y(_01483_));
 sky130_fd_sc_hd__and2b_1 _22509_ (.A_N(_01459_),
    .B(_01464_),
    .X(_01484_));
 sky130_fd_sc_hd__nand2_1 _22510_ (.A(_01451_),
    .B(_01452_),
    .Y(_01485_));
 sky130_fd_sc_hd__o21ai_1 _22511_ (.A1(_10888_),
    .A2(_00933_),
    .B1(_01456_),
    .Y(_01486_));
 sky130_fd_sc_hd__a31o_1 _22512_ (.A1(_01425_),
    .A2(_01443_),
    .A3(_01444_),
    .B1(_01423_),
    .X(_01487_));
 sky130_fd_sc_hd__and4_1 _22513_ (.A(net52),
    .B(net53),
    .C(net54),
    .D(net25),
    .X(_01488_));
 sky130_fd_sc_hd__nand4_4 _22514_ (.A(net52),
    .B(net53),
    .C(net54),
    .D(net25),
    .Y(_01489_));
 sky130_fd_sc_hd__nand2_1 _22515_ (.A(net56),
    .B(net25),
    .Y(_01490_));
 sky130_fd_sc_hd__nand2_1 _22516_ (.A(_02218_),
    .B(net57),
    .Y(_01491_));
 sky130_fd_sc_hd__nand4_4 _22517_ (.A(_02218_),
    .B(net56),
    .C(net57),
    .D(net25),
    .Y(_01492_));
 sky130_fd_sc_hd__a22o_1 _22518_ (.A1(net56),
    .A2(net25),
    .B1(_02218_),
    .B2(net57),
    .X(_01494_));
 sky130_fd_sc_hd__a22oi_4 _22519_ (.A1(_01433_),
    .A2(_01489_),
    .B1(_01492_),
    .B2(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__o2111a_2 _22520_ (.A1(_02207_),
    .A2(_01293_),
    .B1(_01433_),
    .C1(_01492_),
    .D1(_01494_),
    .X(_01496_));
 sky130_fd_sc_hd__o221a_1 _22521_ (.A1(_02207_),
    .A2(_01293_),
    .B1(_01495_),
    .B2(_01496_),
    .C1(_01435_),
    .X(_01497_));
 sky130_fd_sc_hd__o221ai_4 _22522_ (.A1(_02207_),
    .A2(_01293_),
    .B1(_01495_),
    .B2(_01496_),
    .C1(_01435_),
    .Y(_01498_));
 sky130_fd_sc_hd__a211oi_2 _22523_ (.A1(_01435_),
    .A2(_01489_),
    .B1(_01495_),
    .C1(_01496_),
    .Y(_01499_));
 sky130_fd_sc_hd__o21bai_2 _22524_ (.A1(_01497_),
    .A2(_01499_),
    .B1_N(_01427_),
    .Y(_01500_));
 sky130_fd_sc_hd__nand3b_2 _22525_ (.A_N(_01499_),
    .B(_01427_),
    .C(_01498_),
    .Y(_01501_));
 sky130_fd_sc_hd__nand3_2 _22526_ (.A(_01425_),
    .B(_01500_),
    .C(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__a22o_1 _22527_ (.A1(_01384_),
    .A2(_01422_),
    .B1(_01500_),
    .B2(_01501_),
    .X(_01503_));
 sky130_fd_sc_hd__a21o_1 _22528_ (.A1(_01500_),
    .A2(_01501_),
    .B1(_01426_),
    .X(_01505_));
 sky130_fd_sc_hd__o211ai_1 _22529_ (.A1(_01386_),
    .A2(_01423_),
    .B1(_01500_),
    .C1(_01501_),
    .Y(_01506_));
 sky130_fd_sc_hd__o211ai_2 _22530_ (.A1(_00799_),
    .A2(_00929_),
    .B1(_01502_),
    .C1(_01503_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand4_1 _22531_ (.A(_00800_),
    .B(_00931_),
    .C(_01505_),
    .D(_01506_),
    .Y(_01508_));
 sky130_fd_sc_hd__nand3_1 _22532_ (.A(_01503_),
    .B(_01052_),
    .C(_01502_),
    .Y(_01509_));
 sky130_fd_sc_hd__o211ai_1 _22533_ (.A1(_00799_),
    .A2(_00929_),
    .B1(_01505_),
    .C1(_01506_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand3_1 _22534_ (.A(_01487_),
    .B(_01507_),
    .C(_01508_),
    .Y(_01511_));
 sky130_fd_sc_hd__nand4_1 _22535_ (.A(_01422_),
    .B(_01447_),
    .C(_01509_),
    .D(_01510_),
    .Y(_01512_));
 sky130_fd_sc_hd__nand2_1 _22536_ (.A(_01511_),
    .B(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hd__xnor2_1 _22537_ (.A(_01050_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__a21oi_1 _22538_ (.A1(_01046_),
    .A2(_01456_),
    .B1(_01514_),
    .Y(_01516_));
 sky130_fd_sc_hd__xor2_1 _22539_ (.A(_01486_),
    .B(_01514_),
    .X(_01517_));
 sky130_fd_sc_hd__a21oi_1 _22540_ (.A1(_01451_),
    .A2(_01452_),
    .B1(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__xor2_1 _22541_ (.A(_01485_),
    .B(_01517_),
    .X(_01519_));
 sky130_fd_sc_hd__nor2_1 _22542_ (.A(_01484_),
    .B(_01519_),
    .Y(_01520_));
 sky130_fd_sc_hd__nand2_1 _22543_ (.A(_01519_),
    .B(_01484_),
    .Y(_01521_));
 sky130_fd_sc_hd__nand2b_1 _22544_ (.A_N(_01520_),
    .B(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__or3b_1 _22545_ (.A(_01481_),
    .B(_01520_),
    .C_N(_01521_),
    .X(_01523_));
 sky130_fd_sc_hd__nand2_1 _22546_ (.A(_01522_),
    .B(_01481_),
    .Y(_01524_));
 sky130_fd_sc_hd__a21bo_1 _22547_ (.A1(_01420_),
    .A2(_01465_),
    .B1_N(_01466_),
    .X(_01525_));
 sky130_fd_sc_hd__a21oi_1 _22548_ (.A1(_01523_),
    .A2(_01524_),
    .B1(_01525_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand3_1 _22549_ (.A(_01523_),
    .B(_01524_),
    .C(_01525_),
    .Y(_01528_));
 sky130_fd_sc_hd__nand2b_1 _22550_ (.A_N(_01527_),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__o211a_1 _22551_ (.A1(_01471_),
    .A2(_01478_),
    .B1(_01529_),
    .C1(_01469_),
    .X(_01530_));
 sky130_fd_sc_hd__o21ba_1 _22552_ (.A1(_01470_),
    .A2(_01479_),
    .B1_N(_01529_),
    .X(_01531_));
 sky130_fd_sc_hd__nor2_1 _22553_ (.A(_01530_),
    .B(_01531_),
    .Y(net122));
 sky130_fd_sc_hd__or2_1 _22554_ (.A(_01480_),
    .B(_01529_),
    .X(_01532_));
 sky130_fd_sc_hd__o21bai_1 _22555_ (.A1(_01477_),
    .A2(_01476_),
    .B1_N(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__a21o_1 _22556_ (.A1(_01469_),
    .A2(_01528_),
    .B1(_01527_),
    .X(_01534_));
 sky130_fd_sc_hd__a21oi_1 _22557_ (.A1(_01427_),
    .A2(_01498_),
    .B1(_01499_),
    .Y(_01535_));
 sky130_fd_sc_hd__or2_1 _22558_ (.A(_01516_),
    .B(_01518_),
    .X(_01537_));
 sky130_fd_sc_hd__nand2_1 _22559_ (.A(_01507_),
    .B(_01511_),
    .Y(_01538_));
 sky130_fd_sc_hd__a31o_1 _22560_ (.A1(_01049_),
    .A2(_01511_),
    .A3(_01512_),
    .B1(_01045_),
    .X(_01539_));
 sky130_fd_sc_hd__nand2_1 _22561_ (.A(_01422_),
    .B(_01502_),
    .Y(_01540_));
 sky130_fd_sc_hd__a31oi_1 _22562_ (.A1(_01433_),
    .A2(_01492_),
    .A3(_01494_),
    .B1(_01488_),
    .Y(_01541_));
 sky130_fd_sc_hd__o21ai_2 _22563_ (.A1(net25),
    .A2(_02240_),
    .B1(_01490_),
    .Y(_01542_));
 sky130_fd_sc_hd__a21oi_1 _22564_ (.A1(_01433_),
    .A2(_01489_),
    .B1(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21o_1 _22565_ (.A1(_01433_),
    .A2(_01489_),
    .B1(_01542_),
    .X(_01544_));
 sky130_fd_sc_hd__o221a_1 _22566_ (.A1(_02207_),
    .A2(_01293_),
    .B1(_01360_),
    .B2(_01431_),
    .C1(_01542_),
    .X(_01545_));
 sky130_fd_sc_hd__o221ai_2 _22567_ (.A1(_02207_),
    .A2(_01293_),
    .B1(_01431_),
    .B2(_01360_),
    .C1(_01542_),
    .Y(_01546_));
 sky130_fd_sc_hd__o21ai_1 _22568_ (.A1(_01543_),
    .A2(_01545_),
    .B1(_01541_),
    .Y(_01548_));
 sky130_fd_sc_hd__o211ai_2 _22569_ (.A1(_01488_),
    .A2(_01496_),
    .B1(_01544_),
    .C1(_01546_),
    .Y(_01549_));
 sky130_fd_sc_hd__nand3b_1 _22570_ (.A_N(_01492_),
    .B(_01548_),
    .C(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__o2bb2ai_1 _22571_ (.A1_N(_01548_),
    .A2_N(_01549_),
    .B1(_01490_),
    .B2(_01491_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_1 _22572_ (.A(_01550_),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__xor2_1 _22573_ (.A(_01426_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__xor2_1 _22574_ (.A(_01052_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__a21oi_1 _22575_ (.A1(_01422_),
    .A2(_01502_),
    .B1(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__xnor2_1 _22576_ (.A(_01540_),
    .B(_01554_),
    .Y(_01556_));
 sky130_fd_sc_hd__xor2_1 _22577_ (.A(_01049_),
    .B(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__xnor2_1 _22578_ (.A(_01539_),
    .B(_01557_),
    .Y(_01559_));
 sky130_fd_sc_hd__a21o_1 _22579_ (.A1(_01507_),
    .A2(_01511_),
    .B1(_01559_),
    .X(_01560_));
 sky130_fd_sc_hd__xnor2_1 _22580_ (.A(_01538_),
    .B(_01559_),
    .Y(_01561_));
 sky130_fd_sc_hd__o21ai_1 _22581_ (.A1(_01516_),
    .A2(_01518_),
    .B1(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__xnor2_1 _22582_ (.A(_01537_),
    .B(_01561_),
    .Y(_01563_));
 sky130_fd_sc_hd__xor2_1 _22583_ (.A(_01535_),
    .B(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__inv_2 _22584_ (.A(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__a21oi_1 _22585_ (.A1(_01483_),
    .A2(_01521_),
    .B1(_01520_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_1 _22586_ (.A(_01565_),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__or2_1 _22587_ (.A(_01566_),
    .B(_01564_),
    .X(_01568_));
 sky130_fd_sc_hd__nand2_1 _22588_ (.A(_01564_),
    .B(_01566_),
    .Y(_01570_));
 sky130_fd_sc_hd__a22oi_1 _22589_ (.A1(_01568_),
    .A2(_01570_),
    .B1(_01533_),
    .B2(_01534_),
    .Y(_01571_));
 sky130_fd_sc_hd__a22o_1 _22590_ (.A1(_01568_),
    .A2(_01570_),
    .B1(_01533_),
    .B2(_01534_),
    .X(_01572_));
 sky130_fd_sc_hd__and4_1 _22591_ (.A(_01533_),
    .B(_01534_),
    .C(_01568_),
    .D(_01570_),
    .X(_01573_));
 sky130_fd_sc_hd__nor2_1 _22592_ (.A(_01571_),
    .B(_01573_),
    .Y(net123));
 sky130_fd_sc_hd__o21ai_1 _22593_ (.A1(_01535_),
    .A2(_01563_),
    .B1(_01562_),
    .Y(_01574_));
 sky130_fd_sc_hd__a21boi_1 _22594_ (.A1(_01539_),
    .A2(_01557_),
    .B1_N(_01560_),
    .Y(_01575_));
 sky130_fd_sc_hd__o32a_1 _22595_ (.A1(_09386_),
    .A2(_10752_),
    .A3(_00933_),
    .B1(_01050_),
    .B2(_01556_),
    .X(_01576_));
 sky130_fd_sc_hd__a21o_1 _22596_ (.A1(_01384_),
    .A2(_01552_),
    .B1(_01423_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _22597_ (.A0(_01543_),
    .A1(_01542_),
    .S(_01488_),
    .X(_01578_));
 sky130_fd_sc_hd__a21oi_1 _22598_ (.A1(_01549_),
    .A2(_01550_),
    .B1(_01578_),
    .Y(_01580_));
 sky130_fd_sc_hd__a21oi_1 _22599_ (.A1(_01489_),
    .A2(_01543_),
    .B1(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__xnor2_1 _22600_ (.A(_01577_),
    .B(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__xor2_1 _22601_ (.A(_01053_),
    .B(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__xor2_1 _22602_ (.A(_01576_),
    .B(_01583_),
    .X(_01584_));
 sky130_fd_sc_hd__a21o_1 _22603_ (.A1(_01053_),
    .A2(_01553_),
    .B1(_01555_),
    .X(_01585_));
 sky130_fd_sc_hd__xnor2_1 _22604_ (.A(_01584_),
    .B(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hd__xnor2_1 _22605_ (.A(_01575_),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__xnor2_1 _22606_ (.A(_01574_),
    .B(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__o211ai_1 _22607_ (.A1(_01565_),
    .A2(_01566_),
    .B1(_01588_),
    .C1(_01572_),
    .Y(_01589_));
 sky130_fd_sc_hd__o21bai_1 _22608_ (.A1(_01567_),
    .A2(_01571_),
    .B1_N(_01588_),
    .Y(_01591_));
 sky130_fd_sc_hd__nand2_1 _22609_ (.A(_01589_),
    .B(_01591_),
    .Y(net124));
 sky130_fd_sc_hd__and3_1 _22610_ (.A(_05152_),
    .B(_06171_),
    .C(_06182_),
    .X(_01592_));
 sky130_fd_sc_hd__nor2_1 _22611_ (.A(_06225_),
    .B(_01592_),
    .Y(net128));
 sky130_fd_sc_hd__o22a_1 _22612_ (.A1(_01737_),
    .A2(_01824_),
    .B1(_01846_),
    .B2(_01759_),
    .X(_01593_));
 sky130_fd_sc_hd__a31oi_2 _22613_ (.A1(net44),
    .A2(net12),
    .A3(net65),
    .B1(_01593_),
    .Y(net76));
 sky130_fd_sc_hd__xor2_1 _22614_ (.A(_02272_),
    .B(_02327_),
    .X(net87));
 sky130_fd_sc_hd__a2bb2o_1 _22615_ (.A1_N(_02272_),
    .A2_N(_02327_),
    .B1(_02436_),
    .B2(_02447_),
    .X(_01594_));
 sky130_fd_sc_hd__and2_1 _22616_ (.A(_02458_),
    .B(_01594_),
    .X(net98));
 sky130_fd_sc_hd__xor2_1 _22617_ (.A(_02458_),
    .B(_02688_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_16 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_16 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_16 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_16 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_16 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_16 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_16 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_16 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_16 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_16 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_16 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_16 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_16 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_16 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_16 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_16 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_16 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_16 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_16 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_16 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_16 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_16 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_16 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_16 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_16 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_16 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_16 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_16 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_16 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_16 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_16 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_16 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_16 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_16 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_16 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_16 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_16 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_16 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_16 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_16 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_16 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_16 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_16 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_16 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_16 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_16 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_16 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_16 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_16 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_16 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_12 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_12 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_16 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_16 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_16 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_16 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_16 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_16 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_16 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(P[0]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(P[10]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(P[11]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(P[12]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(P[13]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(P[14]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(P[15]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(P[16]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(P[17]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(P[18]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(P[19]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(P[1]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(P[20]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(P[21]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(P[22]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(P[23]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(P[24]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(P[25]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(P[26]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(P[27]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(P[28]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(P[29]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(P[2]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(P[30]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(P[31]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(P[32]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(P[33]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(P[34]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(P[35]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(P[36]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(P[37]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(P[38]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(P[39]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(P[3]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(P[40]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(P[41]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(P[42]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(P[43]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(P[44]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(P[45]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(P[46]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(P[47]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(P[48]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(P[49]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(P[4]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(P[50]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(P[51]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(P[52]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(P[53]));
 sky130_fd_sc_hd__buf_1 output114 (.A(net114),
    .X(P[54]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(P[55]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(P[56]));
 sky130_fd_sc_hd__buf_1 output117 (.A(net117),
    .X(P[57]));
 sky130_fd_sc_hd__buf_1 output118 (.A(net118),
    .X(P[58]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(P[59]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(P[5]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(P[60]));
 sky130_fd_sc_hd__buf_1 output122 (.A(net122),
    .X(P[61]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(P[62]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(P[63]));
 sky130_fd_sc_hd__buf_1 output125 (.A(net125),
    .X(P[6]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(P[7]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(P[8]));
 sky130_fd_sc_hd__buf_1 output128 (.A(net128),
    .X(P[9]));
endmodule
