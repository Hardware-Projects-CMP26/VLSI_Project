module carry_bypass_adder (Cin,
    Cout,
    Overflow,
    A,
    B,
    SUM);
 input Cin;
 output Cout;
 output Overflow;
 input [31:0] A;
 input [31:0] B;
 output [31:0] SUM;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire \ripple_loop[0].R.fa0.SUM ;
 wire \ripple_loop[0].R.fa31.SUM ;
 wire \ripple_loop[0].R.fa[1].SUM ;
 wire \ripple_loop[0].R.fa[2].SUM ;
 wire \ripple_loop[1].R.fa0.SUM ;
 wire \ripple_loop[1].R.fa31.SUM ;
 wire \ripple_loop[1].R.fa[1].SUM ;
 wire \ripple_loop[1].R.fa[2].SUM ;
 wire \ripple_loop[2].R.fa0.SUM ;
 wire \ripple_loop[2].R.fa31.SUM ;
 wire \ripple_loop[2].R.fa[1].SUM ;
 wire \ripple_loop[2].R.fa[2].SUM ;
 wire \ripple_loop[3].R.fa0.SUM ;
 wire \ripple_loop[3].R.fa31.SUM ;
 wire \ripple_loop[3].R.fa[1].SUM ;
 wire \ripple_loop[3].R.fa[2].SUM ;
 wire \ripple_loop[4].R.fa0.SUM ;
 wire \ripple_loop[4].R.fa31.SUM ;
 wire \ripple_loop[4].R.fa[1].SUM ;
 wire \ripple_loop[4].R.fa[2].SUM ;
 wire \ripple_loop[5].R.fa0.SUM ;
 wire \ripple_loop[5].R.fa31.SUM ;
 wire \ripple_loop[5].R.fa[1].SUM ;
 wire \ripple_loop[5].R.fa[2].SUM ;
 wire \ripple_loop[6].R.fa0.SUM ;
 wire \ripple_loop[6].R.fa31.SUM ;
 wire \ripple_loop[6].R.fa[1].SUM ;
 wire \ripple_loop[6].R.fa[2].SUM ;
 wire \ripple_loop[7].R.fa0.SUM ;
 wire \ripple_loop[7].R.fa31.SUM ;
 wire \ripple_loop[7].R.fa[1].SUM ;
 wire \ripple_loop[7].R.fa[2].SUM ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__nor2_1 _143_ (.A(net57),
    .B(net25),
    .Y(_000_));
 sky130_fd_sc_hd__or2_1 _144_ (.A(net57),
    .B(net25),
    .X(_001_));
 sky130_fd_sc_hd__and2_1 _145_ (.A(net57),
    .B(net25),
    .X(_002_));
 sky130_fd_sc_hd__nor2_1 _146_ (.A(_000_),
    .B(_002_),
    .Y(_003_));
 sky130_fd_sc_hd__and2_1 _147_ (.A(net56),
    .B(net24),
    .X(_004_));
 sky130_fd_sc_hd__nor2_1 _148_ (.A(net56),
    .B(net24),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_1 _149_ (.A(_004_),
    .B(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__or2_1 _150_ (.A(_004_),
    .B(_005_),
    .X(_007_));
 sky130_fd_sc_hd__nand2_1 _151_ (.A(net54),
    .B(net22),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_1 _152_ (.A(net53),
    .B(net21),
    .Y(_009_));
 sky130_fd_sc_hd__or2_1 _153_ (.A(net53),
    .B(net21),
    .X(_010_));
 sky130_fd_sc_hd__and2_1 _154_ (.A(_009_),
    .B(_010_),
    .X(_011_));
 sky130_fd_sc_hd__and2_1 _155_ (.A(net52),
    .B(net20),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _156_ (.A(net51),
    .B(net19),
    .X(_013_));
 sky130_fd_sc_hd__nor2_1 _157_ (.A(net51),
    .B(net19),
    .Y(_014_));
 sky130_fd_sc_hd__nor2_1 _158_ (.A(_013_),
    .B(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__and2_1 _159_ (.A(net50),
    .B(net18),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _160_ (.A(net49),
    .B(net17),
    .X(_017_));
 sky130_fd_sc_hd__nor2_1 _161_ (.A(net49),
    .B(net17),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _162_ (.A(_017_),
    .B(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__and2_1 _163_ (.A(net48),
    .B(net16),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _164_ (.A(net47),
    .B(net15),
    .X(_021_));
 sky130_fd_sc_hd__nor2_1 _165_ (.A(net47),
    .B(net15),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_1 _166_ (.A(_021_),
    .B(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__and2_1 _167_ (.A(net46),
    .B(net14),
    .X(_024_));
 sky130_fd_sc_hd__and2_1 _168_ (.A(net45),
    .B(net13),
    .X(_025_));
 sky130_fd_sc_hd__nor2_1 _169_ (.A(net45),
    .B(net13),
    .Y(_026_));
 sky130_fd_sc_hd__nor2_1 _170_ (.A(_025_),
    .B(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__and2_1 _171_ (.A(net43),
    .B(net11),
    .X(_028_));
 sky130_fd_sc_hd__and2_1 _172_ (.A(net42),
    .B(net10),
    .X(_029_));
 sky130_fd_sc_hd__nor2_1 _173_ (.A(net42),
    .B(net10),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_1 _174_ (.A(_029_),
    .B(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__and2_1 _175_ (.A(net41),
    .B(net9),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _176_ (.A(net40),
    .B(net8),
    .X(_033_));
 sky130_fd_sc_hd__nor2_1 _177_ (.A(net40),
    .B(net8),
    .Y(_034_));
 sky130_fd_sc_hd__nor2_1 _178_ (.A(_033_),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__and2_1 _179_ (.A(net39),
    .B(net7),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _180_ (.A(net38),
    .B(net6),
    .X(_037_));
 sky130_fd_sc_hd__nor2_1 _181_ (.A(net38),
    .B(net6),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _182_ (.A(_037_),
    .B(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__and2_1 _183_ (.A(net37),
    .B(net5),
    .X(_040_));
 sky130_fd_sc_hd__and2_1 _184_ (.A(net36),
    .B(net4),
    .X(_041_));
 sky130_fd_sc_hd__nor2_1 _185_ (.A(net36),
    .B(net4),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_1 _186_ (.A(_041_),
    .B(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__and2_1 _187_ (.A(net35),
    .B(net3),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _188_ (.A(net34),
    .B(net2),
    .X(_045_));
 sky130_fd_sc_hd__nor2_1 _189_ (.A(net34),
    .B(net2),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _190_ (.A(_045_),
    .B(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__and2_1 _191_ (.A(net64),
    .B(net32),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _192_ (.A(net63),
    .B(net31),
    .X(_049_));
 sky130_fd_sc_hd__nor2_1 _193_ (.A(net63),
    .B(net31),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _194_ (.A(_049_),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__and2_1 _195_ (.A(net62),
    .B(net30),
    .X(_052_));
 sky130_fd_sc_hd__and2_1 _196_ (.A(net61),
    .B(net29),
    .X(_053_));
 sky130_fd_sc_hd__nor2_1 _197_ (.A(net61),
    .B(net29),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _198_ (.A(_053_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__and2_1 _199_ (.A(net60),
    .B(net28),
    .X(_056_));
 sky130_fd_sc_hd__and2_1 _200_ (.A(net59),
    .B(net27),
    .X(_057_));
 sky130_fd_sc_hd__nor2_1 _201_ (.A(net59),
    .B(net27),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _202_ (.A(_057_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__and2_1 _203_ (.A(net58),
    .B(net26),
    .X(_060_));
 sky130_fd_sc_hd__and2_1 _204_ (.A(net55),
    .B(net23),
    .X(_061_));
 sky130_fd_sc_hd__nand2_1 _205_ (.A(net55),
    .B(net23),
    .Y(_062_));
 sky130_fd_sc_hd__or2_1 _206_ (.A(net55),
    .B(net23),
    .X(_063_));
 sky130_fd_sc_hd__or2_1 _207_ (.A(net44),
    .B(net12),
    .X(_064_));
 sky130_fd_sc_hd__nand2_1 _208_ (.A(net44),
    .B(net12),
    .Y(_065_));
 sky130_fd_sc_hd__or2_1 _209_ (.A(net33),
    .B(net1),
    .X(_066_));
 sky130_fd_sc_hd__nand2_1 _210_ (.A(net33),
    .B(net1),
    .Y(_067_));
 sky130_fd_sc_hd__o21ai_1 _211_ (.A1(net33),
    .A2(net1),
    .B1(net65),
    .Y(_068_));
 sky130_fd_sc_hd__and2_1 _212_ (.A(_067_),
    .B(_068_),
    .X(_069_));
 sky130_fd_sc_hd__nand3_1 _213_ (.A(_065_),
    .B(_067_),
    .C(_068_),
    .Y(_070_));
 sky130_fd_sc_hd__o2111ai_1 _214_ (.A1(net44),
    .A2(net12),
    .B1(_062_),
    .C1(_063_),
    .D1(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__a31oi_2 _215_ (.A1(_063_),
    .A2(_064_),
    .A3(_070_),
    .B1(_061_),
    .Y(_072_));
 sky130_fd_sc_hd__nor2_1 _216_ (.A(net58),
    .B(net26),
    .Y(_073_));
 sky130_fd_sc_hd__or2_1 _217_ (.A(_060_),
    .B(_073_),
    .X(_074_));
 sky130_fd_sc_hd__o21bai_1 _218_ (.A1(_074_),
    .A2(_072_),
    .B1_N(_060_),
    .Y(_075_));
 sky130_fd_sc_hd__a21oi_1 _219_ (.A1(_075_),
    .A2(_059_),
    .B1(_057_),
    .Y(_076_));
 sky130_fd_sc_hd__nor2_1 _220_ (.A(net60),
    .B(net28),
    .Y(_077_));
 sky130_fd_sc_hd__or2_1 _221_ (.A(_056_),
    .B(_077_),
    .X(_078_));
 sky130_fd_sc_hd__o21bai_1 _222_ (.A1(_078_),
    .A2(_076_),
    .B1_N(_056_),
    .Y(_079_));
 sky130_fd_sc_hd__a21oi_1 _223_ (.A1(_079_),
    .A2(_055_),
    .B1(_053_),
    .Y(_080_));
 sky130_fd_sc_hd__nor2_1 _224_ (.A(net62),
    .B(net30),
    .Y(_081_));
 sky130_fd_sc_hd__or2_1 _225_ (.A(_052_),
    .B(_081_),
    .X(_082_));
 sky130_fd_sc_hd__o21bai_1 _226_ (.A1(_082_),
    .A2(_080_),
    .B1_N(_052_),
    .Y(_083_));
 sky130_fd_sc_hd__a21oi_1 _227_ (.A1(_083_),
    .A2(_051_),
    .B1(_049_),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_1 _228_ (.A(net64),
    .B(net32),
    .Y(_085_));
 sky130_fd_sc_hd__or2_1 _229_ (.A(_048_),
    .B(_085_),
    .X(_086_));
 sky130_fd_sc_hd__o21bai_1 _230_ (.A1(_086_),
    .A2(_084_),
    .B1_N(_048_),
    .Y(_087_));
 sky130_fd_sc_hd__a21oi_1 _231_ (.A1(_087_),
    .A2(_047_),
    .B1(_045_),
    .Y(_088_));
 sky130_fd_sc_hd__nor2_1 _232_ (.A(net35),
    .B(net3),
    .Y(_089_));
 sky130_fd_sc_hd__or2_1 _233_ (.A(_044_),
    .B(_089_),
    .X(_090_));
 sky130_fd_sc_hd__o21bai_1 _234_ (.A1(_090_),
    .A2(_088_),
    .B1_N(_044_),
    .Y(_091_));
 sky130_fd_sc_hd__a21oi_1 _235_ (.A1(_091_),
    .A2(_043_),
    .B1(_041_),
    .Y(_092_));
 sky130_fd_sc_hd__nor2_1 _236_ (.A(net37),
    .B(net5),
    .Y(_093_));
 sky130_fd_sc_hd__or2_1 _237_ (.A(_040_),
    .B(_093_),
    .X(_094_));
 sky130_fd_sc_hd__o21bai_1 _238_ (.A1(_094_),
    .A2(_092_),
    .B1_N(_040_),
    .Y(_095_));
 sky130_fd_sc_hd__a21oi_1 _239_ (.A1(_095_),
    .A2(_039_),
    .B1(_037_),
    .Y(_096_));
 sky130_fd_sc_hd__nor2_1 _240_ (.A(net39),
    .B(net7),
    .Y(_097_));
 sky130_fd_sc_hd__or2_1 _241_ (.A(_036_),
    .B(_097_),
    .X(_098_));
 sky130_fd_sc_hd__o21bai_1 _242_ (.A1(_098_),
    .A2(_096_),
    .B1_N(_036_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _243_ (.A1(_099_),
    .A2(_035_),
    .B1(_033_),
    .Y(_100_));
 sky130_fd_sc_hd__nor2_1 _244_ (.A(net41),
    .B(net9),
    .Y(_101_));
 sky130_fd_sc_hd__or2_1 _245_ (.A(_032_),
    .B(_101_),
    .X(_102_));
 sky130_fd_sc_hd__o21bai_1 _246_ (.A1(_102_),
    .A2(_100_),
    .B1_N(_032_),
    .Y(_103_));
 sky130_fd_sc_hd__a21oi_1 _247_ (.A1(_103_),
    .A2(_031_),
    .B1(_029_),
    .Y(_104_));
 sky130_fd_sc_hd__nor2_1 _248_ (.A(net43),
    .B(net11),
    .Y(_105_));
 sky130_fd_sc_hd__or2_1 _249_ (.A(_028_),
    .B(_105_),
    .X(_106_));
 sky130_fd_sc_hd__o21bai_1 _250_ (.A1(_106_),
    .A2(_104_),
    .B1_N(_028_),
    .Y(_107_));
 sky130_fd_sc_hd__a21oi_1 _251_ (.A1(_107_),
    .A2(_027_),
    .B1(_025_),
    .Y(_108_));
 sky130_fd_sc_hd__nor2_1 _252_ (.A(net46),
    .B(net14),
    .Y(_109_));
 sky130_fd_sc_hd__or2_1 _253_ (.A(_024_),
    .B(_109_),
    .X(_110_));
 sky130_fd_sc_hd__o21bai_1 _254_ (.A1(_110_),
    .A2(_108_),
    .B1_N(_024_),
    .Y(_111_));
 sky130_fd_sc_hd__a21oi_1 _255_ (.A1(_111_),
    .A2(_023_),
    .B1(_021_),
    .Y(_112_));
 sky130_fd_sc_hd__nor2_1 _256_ (.A(net48),
    .B(net16),
    .Y(_113_));
 sky130_fd_sc_hd__or2_1 _257_ (.A(_020_),
    .B(_113_),
    .X(_114_));
 sky130_fd_sc_hd__o21bai_1 _258_ (.A1(_114_),
    .A2(_112_),
    .B1_N(_020_),
    .Y(_115_));
 sky130_fd_sc_hd__a21oi_1 _259_ (.A1(_115_),
    .A2(_019_),
    .B1(_017_),
    .Y(_116_));
 sky130_fd_sc_hd__nor2_1 _260_ (.A(net50),
    .B(net18),
    .Y(_117_));
 sky130_fd_sc_hd__or2_1 _261_ (.A(_016_),
    .B(_117_),
    .X(_118_));
 sky130_fd_sc_hd__o21bai_1 _262_ (.A1(_118_),
    .A2(_116_),
    .B1_N(_016_),
    .Y(_119_));
 sky130_fd_sc_hd__a21oi_1 _263_ (.A1(_119_),
    .A2(_015_),
    .B1(_013_),
    .Y(_120_));
 sky130_fd_sc_hd__nor2_1 _264_ (.A(net52),
    .B(net20),
    .Y(_121_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(_012_),
    .B(_121_),
    .X(_122_));
 sky130_fd_sc_hd__o21bai_2 _266_ (.A1(_122_),
    .A2(_120_),
    .B1_N(_012_),
    .Y(_123_));
 sky130_fd_sc_hd__nand2_1 _267_ (.A(_123_),
    .B(_011_),
    .Y(_124_));
 sky130_fd_sc_hd__a21boi_1 _268_ (.A1(_123_),
    .A2(_011_),
    .B1_N(_009_),
    .Y(_125_));
 sky130_fd_sc_hd__and2b_1 _269_ (.A_N(net54),
    .B(net22),
    .X(_126_));
 sky130_fd_sc_hd__and2b_1 _270_ (.A_N(net22),
    .B(net54),
    .X(_127_));
 sky130_fd_sc_hd__nor2_1 _271_ (.A(_126_),
    .B(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__o2bb2ai_1 _272_ (.A1_N(_009_),
    .A2_N(_124_),
    .B1(_126_),
    .B2(_127_),
    .Y(_129_));
 sky130_fd_sc_hd__o21ai_1 _273_ (.A1(_128_),
    .A2(_125_),
    .B1(_008_),
    .Y(_130_));
 sky130_fd_sc_hd__a21oi_2 _274_ (.A1(_008_),
    .A2(_129_),
    .B1(_007_),
    .Y(_131_));
 sky130_fd_sc_hd__nand2_1 _275_ (.A(_130_),
    .B(_006_),
    .Y(_132_));
 sky130_fd_sc_hd__a21oi_1 _276_ (.A1(_130_),
    .A2(_006_),
    .B1(_004_),
    .Y(_133_));
 sky130_fd_sc_hd__o22ai_1 _277_ (.A1(_000_),
    .A2(_002_),
    .B1(_004_),
    .B2(_131_),
    .Y(_134_));
 sky130_fd_sc_hd__nand3b_1 _278_ (.A_N(_004_),
    .B(_132_),
    .C(_003_),
    .Y(_135_));
 sky130_fd_sc_hd__nand2_1 _279_ (.A(_134_),
    .B(_135_),
    .Y(\ripple_loop[7].R.fa31.SUM ));
 sky130_fd_sc_hd__a22o_1 _280_ (.A1(net57),
    .A2(net25),
    .B1(net56),
    .B2(net24),
    .X(_136_));
 sky130_fd_sc_hd__o22a_1 _281_ (.A1(_136_),
    .A2(_131_),
    .B1(_000_),
    .B2(_133_),
    .X(net67));
 sky130_fd_sc_hd__a22o_1 _282_ (.A1(_062_),
    .A2(_063_),
    .B1(_064_),
    .B2(_070_),
    .X(_137_));
 sky130_fd_sc_hd__and2_1 _283_ (.A(_071_),
    .B(_137_),
    .X(\ripple_loop[0].R.fa[2].SUM ));
 sky130_fd_sc_hd__and3_1 _284_ (.A(_064_),
    .B(_065_),
    .C(_069_),
    .X(_138_));
 sky130_fd_sc_hd__a21oi_1 _285_ (.A1(_064_),
    .A2(_065_),
    .B1(_069_),
    .Y(_139_));
 sky130_fd_sc_hd__or2_1 _286_ (.A(_138_),
    .B(_139_),
    .X(\ripple_loop[0].R.fa[1].SUM ));
 sky130_fd_sc_hd__xor2_1 _287_ (.A(_072_),
    .B(_074_),
    .X(\ripple_loop[0].R.fa31.SUM ));
 sky130_fd_sc_hd__and3_1 _288_ (.A(net65),
    .B(net33),
    .C(net1),
    .X(_140_));
 sky130_fd_sc_hd__o22a_1 _289_ (.A1(net65),
    .A2(_066_),
    .B1(_140_),
    .B2(_069_),
    .X(\ripple_loop[0].R.fa0.SUM ));
 sky130_fd_sc_hd__xor2_1 _290_ (.A(_055_),
    .B(_079_),
    .X(\ripple_loop[1].R.fa[2].SUM ));
 sky130_fd_sc_hd__xor2_1 _291_ (.A(_076_),
    .B(_078_),
    .X(\ripple_loop[1].R.fa[1].SUM ));
 sky130_fd_sc_hd__xor2_1 _292_ (.A(_080_),
    .B(_082_),
    .X(\ripple_loop[1].R.fa31.SUM ));
 sky130_fd_sc_hd__xor2_1 _293_ (.A(_059_),
    .B(_075_),
    .X(\ripple_loop[1].R.fa0.SUM ));
 sky130_fd_sc_hd__xor2_1 _294_ (.A(_047_),
    .B(_087_),
    .X(\ripple_loop[2].R.fa[2].SUM ));
 sky130_fd_sc_hd__xor2_1 _295_ (.A(_084_),
    .B(_086_),
    .X(\ripple_loop[2].R.fa[1].SUM ));
 sky130_fd_sc_hd__xor2_1 _296_ (.A(_088_),
    .B(_090_),
    .X(\ripple_loop[2].R.fa31.SUM ));
 sky130_fd_sc_hd__xor2_1 _297_ (.A(_051_),
    .B(_083_),
    .X(\ripple_loop[2].R.fa0.SUM ));
 sky130_fd_sc_hd__xor2_1 _298_ (.A(_039_),
    .B(_095_),
    .X(\ripple_loop[3].R.fa[2].SUM ));
 sky130_fd_sc_hd__xor2_1 _299_ (.A(_092_),
    .B(_094_),
    .X(\ripple_loop[3].R.fa[1].SUM ));
 sky130_fd_sc_hd__xor2_1 _300_ (.A(_096_),
    .B(_098_),
    .X(\ripple_loop[3].R.fa31.SUM ));
 sky130_fd_sc_hd__xor2_1 _301_ (.A(_043_),
    .B(_091_),
    .X(\ripple_loop[3].R.fa0.SUM ));
 sky130_fd_sc_hd__xor2_1 _302_ (.A(_031_),
    .B(_103_),
    .X(\ripple_loop[4].R.fa[2].SUM ));
 sky130_fd_sc_hd__xor2_1 _303_ (.A(_100_),
    .B(_102_),
    .X(\ripple_loop[4].R.fa[1].SUM ));
 sky130_fd_sc_hd__xor2_1 _304_ (.A(_104_),
    .B(_106_),
    .X(\ripple_loop[4].R.fa31.SUM ));
 sky130_fd_sc_hd__xor2_1 _305_ (.A(_035_),
    .B(_099_),
    .X(\ripple_loop[4].R.fa0.SUM ));
 sky130_fd_sc_hd__xor2_1 _306_ (.A(_023_),
    .B(_111_),
    .X(\ripple_loop[5].R.fa[2].SUM ));
 sky130_fd_sc_hd__xor2_1 _307_ (.A(_108_),
    .B(_110_),
    .X(\ripple_loop[5].R.fa[1].SUM ));
 sky130_fd_sc_hd__xor2_1 _308_ (.A(_112_),
    .B(_114_),
    .X(\ripple_loop[5].R.fa31.SUM ));
 sky130_fd_sc_hd__xor2_1 _309_ (.A(_027_),
    .B(_107_),
    .X(\ripple_loop[5].R.fa0.SUM ));
 sky130_fd_sc_hd__xor2_1 _310_ (.A(_015_),
    .B(_119_),
    .X(\ripple_loop[6].R.fa[2].SUM ));
 sky130_fd_sc_hd__xor2_1 _311_ (.A(_116_),
    .B(_118_),
    .X(\ripple_loop[6].R.fa[1].SUM ));
 sky130_fd_sc_hd__xor2_1 _312_ (.A(_120_),
    .B(_122_),
    .X(\ripple_loop[6].R.fa31.SUM ));
 sky130_fd_sc_hd__xor2_1 _313_ (.A(_019_),
    .B(_115_),
    .X(\ripple_loop[6].R.fa0.SUM ));
 sky130_fd_sc_hd__o221a_1 _314_ (.A1(_004_),
    .A2(_005_),
    .B1(_128_),
    .B2(_125_),
    .C1(_008_),
    .X(_141_));
 sky130_fd_sc_hd__nor2_1 _315_ (.A(_131_),
    .B(_141_),
    .Y(\ripple_loop[7].R.fa[2].SUM ));
 sky130_fd_sc_hd__nand2_1 _316_ (.A(_125_),
    .B(_128_),
    .Y(_142_));
 sky130_fd_sc_hd__and2_1 _317_ (.A(_129_),
    .B(_142_),
    .X(\ripple_loop[7].R.fa[1].SUM ));
 sky130_fd_sc_hd__o31a_1 _318_ (.A1(_002_),
    .A2(_004_),
    .A3(_131_),
    .B1(_001_),
    .X(net66));
 sky130_fd_sc_hd__xor2_1 _319_ (.A(_011_),
    .B(_123_),
    .X(\ripple_loop[7].R.fa0.SUM ));
 sky130_fd_sc_hd__clkbuf_1 _320_ (.A(\ripple_loop[0].R.fa0.SUM ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _321_ (.A(\ripple_loop[0].R.fa[1].SUM ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _322_ (.A(\ripple_loop[0].R.fa[2].SUM ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _323_ (.A(\ripple_loop[0].R.fa31.SUM ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _324_ (.A(\ripple_loop[1].R.fa0.SUM ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _325_ (.A(\ripple_loop[1].R.fa[1].SUM ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _326_ (.A(\ripple_loop[1].R.fa[2].SUM ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _327_ (.A(\ripple_loop[1].R.fa31.SUM ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _328_ (.A(\ripple_loop[2].R.fa0.SUM ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _329_ (.A(\ripple_loop[2].R.fa[1].SUM ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _330_ (.A(\ripple_loop[2].R.fa[2].SUM ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _331_ (.A(\ripple_loop[2].R.fa31.SUM ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _332_ (.A(\ripple_loop[3].R.fa0.SUM ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _333_ (.A(\ripple_loop[3].R.fa[1].SUM ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _334_ (.A(\ripple_loop[3].R.fa[2].SUM ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _335_ (.A(\ripple_loop[3].R.fa31.SUM ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _336_ (.A(\ripple_loop[4].R.fa0.SUM ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _337_ (.A(\ripple_loop[4].R.fa[1].SUM ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _338_ (.A(\ripple_loop[4].R.fa[2].SUM ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _339_ (.A(\ripple_loop[4].R.fa31.SUM ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _340_ (.A(\ripple_loop[5].R.fa0.SUM ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _341_ (.A(\ripple_loop[5].R.fa[1].SUM ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _342_ (.A(\ripple_loop[5].R.fa[2].SUM ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _343_ (.A(\ripple_loop[5].R.fa31.SUM ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _344_ (.A(\ripple_loop[6].R.fa0.SUM ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _345_ (.A(\ripple_loop[6].R.fa[1].SUM ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _346_ (.A(\ripple_loop[6].R.fa[2].SUM ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _347_ (.A(\ripple_loop[6].R.fa31.SUM ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _348_ (.A(\ripple_loop[7].R.fa0.SUM ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _349_ (.A(\ripple_loop[7].R.fa[1].SUM ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _350_ (.A(\ripple_loop[7].R.fa[2].SUM ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _351_ (.A(\ripple_loop[7].R.fa31.SUM ),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(Cin),
    .X(net65));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(Cout));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(Overflow));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(SUM[0]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(SUM[10]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(SUM[11]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(SUM[12]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(SUM[13]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(SUM[14]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(SUM[15]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(SUM[16]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(SUM[17]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(SUM[18]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(SUM[19]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(SUM[1]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(SUM[20]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(SUM[21]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(SUM[22]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(SUM[23]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(SUM[24]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(SUM[25]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(SUM[26]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(SUM[27]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(SUM[28]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(SUM[29]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(SUM[2]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(SUM[30]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(SUM[31]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(SUM[3]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(SUM[4]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(SUM[5]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(SUM[6]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(SUM[7]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(SUM[8]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(SUM[9]));
endmodule
