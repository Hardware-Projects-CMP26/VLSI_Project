module booth_multiplier (multiplicand,
    multiplier,
    product);
 input [31:0] multiplicand;
 input [31:0] multiplier;
 output [63:0] product;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;

 sky130_fd_sc_hd__clkinv_16 _13382_ (.A(net1),
    .Y(_03176_));
 sky130_fd_sc_hd__clkinv_16 _13383_ (.A(net33),
    .Y(_03286_));
 sky130_fd_sc_hd__clkinv_16 _13384_ (.A(net23),
    .Y(_03396_));
 sky130_fd_sc_hd__clkinv_16 _13385_ (.A(net26),
    .Y(_03506_));
 sky130_fd_sc_hd__inv_16 _13386_ (.A(net27),
    .Y(_03616_));
 sky130_fd_sc_hd__inv_12 _13387_ (.A(net28),
    .Y(_03725_));
 sky130_fd_sc_hd__inv_16 _13388_ (.A(net29),
    .Y(_03835_));
 sky130_fd_sc_hd__clkinv_16 _13389_ (.A(net30),
    .Y(_03916_));
 sky130_fd_sc_hd__clkinv_16 _13390_ (.A(net62),
    .Y(_03927_));
 sky130_fd_sc_hd__clkinv_16 _13391_ (.A(net31),
    .Y(_03938_));
 sky130_fd_sc_hd__inv_16 _13392_ (.A(net32),
    .Y(_03949_));
 sky130_fd_sc_hd__inv_16 _13393_ (.A(net2),
    .Y(_03960_));
 sky130_fd_sc_hd__inv_16 _13394_ (.A(net34),
    .Y(_03971_));
 sky130_fd_sc_hd__inv_16 _13395_ (.A(net3),
    .Y(_03982_));
 sky130_fd_sc_hd__inv_16 _13396_ (.A(net35),
    .Y(_03993_));
 sky130_fd_sc_hd__inv_16 _13397_ (.A(net4),
    .Y(_04004_));
 sky130_fd_sc_hd__inv_16 _13398_ (.A(net5),
    .Y(_04015_));
 sky130_fd_sc_hd__inv_16 _13399_ (.A(net6),
    .Y(_04026_));
 sky130_fd_sc_hd__inv_16 _13400_ (.A(net38),
    .Y(_04037_));
 sky130_fd_sc_hd__inv_16 _13401_ (.A(net7),
    .Y(_04048_));
 sky130_fd_sc_hd__inv_16 _13402_ (.A(net8),
    .Y(_04059_));
 sky130_fd_sc_hd__inv_16 _13403_ (.A(net9),
    .Y(_04069_));
 sky130_fd_sc_hd__inv_16 _13404_ (.A(net10),
    .Y(_04080_));
 sky130_fd_sc_hd__inv_16 _13405_ (.A(net11),
    .Y(_04091_));
 sky130_fd_sc_hd__inv_16 _13406_ (.A(net43),
    .Y(_04102_));
 sky130_fd_sc_hd__inv_16 _13407_ (.A(net13),
    .Y(_04113_));
 sky130_fd_sc_hd__inv_16 _13408_ (.A(net45),
    .Y(_04124_));
 sky130_fd_sc_hd__inv_16 _13409_ (.A(net14),
    .Y(_04135_));
 sky130_fd_sc_hd__inv_16 _13410_ (.A(net15),
    .Y(_04146_));
 sky130_fd_sc_hd__clkinv_16 _13411_ (.A(net16),
    .Y(_04157_));
 sky130_fd_sc_hd__inv_8 _13412_ (.A(net17),
    .Y(_04168_));
 sky130_fd_sc_hd__inv_16 _13413_ (.A(net18),
    .Y(_04179_));
 sky130_fd_sc_hd__inv_16 _13414_ (.A(net50),
    .Y(_04190_));
 sky130_fd_sc_hd__inv_16 _13415_ (.A(net19),
    .Y(_04201_));
 sky130_fd_sc_hd__inv_16 _13416_ (.A(net20),
    .Y(_04212_));
 sky130_fd_sc_hd__inv_16 _13417_ (.A(net21),
    .Y(_04223_));
 sky130_fd_sc_hd__inv_4 _13418_ (.A(net53),
    .Y(_04234_));
 sky130_fd_sc_hd__clkinv_16 _13419_ (.A(net22),
    .Y(_04245_));
 sky130_fd_sc_hd__inv_16 _13420_ (.A(net24),
    .Y(_04256_));
 sky130_fd_sc_hd__inv_16 _13421_ (.A(net56),
    .Y(_04266_));
 sky130_fd_sc_hd__clkinv_16 _13422_ (.A(net25),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_1 _13423_ (.A(_03176_),
    .B(_03286_),
    .Y(net65));
 sky130_fd_sc_hd__and2b_2 _13424_ (.A_N(net12),
    .B(net1),
    .X(_04298_));
 sky130_fd_sc_hd__nand2b_2 _13425_ (.A_N(net12),
    .B(net1),
    .Y(_04309_));
 sky130_fd_sc_hd__nor2_8 _13426_ (.A(net44),
    .B(_03286_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand2b_4 _13427_ (.A_N(net44),
    .B(net33),
    .Y(_04331_));
 sky130_fd_sc_hd__and2b_4 _13428_ (.A_N(net44),
    .B(net55),
    .X(_04342_));
 sky130_fd_sc_hd__nand2b_4 _13429_ (.A_N(net44),
    .B(net55),
    .Y(_04353_));
 sky130_fd_sc_hd__and2b_4 _13430_ (.A_N(net55),
    .B(net44),
    .X(_04364_));
 sky130_fd_sc_hd__nand2b_4 _13431_ (.A_N(net55),
    .B(net44),
    .Y(_04375_));
 sky130_fd_sc_hd__a21oi_1 _13432_ (.A1(_04353_),
    .A2(_04375_),
    .B1(_03176_),
    .Y(_04386_));
 sky130_fd_sc_hd__nor2_8 _13433_ (.A(net1),
    .B(net12),
    .Y(_04397_));
 sky130_fd_sc_hd__o21a_4 _13434_ (.A1(net1),
    .A2(net12),
    .B1(net23),
    .X(_04408_));
 sky130_fd_sc_hd__o21ai_4 _13435_ (.A1(net1),
    .A2(net12),
    .B1(net23),
    .Y(_04419_));
 sky130_fd_sc_hd__nor2_4 _13436_ (.A(net12),
    .B(net23),
    .Y(_04430_));
 sky130_fd_sc_hd__nor3_4 _13437_ (.A(net1),
    .B(net12),
    .C(net23),
    .Y(_04441_));
 sky130_fd_sc_hd__nand2_8 _13438_ (.A(_04397_),
    .B(_03396_),
    .Y(_04452_));
 sky130_fd_sc_hd__a21oi_4 _13439_ (.A1(_03176_),
    .A2(_04430_),
    .B1(_04408_),
    .Y(_04463_));
 sky130_fd_sc_hd__a21o_4 _13440_ (.A1(_03176_),
    .A2(_04430_),
    .B1(_04408_),
    .X(_04474_));
 sky130_fd_sc_hd__and2b_4 _13441_ (.A_N(net33),
    .B(net44),
    .X(_04484_));
 sky130_fd_sc_hd__nand2_8 _13442_ (.A(_03286_),
    .B(net44),
    .Y(_04495_));
 sky130_fd_sc_hd__and2b_2 _13443_ (.A_N(net1),
    .B(net12),
    .X(_04506_));
 sky130_fd_sc_hd__nand2b_2 _13444_ (.A_N(net1),
    .B(net12),
    .Y(_04517_));
 sky130_fd_sc_hd__xnor2_4 _13445_ (.A(net1),
    .B(net12),
    .Y(_04528_));
 sky130_fd_sc_hd__nand2_8 _13446_ (.A(_04309_),
    .B(_04517_),
    .Y(_04539_));
 sky130_fd_sc_hd__a22o_1 _13447_ (.A1(net12),
    .A2(_04320_),
    .B1(_04539_),
    .B2(_04484_),
    .X(_04550_));
 sky130_fd_sc_hd__and3_1 _13448_ (.A(_04550_),
    .B(_04463_),
    .C(net33),
    .X(_04561_));
 sky130_fd_sc_hd__a31o_1 _13449_ (.A1(net33),
    .A2(_04419_),
    .A3(_04452_),
    .B1(_04550_),
    .X(_04572_));
 sky130_fd_sc_hd__and2b_1 _13450_ (.A_N(_04561_),
    .B(_04572_),
    .X(_04583_));
 sky130_fd_sc_hd__xor2_1 _13451_ (.A(_04386_),
    .B(_04583_),
    .X(_04594_));
 sky130_fd_sc_hd__and3_2 _13452_ (.A(_04298_),
    .B(_04320_),
    .C(_04594_),
    .X(_04605_));
 sky130_fd_sc_hd__or4b_1 _13453_ (.A(_03176_),
    .B(net12),
    .C(_04331_),
    .D_N(_04594_),
    .X(_04616_));
 sky130_fd_sc_hd__and2b_4 _13454_ (.A_N(net55),
    .B(net58),
    .X(_04627_));
 sky130_fd_sc_hd__nand2b_4 _13455_ (.A_N(net55),
    .B(net58),
    .Y(_04638_));
 sky130_fd_sc_hd__and2b_4 _13456_ (.A_N(net58),
    .B(net55),
    .X(_04649_));
 sky130_fd_sc_hd__nand2b_4 _13457_ (.A_N(net58),
    .B(net55),
    .Y(_04660_));
 sky130_fd_sc_hd__o21ai_1 _13458_ (.A1(_04627_),
    .A2(_04649_),
    .B1(net1),
    .Y(_04671_));
 sky130_fd_sc_hd__a21oi_1 _13459_ (.A1(_04572_),
    .A2(_04386_),
    .B1(_04561_),
    .Y(_04682_));
 sky130_fd_sc_hd__a22o_1 _13460_ (.A1(net12),
    .A2(_04364_),
    .B1(_04539_),
    .B2(_04342_),
    .X(_04693_));
 sky130_fd_sc_hd__o31a_4 _13461_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .B1(net26),
    .X(_04703_));
 sky130_fd_sc_hd__o31ai_2 _13462_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .B1(net26),
    .Y(_04714_));
 sky130_fd_sc_hd__nor2_8 _13463_ (.A(net23),
    .B(net26),
    .Y(_04725_));
 sky130_fd_sc_hd__nor4_4 _13464_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(net26),
    .Y(_04736_));
 sky130_fd_sc_hd__nand2_8 _13465_ (.A(_04397_),
    .B(_04725_),
    .Y(_04747_));
 sky130_fd_sc_hd__nand2_8 _13466_ (.A(net314),
    .B(net267),
    .Y(_04758_));
 sky130_fd_sc_hd__a211o_1 _13467_ (.A1(_03176_),
    .A2(_04430_),
    .B1(_04408_),
    .C1(_04495_),
    .X(_04769_));
 sky130_fd_sc_hd__o221ai_4 _13468_ (.A1(_03396_),
    .A2(_04331_),
    .B1(_04758_),
    .B2(_03286_),
    .C1(_04769_),
    .Y(_04780_));
 sky130_fd_sc_hd__o31a_1 _13469_ (.A1(_03396_),
    .A2(net26),
    .A3(_04331_),
    .B1(_04780_),
    .X(_04791_));
 sky130_fd_sc_hd__xnor2_1 _13470_ (.A(_04693_),
    .B(_04791_),
    .Y(_04802_));
 sky130_fd_sc_hd__or2_1 _13471_ (.A(_04682_),
    .B(_04802_),
    .X(_04813_));
 sky130_fd_sc_hd__nand2_1 _13472_ (.A(_04802_),
    .B(_04682_),
    .Y(_04824_));
 sky130_fd_sc_hd__o2111ai_2 _13473_ (.A1(_04627_),
    .A2(_04649_),
    .B1(_04824_),
    .C1(net1),
    .D1(_04813_),
    .Y(_04835_));
 sky130_fd_sc_hd__and3_1 _13474_ (.A(_04671_),
    .B(_04813_),
    .C(_04824_),
    .X(_04846_));
 sky130_fd_sc_hd__a21oi_2 _13475_ (.A1(_04813_),
    .A2(_04824_),
    .B1(_04671_),
    .Y(_04857_));
 sky130_fd_sc_hd__nor2_1 _13476_ (.A(_04846_),
    .B(_04857_),
    .Y(_04868_));
 sky130_fd_sc_hd__xnor2_1 _13477_ (.A(_04605_),
    .B(_04868_),
    .Y(net98));
 sky130_fd_sc_hd__and2b_4 _13478_ (.A_N(net58),
    .B(net59),
    .X(_04889_));
 sky130_fd_sc_hd__nand2b_4 _13479_ (.A_N(net58),
    .B(net59),
    .Y(_04900_));
 sky130_fd_sc_hd__and2b_4 _13480_ (.A_N(net59),
    .B(net58),
    .X(_04911_));
 sky130_fd_sc_hd__o21a_1 _13481_ (.A1(net305),
    .A2(_04911_),
    .B1(net1),
    .X(_04922_));
 sky130_fd_sc_hd__a22o_1 _13482_ (.A1(net12),
    .A2(_04649_),
    .B1(_04539_),
    .B2(_04627_),
    .X(_04933_));
 sky130_fd_sc_hd__nand2_2 _13483_ (.A(_04933_),
    .B(_04922_),
    .Y(_04943_));
 sky130_fd_sc_hd__a221o_1 _13484_ (.A1(_04539_),
    .A2(net317),
    .B1(_04649_),
    .B2(net12),
    .C1(_04922_),
    .X(_04954_));
 sky130_fd_sc_hd__nand2_1 _13485_ (.A(_04943_),
    .B(_04954_),
    .Y(_04965_));
 sky130_fd_sc_hd__a32oi_4 _13486_ (.A1(net23),
    .A2(_04320_),
    .A3(_03506_),
    .B1(_04780_),
    .B2(_04693_),
    .Y(_04976_));
 sky130_fd_sc_hd__a32o_1 _13487_ (.A1(_04452_),
    .A2(_04342_),
    .A3(_04419_),
    .B1(_04364_),
    .B2(net23),
    .X(_04987_));
 sky130_fd_sc_hd__nand4_4 _13488_ (.A(_04397_),
    .B(_03616_),
    .C(_03506_),
    .D(_03396_),
    .Y(_04998_));
 sky130_fd_sc_hd__o41ai_4 _13489_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .A4(net26),
    .B1(net27),
    .Y(_05009_));
 sky130_fd_sc_hd__nand2_8 _13490_ (.A(net266),
    .B(net302),
    .Y(_05020_));
 sky130_fd_sc_hd__nand3_1 _13491_ (.A(net300),
    .B(net33),
    .C(_04998_),
    .Y(_05031_));
 sky130_fd_sc_hd__and4b_1 _13492_ (.A_N(net44),
    .B(_03616_),
    .C(net33),
    .D(net26),
    .X(_05042_));
 sky130_fd_sc_hd__or4_1 _13493_ (.A(net44),
    .B(net27),
    .C(_03286_),
    .D(_03506_),
    .X(_05053_));
 sky130_fd_sc_hd__o221a_1 _13494_ (.A1(_03506_),
    .A2(_04331_),
    .B1(_04495_),
    .B2(_04758_),
    .C1(_05031_),
    .X(_05064_));
 sky130_fd_sc_hd__o221ai_2 _13495_ (.A1(_03506_),
    .A2(_04331_),
    .B1(_04495_),
    .B2(_04758_),
    .C1(_05031_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand3b_1 _13496_ (.A_N(_04987_),
    .B(_05053_),
    .C(_05075_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21ai_1 _13497_ (.A1(_05042_),
    .A2(_05064_),
    .B1(_04987_),
    .Y(_05097_));
 sky130_fd_sc_hd__a21oi_1 _13498_ (.A1(_05086_),
    .A2(_05097_),
    .B1(_04976_),
    .Y(_05108_));
 sky130_fd_sc_hd__a21o_1 _13499_ (.A1(_05086_),
    .A2(_05097_),
    .B1(_04976_),
    .X(_05119_));
 sky130_fd_sc_hd__nand3_1 _13500_ (.A(_04976_),
    .B(_05086_),
    .C(_05097_),
    .Y(_05130_));
 sky130_fd_sc_hd__nand2_1 _13501_ (.A(_05119_),
    .B(_05130_),
    .Y(_05141_));
 sky130_fd_sc_hd__xnor2_1 _13502_ (.A(_04965_),
    .B(_05141_),
    .Y(_05152_));
 sky130_fd_sc_hd__a21o_2 _13503_ (.A1(_04813_),
    .A2(_04835_),
    .B1(_05152_),
    .X(_05163_));
 sky130_fd_sc_hd__o211ai_2 _13504_ (.A1(_04802_),
    .A2(_04682_),
    .B1(_05152_),
    .C1(_04835_),
    .Y(_05174_));
 sky130_fd_sc_hd__o2111ai_4 _13505_ (.A1(_04846_),
    .A2(_04857_),
    .B1(_05174_),
    .C1(_04605_),
    .D1(_05163_),
    .Y(_05185_));
 sky130_fd_sc_hd__a2bb2o_1 _13506_ (.A1_N(_04616_),
    .A2_N(_04868_),
    .B1(_05163_),
    .B2(_05174_),
    .X(_05195_));
 sky130_fd_sc_hd__and2_1 _13507_ (.A(_05185_),
    .B(_05195_),
    .X(net109));
 sky130_fd_sc_hd__a31oi_1 _13508_ (.A1(_04943_),
    .A2(_04954_),
    .A3(_05130_),
    .B1(_05108_),
    .Y(_05216_));
 sky130_fd_sc_hd__and2b_4 _13509_ (.A_N(net59),
    .B(net60),
    .X(_05227_));
 sky130_fd_sc_hd__nand2b_4 _13510_ (.A_N(net59),
    .B(net60),
    .Y(_05238_));
 sky130_fd_sc_hd__and2b_4 _13511_ (.A_N(net60),
    .B(net59),
    .X(_05249_));
 sky130_fd_sc_hd__nand2b_4 _13512_ (.A_N(net60),
    .B(net59),
    .Y(_05260_));
 sky130_fd_sc_hd__a21oi_2 _13513_ (.A1(_05238_),
    .A2(_05260_),
    .B1(_03176_),
    .Y(_05271_));
 sky130_fd_sc_hd__o21ai_1 _13514_ (.A1(_04298_),
    .A2(_04506_),
    .B1(net305),
    .Y(_05282_));
 sky130_fd_sc_hd__nand2_1 _13515_ (.A(net12),
    .B(_04911_),
    .Y(_05293_));
 sky130_fd_sc_hd__nand3_1 _13516_ (.A(_04419_),
    .B(_04452_),
    .C(net317),
    .Y(_05304_));
 sky130_fd_sc_hd__nand2_1 _13517_ (.A(net23),
    .B(_04649_),
    .Y(_05315_));
 sky130_fd_sc_hd__a22oi_1 _13518_ (.A1(_05282_),
    .A2(_05293_),
    .B1(_05304_),
    .B2(_05315_),
    .Y(_05326_));
 sky130_fd_sc_hd__a22o_1 _13519_ (.A1(_05282_),
    .A2(_05293_),
    .B1(_05304_),
    .B2(_05315_),
    .X(_05337_));
 sky130_fd_sc_hd__nand4_2 _13520_ (.A(_05282_),
    .B(_05293_),
    .C(_05304_),
    .D(_05315_),
    .Y(_05348_));
 sky130_fd_sc_hd__a21bo_1 _13521_ (.A1(_05337_),
    .A2(_05348_),
    .B1_N(_05271_),
    .X(_05359_));
 sky130_fd_sc_hd__nand3b_1 _13522_ (.A_N(_05271_),
    .B(_05337_),
    .C(_05348_),
    .Y(_05370_));
 sky130_fd_sc_hd__nand2_1 _13523_ (.A(_05359_),
    .B(_05370_),
    .Y(_05381_));
 sky130_fd_sc_hd__a21boi_1 _13524_ (.A1(_04987_),
    .A2(_05075_),
    .B1_N(_05053_),
    .Y(_05392_));
 sky130_fd_sc_hd__a32o_1 _13525_ (.A1(net267),
    .A2(_04342_),
    .A3(net314),
    .B1(_04364_),
    .B2(net26),
    .X(_05403_));
 sky130_fd_sc_hd__a31o_4 _13526_ (.A1(_04397_),
    .A2(_04725_),
    .A3(_03616_),
    .B1(_03725_),
    .X(_05414_));
 sky130_fd_sc_hd__nor2_4 _13527_ (.A(net27),
    .B(net28),
    .Y(_05425_));
 sky130_fd_sc_hd__or2_4 _13528_ (.A(net27),
    .B(net28),
    .X(_05436_));
 sky130_fd_sc_hd__nand3_4 _13529_ (.A(_04397_),
    .B(_04725_),
    .C(_05425_),
    .Y(_05446_));
 sky130_fd_sc_hd__o21ai_4 _13530_ (.A1(net267),
    .A2(_05436_),
    .B1(_05414_),
    .Y(_05457_));
 sky130_fd_sc_hd__o211ai_1 _13531_ (.A1(net267),
    .A2(_05436_),
    .B1(net33),
    .C1(_05414_),
    .Y(_05468_));
 sky130_fd_sc_hd__a32oi_4 _13532_ (.A1(net300),
    .A2(_04484_),
    .A3(_04998_),
    .B1(_04320_),
    .B2(net27),
    .Y(_05479_));
 sky130_fd_sc_hd__o21ai_2 _13533_ (.A1(_03286_),
    .A2(_05457_),
    .B1(_05479_),
    .Y(_05490_));
 sky130_fd_sc_hd__and3_1 _13534_ (.A(net27),
    .B(_04320_),
    .C(_03725_),
    .X(_05501_));
 sky130_fd_sc_hd__or4_1 _13535_ (.A(net44),
    .B(net28),
    .C(_03616_),
    .D(_03286_),
    .X(_05512_));
 sky130_fd_sc_hd__nand3_1 _13536_ (.A(_05403_),
    .B(_05490_),
    .C(_05512_),
    .Y(_05523_));
 sky130_fd_sc_hd__a21o_1 _13537_ (.A1(_05490_),
    .A2(_05512_),
    .B1(_05403_),
    .X(_05534_));
 sky130_fd_sc_hd__a21bo_1 _13538_ (.A1(_05490_),
    .A2(_05512_),
    .B1_N(_05403_),
    .X(_05545_));
 sky130_fd_sc_hd__a211o_1 _13539_ (.A1(_05479_),
    .A2(_05468_),
    .B1(_05403_),
    .C1(_05501_),
    .X(_05556_));
 sky130_fd_sc_hd__nand3b_1 _13540_ (.A_N(_05392_),
    .B(_05523_),
    .C(_05534_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand3_1 _13541_ (.A(_05545_),
    .B(_05556_),
    .C(_05392_),
    .Y(_05578_));
 sky130_fd_sc_hd__nand3_1 _13542_ (.A(_05534_),
    .B(_05392_),
    .C(_05523_),
    .Y(_05589_));
 sky130_fd_sc_hd__nand3b_1 _13543_ (.A_N(_05392_),
    .B(_05545_),
    .C(_05556_),
    .Y(_05600_));
 sky130_fd_sc_hd__nand3_1 _13544_ (.A(_05567_),
    .B(_05578_),
    .C(_05381_),
    .Y(_05611_));
 sky130_fd_sc_hd__nand3b_1 _13545_ (.A_N(_05381_),
    .B(_05567_),
    .C(_05578_),
    .Y(_05622_));
 sky130_fd_sc_hd__nand3_1 _13546_ (.A(_05600_),
    .B(_05381_),
    .C(_05589_),
    .Y(_05633_));
 sky130_fd_sc_hd__o2111ai_1 _13547_ (.A1(_04965_),
    .A2(_05141_),
    .B1(_05622_),
    .C1(_05633_),
    .D1(_05119_),
    .Y(_05644_));
 sky130_fd_sc_hd__a21o_1 _13548_ (.A1(_05622_),
    .A2(_05633_),
    .B1(_05216_),
    .X(_05655_));
 sky130_fd_sc_hd__nand2_1 _13549_ (.A(_05644_),
    .B(_05655_),
    .Y(_05666_));
 sky130_fd_sc_hd__xnor2_2 _13550_ (.A(_04943_),
    .B(_05666_),
    .Y(_05677_));
 sky130_fd_sc_hd__and2b_4 _13551_ (.A_N(net60),
    .B(net61),
    .X(_05688_));
 sky130_fd_sc_hd__nand2b_4 _13552_ (.A_N(net60),
    .B(net61),
    .Y(_05699_));
 sky130_fd_sc_hd__and2b_2 _13553_ (.A_N(net61),
    .B(net60),
    .X(_05710_));
 sky130_fd_sc_hd__nand2b_4 _13554_ (.A_N(net61),
    .B(net60),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ai_2 _13555_ (.A1(net299),
    .A2(_05710_),
    .B1(net1),
    .Y(_05731_));
 sky130_fd_sc_hd__a21oi_2 _13556_ (.A1(_05348_),
    .A2(_05271_),
    .B1(_05326_),
    .Y(_05742_));
 sky130_fd_sc_hd__nor2_1 _13557_ (.A(_05731_),
    .B(_05742_),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(_05742_),
    .B(_05731_),
    .Y(_05764_));
 sky130_fd_sc_hd__nand2b_1 _13559_ (.A_N(_05753_),
    .B(_05764_),
    .Y(_05775_));
 sky130_fd_sc_hd__a21boi_1 _13560_ (.A1(_05381_),
    .A2(_05578_),
    .B1_N(_05567_),
    .Y(_05786_));
 sky130_fd_sc_hd__a2bb2o_1 _13561_ (.A1_N(_05403_),
    .A2_N(_05501_),
    .B1(_05479_),
    .B2(_05468_),
    .X(_05797_));
 sky130_fd_sc_hd__a32o_1 _13562_ (.A1(net27),
    .A2(_04320_),
    .A3(_03725_),
    .B1(_05490_),
    .B2(_05403_),
    .X(_05808_));
 sky130_fd_sc_hd__a32o_1 _13563_ (.A1(net300),
    .A2(_04342_),
    .A3(_04998_),
    .B1(_04364_),
    .B2(net27),
    .X(_05819_));
 sky130_fd_sc_hd__a31oi_4 _13564_ (.A1(_04397_),
    .A2(_04725_),
    .A3(_05425_),
    .B1(_03835_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_8 _13565_ (.A(_05446_),
    .B(net29),
    .Y(_05841_));
 sky130_fd_sc_hd__nor3_4 _13566_ (.A(net27),
    .B(net28),
    .C(net29),
    .Y(_05852_));
 sky130_fd_sc_hd__nand4_4 _13567_ (.A(_04397_),
    .B(_04725_),
    .C(_05425_),
    .D(_03835_),
    .Y(_05863_));
 sky130_fd_sc_hd__a21oi_4 _13568_ (.A1(net312),
    .A2(net297),
    .B1(_05830_),
    .Y(_05874_));
 sky130_fd_sc_hd__nand3_1 _13569_ (.A(_05841_),
    .B(_05863_),
    .C(net33),
    .Y(_05885_));
 sky130_fd_sc_hd__nand3_1 _13570_ (.A(_05414_),
    .B(_05446_),
    .C(_04484_),
    .Y(_05896_));
 sky130_fd_sc_hd__or3_1 _13571_ (.A(net44),
    .B(_03725_),
    .C(_03286_),
    .X(_05907_));
 sky130_fd_sc_hd__or4_2 _13572_ (.A(net44),
    .B(net29),
    .C(_03725_),
    .D(_03286_),
    .X(_05918_));
 sky130_fd_sc_hd__nand3_2 _13573_ (.A(_05885_),
    .B(_05896_),
    .C(_05907_),
    .Y(_05929_));
 sky130_fd_sc_hd__a21o_1 _13574_ (.A1(_05918_),
    .A2(_05929_),
    .B1(_05819_),
    .X(_05940_));
 sky130_fd_sc_hd__nand3_1 _13575_ (.A(_05819_),
    .B(_05918_),
    .C(_05929_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand3b_1 _13576_ (.A_N(_05819_),
    .B(_05918_),
    .C(_05929_),
    .Y(_05962_));
 sky130_fd_sc_hd__a21bo_1 _13577_ (.A1(_05918_),
    .A2(_05929_),
    .B1_N(_05819_),
    .X(_05973_));
 sky130_fd_sc_hd__nand3_2 _13578_ (.A(_05973_),
    .B(_05797_),
    .C(_05962_),
    .Y(_05984_));
 sky130_fd_sc_hd__inv_2 _13579_ (.A(_05984_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand3_1 _13580_ (.A(_05808_),
    .B(_05940_),
    .C(_05951_),
    .Y(_06006_));
 sky130_fd_sc_hd__o2bb2a_1 _13581_ (.A1_N(net12),
    .A2_N(_05249_),
    .B1(_05238_),
    .B2(_04528_),
    .X(_06017_));
 sky130_fd_sc_hd__a22o_1 _13582_ (.A1(net12),
    .A2(_05249_),
    .B1(_04539_),
    .B2(_05227_),
    .X(_06027_));
 sky130_fd_sc_hd__a22oi_2 _13583_ (.A1(_04463_),
    .A2(net305),
    .B1(_04911_),
    .B2(net23),
    .Y(_06038_));
 sky130_fd_sc_hd__a32o_1 _13584_ (.A1(_04419_),
    .A2(_04452_),
    .A3(net305),
    .B1(_04911_),
    .B2(net23),
    .X(_06049_));
 sky130_fd_sc_hd__a32o_1 _13585_ (.A1(net267),
    .A2(net317),
    .A3(net314),
    .B1(_04649_),
    .B2(net26),
    .X(_06060_));
 sky130_fd_sc_hd__nand2_1 _13586_ (.A(_06049_),
    .B(_06060_),
    .Y(_06071_));
 sky130_fd_sc_hd__o221ai_4 _13587_ (.A1(_03506_),
    .A2(_04660_),
    .B1(_04758_),
    .B2(_04638_),
    .C1(_06038_),
    .Y(_06082_));
 sky130_fd_sc_hd__and3_1 _13588_ (.A(_06071_),
    .B(_06082_),
    .C(_06017_),
    .X(_06093_));
 sky130_fd_sc_hd__nand3_1 _13589_ (.A(_06071_),
    .B(_06082_),
    .C(_06017_),
    .Y(_06104_));
 sky130_fd_sc_hd__a21oi_1 _13590_ (.A1(_06071_),
    .A2(_06082_),
    .B1(_06017_),
    .Y(_06115_));
 sky130_fd_sc_hd__a21o_1 _13591_ (.A1(_06071_),
    .A2(_06082_),
    .B1(_06017_),
    .X(_06126_));
 sky130_fd_sc_hd__nand2_1 _13592_ (.A(_06104_),
    .B(_06126_),
    .Y(_06137_));
 sky130_fd_sc_hd__o211a_1 _13593_ (.A1(_06093_),
    .A2(_06115_),
    .B1(_05984_),
    .C1(_06006_),
    .X(_06148_));
 sky130_fd_sc_hd__a21oi_1 _13594_ (.A1(_05984_),
    .A2(_06006_),
    .B1(_06137_),
    .Y(_06159_));
 sky130_fd_sc_hd__a211o_1 _13595_ (.A1(_05567_),
    .A2(_05611_),
    .B1(_06148_),
    .C1(_06159_),
    .X(_06170_));
 sky130_fd_sc_hd__o21a_1 _13596_ (.A1(_06148_),
    .A2(_06159_),
    .B1(_05786_),
    .X(_06181_));
 sky130_fd_sc_hd__o21ai_1 _13597_ (.A1(_06148_),
    .A2(_06159_),
    .B1(_05786_),
    .Y(_06192_));
 sky130_fd_sc_hd__nand3_1 _13598_ (.A(_05775_),
    .B(_06170_),
    .C(_06192_),
    .Y(_06203_));
 sky130_fd_sc_hd__a21o_1 _13599_ (.A1(_06170_),
    .A2(_06192_),
    .B1(_05775_),
    .X(_06214_));
 sky130_fd_sc_hd__and2_1 _13600_ (.A(_06203_),
    .B(_06214_),
    .X(_06225_));
 sky130_fd_sc_hd__a32o_1 _13601_ (.A1(_05216_),
    .A2(_05622_),
    .A3(_05633_),
    .B1(_05655_),
    .B2(_04943_),
    .X(_06236_));
 sky130_fd_sc_hd__a21oi_2 _13602_ (.A1(_06203_),
    .A2(_06214_),
    .B1(_06236_),
    .Y(_06247_));
 sky130_fd_sc_hd__nor2_1 _13603_ (.A(_05163_),
    .B(_05677_),
    .Y(_06258_));
 sky130_fd_sc_hd__xnor2_2 _13604_ (.A(_05163_),
    .B(_05677_),
    .Y(_06269_));
 sky130_fd_sc_hd__xor2_1 _13605_ (.A(_05185_),
    .B(_06269_),
    .X(net120));
 sky130_fd_sc_hd__nand2_1 _13606_ (.A(_06225_),
    .B(_06236_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand2b_1 _13607_ (.A_N(_06247_),
    .B(_06290_),
    .Y(_06301_));
 sky130_fd_sc_hd__o22a_1 _13608_ (.A1(_05163_),
    .A2(_05677_),
    .B1(_06269_),
    .B2(_05185_),
    .X(_06312_));
 sky130_fd_sc_hd__xor2_1 _13609_ (.A(_06301_),
    .B(_06312_),
    .X(net125));
 sky130_fd_sc_hd__o32a_1 _13610_ (.A1(_05238_),
    .A2(_04441_),
    .A3(_04408_),
    .B1(_03396_),
    .B2(_05260_),
    .X(_06332_));
 sky130_fd_sc_hd__nand3_1 _13611_ (.A(net314),
    .B(net267),
    .C(net305),
    .Y(_06343_));
 sky130_fd_sc_hd__nand2_1 _13612_ (.A(net26),
    .B(_04911_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand3_1 _13613_ (.A(net300),
    .B(net317),
    .C(_04998_),
    .Y(_06365_));
 sky130_fd_sc_hd__or3b_1 _13614_ (.A(net58),
    .B(_03616_),
    .C_N(net55),
    .X(_06376_));
 sky130_fd_sc_hd__a22oi_1 _13615_ (.A1(_06343_),
    .A2(_06354_),
    .B1(_06365_),
    .B2(_06376_),
    .Y(_06387_));
 sky130_fd_sc_hd__a22o_1 _13616_ (.A1(_06343_),
    .A2(_06354_),
    .B1(_06365_),
    .B2(_06376_),
    .X(_06398_));
 sky130_fd_sc_hd__o2111a_1 _13617_ (.A1(_03616_),
    .A2(_04660_),
    .B1(_06343_),
    .C1(_06354_),
    .D1(_06365_),
    .X(_06409_));
 sky130_fd_sc_hd__nor3_1 _13618_ (.A(_06332_),
    .B(_06387_),
    .C(_06409_),
    .Y(_06420_));
 sky130_fd_sc_hd__o21a_1 _13619_ (.A1(_06387_),
    .A2(_06409_),
    .B1(_06332_),
    .X(_06431_));
 sky130_fd_sc_hd__nor2_1 _13620_ (.A(_06420_),
    .B(_06431_),
    .Y(_06442_));
 sky130_fd_sc_hd__or3b_1 _13621_ (.A(net55),
    .B(_03725_),
    .C_N(net44),
    .X(_06453_));
 sky130_fd_sc_hd__o211ai_1 _13622_ (.A1(net267),
    .A2(_05436_),
    .B1(_04342_),
    .C1(_05414_),
    .Y(_06464_));
 sky130_fd_sc_hd__a32o_1 _13623_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_04342_),
    .B1(_04364_),
    .B2(net28),
    .X(_06475_));
 sky130_fd_sc_hd__nand2_8 _13624_ (.A(net265),
    .B(net30),
    .Y(_06486_));
 sky130_fd_sc_hd__nor4_4 _13625_ (.A(net27),
    .B(net28),
    .C(net29),
    .D(net30),
    .Y(_06497_));
 sky130_fd_sc_hd__nand3_4 _13626_ (.A(_05425_),
    .B(_03916_),
    .C(_03835_),
    .Y(_06508_));
 sky130_fd_sc_hd__nor2_8 _13627_ (.A(net267),
    .B(_06508_),
    .Y(_06519_));
 sky130_fd_sc_hd__nand4_4 _13628_ (.A(_04441_),
    .B(_05852_),
    .C(_03506_),
    .D(_03916_),
    .Y(_06530_));
 sky130_fd_sc_hd__a22oi_4 _13629_ (.A1(net309),
    .A2(net295),
    .B1(_05863_),
    .B2(net30),
    .Y(_06541_));
 sky130_fd_sc_hd__a32o_4 _13630_ (.A1(_06497_),
    .A2(_03506_),
    .A3(_04441_),
    .B1(_05863_),
    .B2(net30),
    .X(_06552_));
 sky130_fd_sc_hd__o211ai_1 _13631_ (.A1(net267),
    .A2(_06508_),
    .B1(net33),
    .C1(_06486_),
    .Y(_06563_));
 sky130_fd_sc_hd__nor2_1 _13632_ (.A(_03835_),
    .B(_04331_),
    .Y(_06574_));
 sky130_fd_sc_hd__or3_1 _13633_ (.A(net44),
    .B(_03835_),
    .C(_03286_),
    .X(_06585_));
 sky130_fd_sc_hd__nand3_1 _13634_ (.A(_05841_),
    .B(_05863_),
    .C(_04484_),
    .Y(_06596_));
 sky130_fd_sc_hd__nand3_2 _13635_ (.A(_06563_),
    .B(_06585_),
    .C(_06596_),
    .Y(_06607_));
 sky130_fd_sc_hd__nand4_1 _13636_ (.A(_06486_),
    .B(_06530_),
    .C(_06574_),
    .D(net33),
    .Y(_06618_));
 sky130_fd_sc_hd__a21oi_1 _13637_ (.A1(_06607_),
    .A2(_06618_),
    .B1(_06475_),
    .Y(_06628_));
 sky130_fd_sc_hd__a21o_1 _13638_ (.A1(_06607_),
    .A2(_06618_),
    .B1(_06475_),
    .X(_06639_));
 sky130_fd_sc_hd__a32oi_2 _13639_ (.A1(net33),
    .A2(_06541_),
    .A3(_06574_),
    .B1(_06453_),
    .B2(_06464_),
    .Y(_06650_));
 sky130_fd_sc_hd__nand2_1 _13640_ (.A(_06650_),
    .B(_06607_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand2_1 _13641_ (.A(_05819_),
    .B(_05929_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_1 _13642_ (.A(_05918_),
    .B(_06672_),
    .Y(_06683_));
 sky130_fd_sc_hd__a221oi_2 _13643_ (.A1(_06650_),
    .A2(_06607_),
    .B1(_05918_),
    .B2(_06672_),
    .C1(_06628_),
    .Y(_06694_));
 sky130_fd_sc_hd__nand3_1 _13644_ (.A(_06683_),
    .B(_06661_),
    .C(_06639_),
    .Y(_06705_));
 sky130_fd_sc_hd__a21oi_1 _13645_ (.A1(_06639_),
    .A2(_06661_),
    .B1(_06683_),
    .Y(_06716_));
 sky130_fd_sc_hd__a21o_1 _13646_ (.A1(_06639_),
    .A2(_06661_),
    .B1(_06683_),
    .X(_06727_));
 sky130_fd_sc_hd__nand3_2 _13647_ (.A(_06727_),
    .B(_06442_),
    .C(_06705_),
    .Y(_06738_));
 sky130_fd_sc_hd__inv_2 _13648_ (.A(_06738_),
    .Y(_06749_));
 sky130_fd_sc_hd__o22ai_2 _13649_ (.A1(_06420_),
    .A2(_06431_),
    .B1(_06694_),
    .B2(_06716_),
    .Y(_06760_));
 sky130_fd_sc_hd__a311oi_2 _13650_ (.A1(_05808_),
    .A2(_05940_),
    .A3(_05951_),
    .B1(_06093_),
    .C1(_06115_),
    .Y(_06771_));
 sky130_fd_sc_hd__a21bo_1 _13651_ (.A1(_05984_),
    .A2(_06137_),
    .B1_N(_06006_),
    .X(_06782_));
 sky130_fd_sc_hd__o2bb2ai_2 _13652_ (.A1_N(_06738_),
    .A2_N(_06760_),
    .B1(_06771_),
    .B2(_05995_),
    .Y(_06793_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(_06782_),
    .B(_06760_),
    .Y(_06804_));
 sky130_fd_sc_hd__nand3_1 _13654_ (.A(_06782_),
    .B(_06760_),
    .C(_06738_),
    .Y(_06815_));
 sky130_fd_sc_hd__and2b_4 _13655_ (.A_N(net61),
    .B(net62),
    .X(_06826_));
 sky130_fd_sc_hd__nand2b_4 _13656_ (.A_N(net61),
    .B(net62),
    .Y(_06837_));
 sky130_fd_sc_hd__and2b_4 _13657_ (.A_N(net62),
    .B(net61),
    .X(_06848_));
 sky130_fd_sc_hd__nand2_8 _13658_ (.A(_03927_),
    .B(net61),
    .Y(_06859_));
 sky130_fd_sc_hd__a21oi_4 _13659_ (.A1(_06837_),
    .A2(_06859_),
    .B1(_03176_),
    .Y(_06870_));
 sky130_fd_sc_hd__a22o_1 _13660_ (.A1(net12),
    .A2(_05710_),
    .B1(_04539_),
    .B2(net299),
    .X(_06881_));
 sky130_fd_sc_hd__nand2_1 _13661_ (.A(_06881_),
    .B(_06870_),
    .Y(_06892_));
 sky130_fd_sc_hd__a221o_1 _13662_ (.A1(_04539_),
    .A2(net299),
    .B1(_05710_),
    .B2(net12),
    .C1(_06870_),
    .X(_06903_));
 sky130_fd_sc_hd__nand2_1 _13663_ (.A(_06892_),
    .B(_06903_),
    .Y(_06914_));
 sky130_fd_sc_hd__a21boi_2 _13664_ (.A1(_06027_),
    .A2(_06082_),
    .B1_N(_06071_),
    .Y(_06925_));
 sky130_fd_sc_hd__nor2_1 _13665_ (.A(_06914_),
    .B(_06925_),
    .Y(_06936_));
 sky130_fd_sc_hd__and2_1 _13666_ (.A(_06914_),
    .B(_06925_),
    .X(_06946_));
 sky130_fd_sc_hd__nor2_1 _13667_ (.A(_06936_),
    .B(_06946_),
    .Y(_06957_));
 sky130_fd_sc_hd__o2bb2ai_1 _13668_ (.A1_N(_06793_),
    .A2_N(_06815_),
    .B1(_06936_),
    .B2(_06946_),
    .Y(_06968_));
 sky130_fd_sc_hd__nand3_1 _13669_ (.A(_06793_),
    .B(_06815_),
    .C(_06957_),
    .Y(_06979_));
 sky130_fd_sc_hd__o21ai_1 _13670_ (.A1(_05775_),
    .A2(_06181_),
    .B1(_06170_),
    .Y(_06990_));
 sky130_fd_sc_hd__a21o_1 _13671_ (.A1(_06968_),
    .A2(_06979_),
    .B1(_06990_),
    .X(_07001_));
 sky130_fd_sc_hd__nand3_2 _13672_ (.A(_06990_),
    .B(_06979_),
    .C(_06968_),
    .Y(_07012_));
 sky130_fd_sc_hd__o2bb2ai_2 _13673_ (.A1_N(_07001_),
    .A2_N(_07012_),
    .B1(_05731_),
    .B2(_05742_),
    .Y(_07023_));
 sky130_fd_sc_hd__nand3_2 _13674_ (.A(_07001_),
    .B(_07012_),
    .C(_05753_),
    .Y(_07034_));
 sky130_fd_sc_hd__and4_1 _13675_ (.A(_06258_),
    .B(_06290_),
    .C(_07023_),
    .D(_07034_),
    .X(_07045_));
 sky130_fd_sc_hd__inv_2 _13676_ (.A(_07045_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand3_1 _13677_ (.A(_07023_),
    .B(_07034_),
    .C(_06247_),
    .Y(_07067_));
 sky130_fd_sc_hd__inv_2 _13678_ (.A(_07067_),
    .Y(_07078_));
 sky130_fd_sc_hd__a2bb2o_1 _13679_ (.A1_N(_06225_),
    .A2_N(_06236_),
    .B1(_07023_),
    .B2(_07034_),
    .X(_07089_));
 sky130_fd_sc_hd__a22o_1 _13680_ (.A1(_06290_),
    .A2(_06258_),
    .B1(_07089_),
    .B2(_07067_),
    .X(_07100_));
 sky130_fd_sc_hd__and2_1 _13681_ (.A(_07056_),
    .B(_07100_),
    .X(_07111_));
 sky130_fd_sc_hd__nor3_1 _13682_ (.A(_05185_),
    .B(_06269_),
    .C(_06301_),
    .Y(_07122_));
 sky130_fd_sc_hd__or4b_1 _13683_ (.A(_05185_),
    .B(_06269_),
    .C(_06301_),
    .D_N(_07111_),
    .X(_07133_));
 sky130_fd_sc_hd__xor2_1 _13684_ (.A(_07111_),
    .B(_07122_),
    .X(net126));
 sky130_fd_sc_hd__a21bo_2 _13685_ (.A1(_07001_),
    .A2(_05753_),
    .B1_N(_07012_),
    .X(_07154_));
 sky130_fd_sc_hd__a21boi_1 _13686_ (.A1(_07001_),
    .A2(_05753_),
    .B1_N(_07012_),
    .Y(_07165_));
 sky130_fd_sc_hd__a21oi_1 _13687_ (.A1(_06727_),
    .A2(_06442_),
    .B1(_06694_),
    .Y(_07176_));
 sky130_fd_sc_hd__a21o_1 _13688_ (.A1(_06727_),
    .A2(_06442_),
    .B1(_06694_),
    .X(_07187_));
 sky130_fd_sc_hd__and3_1 _13689_ (.A(_05841_),
    .B(_05863_),
    .C(_04342_),
    .X(_07198_));
 sky130_fd_sc_hd__nor2_1 _13690_ (.A(_03835_),
    .B(_04375_),
    .Y(_07209_));
 sky130_fd_sc_hd__a31o_1 _13691_ (.A1(_05841_),
    .A2(_05863_),
    .A3(_04342_),
    .B1(_07209_),
    .X(_07220_));
 sky130_fd_sc_hd__a41oi_2 _13692_ (.A1(_04441_),
    .A2(_05852_),
    .A3(_03506_),
    .A4(_03916_),
    .B1(_03938_),
    .Y(_07231_));
 sky130_fd_sc_hd__a41o_4 _13693_ (.A1(_04441_),
    .A2(_05852_),
    .A3(_03506_),
    .A4(_03916_),
    .B1(_03938_),
    .X(_07242_));
 sky130_fd_sc_hd__nand4_4 _13694_ (.A(_04736_),
    .B(_05852_),
    .C(_03916_),
    .D(_03938_),
    .Y(_07253_));
 sky130_fd_sc_hd__nand2_8 _13695_ (.A(_07242_),
    .B(net258),
    .Y(_07263_));
 sky130_fd_sc_hd__nand3_1 _13696_ (.A(_07242_),
    .B(net258),
    .C(net33),
    .Y(_07274_));
 sky130_fd_sc_hd__o211ai_1 _13697_ (.A1(net267),
    .A2(_06508_),
    .B1(_04484_),
    .C1(_06486_),
    .Y(_07285_));
 sky130_fd_sc_hd__nor2_1 _13698_ (.A(_03916_),
    .B(_04331_),
    .Y(_07296_));
 sky130_fd_sc_hd__or3_1 _13699_ (.A(net44),
    .B(_03916_),
    .C(_03286_),
    .X(_07307_));
 sky130_fd_sc_hd__and4_1 _13700_ (.A(_07242_),
    .B(net258),
    .C(_07296_),
    .D(net33),
    .X(_07318_));
 sky130_fd_sc_hd__nand4_2 _13701_ (.A(_07242_),
    .B(net258),
    .C(_07296_),
    .D(net33),
    .Y(_07329_));
 sky130_fd_sc_hd__nand3_2 _13702_ (.A(_07274_),
    .B(_07285_),
    .C(_07307_),
    .Y(_07340_));
 sky130_fd_sc_hd__a21oi_1 _13703_ (.A1(_07329_),
    .A2(_07340_),
    .B1(_07220_),
    .Y(_07351_));
 sky130_fd_sc_hd__a21o_1 _13704_ (.A1(_07329_),
    .A2(_07340_),
    .B1(_07220_),
    .X(_07362_));
 sky130_fd_sc_hd__o211a_1 _13705_ (.A1(_07198_),
    .A2(_07209_),
    .B1(_07329_),
    .C1(_07340_),
    .X(_07373_));
 sky130_fd_sc_hd__o211ai_2 _13706_ (.A1(_07198_),
    .A2(_07209_),
    .B1(_07329_),
    .C1(_07340_),
    .Y(_07384_));
 sky130_fd_sc_hd__a32o_1 _13707_ (.A1(net33),
    .A2(_06541_),
    .A3(_06574_),
    .B1(_06607_),
    .B2(_06475_),
    .X(_07395_));
 sky130_fd_sc_hd__o21bai_4 _13708_ (.A1(_07351_),
    .A2(_07373_),
    .B1_N(_07395_),
    .Y(_07406_));
 sky130_fd_sc_hd__nand3_4 _13709_ (.A(_07362_),
    .B(_07384_),
    .C(_07395_),
    .Y(_07417_));
 sky130_fd_sc_hd__o32a_4 _13710_ (.A1(_05238_),
    .A2(_04736_),
    .A3(_04703_),
    .B1(_03506_),
    .B2(_05260_),
    .X(_07428_));
 sky130_fd_sc_hd__a32oi_4 _13711_ (.A1(net300),
    .A2(net305),
    .A3(_04998_),
    .B1(_04911_),
    .B2(net27),
    .Y(_07439_));
 sky130_fd_sc_hd__o211ai_2 _13712_ (.A1(net267),
    .A2(_05436_),
    .B1(net317),
    .C1(_05414_),
    .Y(_07450_));
 sky130_fd_sc_hd__or3b_2 _13713_ (.A(net58),
    .B(_03725_),
    .C_N(net55),
    .X(_07461_));
 sky130_fd_sc_hd__a21oi_2 _13714_ (.A1(_07450_),
    .A2(_07461_),
    .B1(_07439_),
    .Y(_07472_));
 sky130_fd_sc_hd__a21o_1 _13715_ (.A1(_07450_),
    .A2(_07461_),
    .B1(_07439_),
    .X(_07483_));
 sky130_fd_sc_hd__o221a_1 _13716_ (.A1(_03725_),
    .A2(_04660_),
    .B1(_05457_),
    .B2(_04638_),
    .C1(_07439_),
    .X(_07494_));
 sky130_fd_sc_hd__o221ai_4 _13717_ (.A1(_03725_),
    .A2(_04660_),
    .B1(_05457_),
    .B2(_04638_),
    .C1(_07439_),
    .Y(_07505_));
 sky130_fd_sc_hd__o21a_1 _13718_ (.A1(_07472_),
    .A2(_07494_),
    .B1(_07428_),
    .X(_07516_));
 sky130_fd_sc_hd__nor3_1 _13719_ (.A(_07428_),
    .B(_07472_),
    .C(_07494_),
    .Y(_07527_));
 sky130_fd_sc_hd__a21oi_1 _13720_ (.A1(_07483_),
    .A2(_07505_),
    .B1(_07428_),
    .Y(_07538_));
 sky130_fd_sc_hd__a21o_1 _13721_ (.A1(_07483_),
    .A2(_07505_),
    .B1(_07428_),
    .X(_07549_));
 sky130_fd_sc_hd__and3_1 _13722_ (.A(_07483_),
    .B(_07505_),
    .C(_07428_),
    .X(_07560_));
 sky130_fd_sc_hd__nand3_1 _13723_ (.A(_07483_),
    .B(_07505_),
    .C(_07428_),
    .Y(_07571_));
 sky130_fd_sc_hd__nand2_1 _13724_ (.A(_07549_),
    .B(_07571_),
    .Y(_07582_));
 sky130_fd_sc_hd__o2bb2ai_1 _13725_ (.A1_N(_07406_),
    .A2_N(_07417_),
    .B1(_07516_),
    .B2(_07527_),
    .Y(_07593_));
 sky130_fd_sc_hd__nand3_2 _13726_ (.A(_07406_),
    .B(_07417_),
    .C(_07582_),
    .Y(_07603_));
 sky130_fd_sc_hd__nand4_1 _13727_ (.A(_07406_),
    .B(_07417_),
    .C(_07549_),
    .D(_07571_),
    .Y(_07614_));
 sky130_fd_sc_hd__o2bb2ai_1 _13728_ (.A1_N(_07406_),
    .A2_N(_07417_),
    .B1(_07538_),
    .B2(_07560_),
    .Y(_07625_));
 sky130_fd_sc_hd__nand3_2 _13729_ (.A(_07625_),
    .B(_07176_),
    .C(_07614_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand3_2 _13730_ (.A(_07187_),
    .B(_07593_),
    .C(_07603_),
    .Y(_07647_));
 sky130_fd_sc_hd__and2_4 _13731_ (.A(_03927_),
    .B(net63),
    .X(_07658_));
 sky130_fd_sc_hd__nand2_8 _13732_ (.A(_03927_),
    .B(net63),
    .Y(_07669_));
 sky130_fd_sc_hd__nor2_8 _13733_ (.A(net63),
    .B(_03927_),
    .Y(_07680_));
 sky130_fd_sc_hd__or2_4 _13734_ (.A(net63),
    .B(_03927_),
    .X(_07691_));
 sky130_fd_sc_hd__nor2_1 _13735_ (.A(_07658_),
    .B(_07680_),
    .Y(_07702_));
 sky130_fd_sc_hd__a22oi_2 _13736_ (.A1(net12),
    .A2(_06848_),
    .B1(_04539_),
    .B2(net292),
    .Y(_07713_));
 sky130_fd_sc_hd__o2bb2ai_1 _13737_ (.A1_N(net12),
    .A2_N(_06848_),
    .B1(_06837_),
    .B2(_04528_),
    .Y(_07724_));
 sky130_fd_sc_hd__nand2_1 _13738_ (.A(net23),
    .B(_05710_),
    .Y(_07735_));
 sky130_fd_sc_hd__o31ai_1 _13739_ (.A1(_05699_),
    .A2(_04441_),
    .A3(_04408_),
    .B1(_07735_),
    .Y(_07746_));
 sky130_fd_sc_hd__o221a_1 _13740_ (.A1(_04474_),
    .A2(_05699_),
    .B1(net298),
    .B2(_03396_),
    .C1(_07713_),
    .X(_07757_));
 sky130_fd_sc_hd__o211ai_4 _13741_ (.A1(_04474_),
    .A2(_05699_),
    .B1(_07735_),
    .C1(_07713_),
    .Y(_07768_));
 sky130_fd_sc_hd__nand2_2 _13742_ (.A(_07724_),
    .B(_07746_),
    .Y(_07779_));
 sky130_fd_sc_hd__o2111ai_4 _13743_ (.A1(_07658_),
    .A2(_07680_),
    .B1(net1),
    .C1(_07768_),
    .D1(_07779_),
    .Y(_07790_));
 sky130_fd_sc_hd__o2bb2ai_2 _13744_ (.A1_N(_07768_),
    .A2_N(_07779_),
    .B1(_03176_),
    .B2(_07702_),
    .Y(_07801_));
 sky130_fd_sc_hd__o21ai_2 _13745_ (.A1(_06332_),
    .A2(_06409_),
    .B1(_06398_),
    .Y(_07812_));
 sky130_fd_sc_hd__a21oi_2 _13746_ (.A1(_07790_),
    .A2(_07801_),
    .B1(_07812_),
    .Y(_07823_));
 sky130_fd_sc_hd__a21o_1 _13747_ (.A1(_07790_),
    .A2(_07801_),
    .B1(_07812_),
    .X(_07834_));
 sky130_fd_sc_hd__and2_1 _13748_ (.A(_07812_),
    .B(_07801_),
    .X(_07845_));
 sky130_fd_sc_hd__and3_4 _13749_ (.A(_07812_),
    .B(_07801_),
    .C(_07790_),
    .X(_07856_));
 sky130_fd_sc_hd__o2bb2a_1 _13750_ (.A1_N(_06870_),
    .A2_N(_06881_),
    .B1(_07823_),
    .B2(_07856_),
    .X(_07867_));
 sky130_fd_sc_hd__o21ai_1 _13751_ (.A1(_07823_),
    .A2(_07856_),
    .B1(_06892_),
    .Y(_07878_));
 sky130_fd_sc_hd__nor3_1 _13752_ (.A(_06892_),
    .B(_07823_),
    .C(_07856_),
    .Y(_07889_));
 sky130_fd_sc_hd__a211o_1 _13753_ (.A1(_07845_),
    .A2(_07790_),
    .B1(_06892_),
    .C1(_07823_),
    .X(_07900_));
 sky130_fd_sc_hd__o211a_1 _13754_ (.A1(_07823_),
    .A2(_07856_),
    .B1(_06870_),
    .C1(_06881_),
    .X(_07911_));
 sky130_fd_sc_hd__a211oi_1 _13755_ (.A1(_06870_),
    .A2(_06881_),
    .B1(_07823_),
    .C1(_07856_),
    .Y(_07922_));
 sky130_fd_sc_hd__nor2_1 _13756_ (.A(_07867_),
    .B(_07889_),
    .Y(_07933_));
 sky130_fd_sc_hd__nand2_1 _13757_ (.A(_07878_),
    .B(_07900_),
    .Y(_07944_));
 sky130_fd_sc_hd__o2bb2ai_1 _13758_ (.A1_N(_07636_),
    .A2_N(_07647_),
    .B1(_07867_),
    .B2(_07889_),
    .Y(_07955_));
 sky130_fd_sc_hd__o211ai_1 _13759_ (.A1(_07911_),
    .A2(_07922_),
    .B1(_07636_),
    .C1(_07647_),
    .Y(_07965_));
 sky130_fd_sc_hd__o211ai_1 _13760_ (.A1(_07867_),
    .A2(_07889_),
    .B1(_07636_),
    .C1(_07647_),
    .Y(_07976_));
 sky130_fd_sc_hd__o2bb2ai_1 _13761_ (.A1_N(_07636_),
    .A2_N(_07647_),
    .B1(_07911_),
    .B2(_07922_),
    .Y(_07987_));
 sky130_fd_sc_hd__a21boi_1 _13762_ (.A1(_06793_),
    .A2(_06957_),
    .B1_N(_06815_),
    .Y(_07998_));
 sky130_fd_sc_hd__o2bb2ai_1 _13763_ (.A1_N(_06957_),
    .A2_N(_06793_),
    .B1(_06749_),
    .B2(_06804_),
    .Y(_08009_));
 sky130_fd_sc_hd__nand3_2 _13764_ (.A(_07998_),
    .B(_07987_),
    .C(_07976_),
    .Y(_08020_));
 sky130_fd_sc_hd__nand3_2 _13765_ (.A(_07955_),
    .B(_07965_),
    .C(_08009_),
    .Y(_08031_));
 sky130_fd_sc_hd__nand3_1 _13766_ (.A(_08020_),
    .B(_08031_),
    .C(_06936_),
    .Y(_08042_));
 sky130_fd_sc_hd__a2bb2o_1 _13767_ (.A1_N(_06914_),
    .A2_N(_06925_),
    .B1(_08020_),
    .B2(_08031_),
    .X(_08053_));
 sky130_fd_sc_hd__a21bo_1 _13768_ (.A1(_08020_),
    .A2(_08031_),
    .B1_N(_06936_),
    .X(_08064_));
 sky130_fd_sc_hd__o211ai_2 _13769_ (.A1(_06914_),
    .A2(_06925_),
    .B1(_08020_),
    .C1(_08031_),
    .Y(_08075_));
 sky130_fd_sc_hd__nand2_2 _13770_ (.A(_08064_),
    .B(_08075_),
    .Y(_08086_));
 sky130_fd_sc_hd__nand3_2 _13771_ (.A(_07154_),
    .B(_08042_),
    .C(_08053_),
    .Y(_08097_));
 sky130_fd_sc_hd__and3_1 _13772_ (.A(_07165_),
    .B(_08064_),
    .C(_08075_),
    .X(_08108_));
 sky130_fd_sc_hd__nand3_2 _13773_ (.A(_07165_),
    .B(_08064_),
    .C(_08075_),
    .Y(_08119_));
 sky130_fd_sc_hd__a32oi_2 _13774_ (.A1(_06247_),
    .A2(_07023_),
    .A3(_07034_),
    .B1(_08097_),
    .B2(_08119_),
    .Y(_08130_));
 sky130_fd_sc_hd__a32o_1 _13775_ (.A1(_06247_),
    .A2(_07023_),
    .A3(_07034_),
    .B1(_08097_),
    .B2(_08119_),
    .X(_08141_));
 sky130_fd_sc_hd__a21oi_1 _13776_ (.A1(_07078_),
    .A2(_08119_),
    .B1(_08130_),
    .Y(_08152_));
 sky130_fd_sc_hd__nand2_1 _13777_ (.A(_08141_),
    .B(_07045_),
    .Y(_08163_));
 sky130_fd_sc_hd__xor2_1 _13778_ (.A(_07056_),
    .B(_08152_),
    .X(_08174_));
 sky130_fd_sc_hd__nand4_1 _13779_ (.A(_08152_),
    .B(_07100_),
    .C(_07056_),
    .D(_07122_),
    .Y(_08185_));
 sky130_fd_sc_hd__nand2_1 _13780_ (.A(_07133_),
    .B(_08174_),
    .Y(_08196_));
 sky130_fd_sc_hd__and2_1 _13781_ (.A(_08185_),
    .B(_08196_),
    .X(net127));
 sky130_fd_sc_hd__nand2_1 _13782_ (.A(_08020_),
    .B(_06936_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_1 _13783_ (.A(_08031_),
    .B(_08217_),
    .Y(_08228_));
 sky130_fd_sc_hd__a21boi_1 _13784_ (.A1(_08020_),
    .A2(_06936_),
    .B1_N(_08031_),
    .Y(_08239_));
 sky130_fd_sc_hd__and2b_4 _13785_ (.A_N(net63),
    .B(net64),
    .X(_08250_));
 sky130_fd_sc_hd__nand2b_4 _13786_ (.A_N(net63),
    .B(net64),
    .Y(_08261_));
 sky130_fd_sc_hd__and2b_4 _13787_ (.A_N(net64),
    .B(net63),
    .X(_08272_));
 sky130_fd_sc_hd__nand2b_4 _13788_ (.A_N(net64),
    .B(net63),
    .Y(_08283_));
 sky130_fd_sc_hd__a21oi_4 _13789_ (.A1(_08261_),
    .A2(_08283_),
    .B1(_03176_),
    .Y(_08294_));
 sky130_fd_sc_hd__and3_2 _13790_ (.A(_07834_),
    .B(_06870_),
    .C(_06881_),
    .X(_08305_));
 sky130_fd_sc_hd__o221a_1 _13791_ (.A1(_08250_),
    .A2(_08272_),
    .B1(_08305_),
    .B2(_07856_),
    .C1(net1),
    .X(_08316_));
 sky130_fd_sc_hd__o21ai_2 _13792_ (.A1(_07856_),
    .A2(_08305_),
    .B1(_08294_),
    .Y(_08327_));
 sky130_fd_sc_hd__a311o_1 _13793_ (.A1(_07834_),
    .A2(_06870_),
    .A3(_06881_),
    .B1(_07856_),
    .C1(_08294_),
    .X(_08338_));
 sky130_fd_sc_hd__and2_1 _13794_ (.A(_08327_),
    .B(_08338_),
    .X(_08349_));
 sky130_fd_sc_hd__nand2_1 _13795_ (.A(_08327_),
    .B(_08338_),
    .Y(_08359_));
 sky130_fd_sc_hd__a32oi_2 _13796_ (.A1(_07187_),
    .A2(_07593_),
    .A3(_07603_),
    .B1(_07933_),
    .B2(_07636_),
    .Y(_08370_));
 sky130_fd_sc_hd__a21boi_1 _13797_ (.A1(_07647_),
    .A2(_07944_),
    .B1_N(_07636_),
    .Y(_08381_));
 sky130_fd_sc_hd__a32o_1 _13798_ (.A1(_04998_),
    .A2(net300),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net27),
    .X(_08392_));
 sky130_fd_sc_hd__a31oi_4 _13799_ (.A1(_04397_),
    .A2(_04725_),
    .A3(_05425_),
    .B1(_04900_),
    .Y(_08403_));
 sky130_fd_sc_hd__a22oi_2 _13800_ (.A1(net28),
    .A2(_04911_),
    .B1(_05414_),
    .B2(_08403_),
    .Y(_08414_));
 sky130_fd_sc_hd__a22o_1 _13801_ (.A1(net28),
    .A2(_04911_),
    .B1(_05414_),
    .B2(_08403_),
    .X(_08425_));
 sky130_fd_sc_hd__a31o_1 _13802_ (.A1(_04441_),
    .A2(net297),
    .A3(_03506_),
    .B1(_04638_),
    .X(_08436_));
 sky130_fd_sc_hd__nand3_1 _13803_ (.A(_05841_),
    .B(_05863_),
    .C(net317),
    .Y(_08447_));
 sky130_fd_sc_hd__o22ai_2 _13804_ (.A1(_03835_),
    .A2(net316),
    .B1(_05830_),
    .B2(_08436_),
    .Y(_08458_));
 sky130_fd_sc_hd__nand2_1 _13805_ (.A(_08425_),
    .B(_08458_),
    .Y(_08469_));
 sky130_fd_sc_hd__o211a_1 _13806_ (.A1(_03835_),
    .A2(_04660_),
    .B1(_08447_),
    .C1(_08414_),
    .X(_08480_));
 sky130_fd_sc_hd__o211ai_2 _13807_ (.A1(_03835_),
    .A2(_04660_),
    .B1(_08447_),
    .C1(_08414_),
    .Y(_08491_));
 sky130_fd_sc_hd__a21oi_1 _13808_ (.A1(_08469_),
    .A2(_08491_),
    .B1(_08392_),
    .Y(_08502_));
 sky130_fd_sc_hd__and3_1 _13809_ (.A(_08392_),
    .B(_08469_),
    .C(_08491_),
    .X(_08513_));
 sky130_fd_sc_hd__and3b_1 _13810_ (.A_N(_08392_),
    .B(_08469_),
    .C(_08491_),
    .X(_08524_));
 sky130_fd_sc_hd__a21boi_1 _13811_ (.A1(_08469_),
    .A2(_08491_),
    .B1_N(_08392_),
    .Y(_08535_));
 sky130_fd_sc_hd__nor2_1 _13812_ (.A(_08502_),
    .B(_08513_),
    .Y(_08546_));
 sky130_fd_sc_hd__a21oi_1 _13813_ (.A1(_07220_),
    .A2(_07340_),
    .B1(_07318_),
    .Y(_08557_));
 sky130_fd_sc_hd__nor2_1 _13814_ (.A(_03916_),
    .B(_04375_),
    .Y(_08568_));
 sky130_fd_sc_hd__o311a_1 _13815_ (.A1(net26),
    .A2(_04452_),
    .A3(_06508_),
    .B1(_04342_),
    .C1(_06486_),
    .X(_08579_));
 sky130_fd_sc_hd__a31o_2 _13816_ (.A1(_06486_),
    .A2(_06530_),
    .A3(_04342_),
    .B1(_08568_),
    .X(_08590_));
 sky130_fd_sc_hd__nor2_1 _13817_ (.A(_03938_),
    .B(_04331_),
    .Y(_08601_));
 sky130_fd_sc_hd__or3_1 _13818_ (.A(net44),
    .B(net32),
    .C(_03286_),
    .X(_08612_));
 sky130_fd_sc_hd__and3_2 _13819_ (.A(net31),
    .B(_04320_),
    .C(_03949_),
    .X(_08623_));
 sky130_fd_sc_hd__or4_1 _13820_ (.A(net44),
    .B(net32),
    .C(_03938_),
    .D(_03286_),
    .X(_08634_));
 sky130_fd_sc_hd__nor2_8 _13821_ (.A(net31),
    .B(net32),
    .Y(_08645_));
 sky130_fd_sc_hd__or2_4 _13822_ (.A(net31),
    .B(net32),
    .X(_08656_));
 sky130_fd_sc_hd__and3_2 _13823_ (.A(net311),
    .B(net295),
    .C(_08645_),
    .X(_08667_));
 sky130_fd_sc_hd__nand4_2 _13824_ (.A(net311),
    .B(net297),
    .C(_08645_),
    .D(_03916_),
    .Y(_08678_));
 sky130_fd_sc_hd__a41oi_4 _13825_ (.A1(net309),
    .A2(net297),
    .A3(_03916_),
    .A4(_03938_),
    .B1(_03949_),
    .Y(_08689_));
 sky130_fd_sc_hd__a41o_4 _13826_ (.A1(_04736_),
    .A2(_05852_),
    .A3(_03916_),
    .A4(_03938_),
    .B1(_03949_),
    .X(_08700_));
 sky130_fd_sc_hd__o21ai_4 _13827_ (.A1(_06530_),
    .A2(_08656_),
    .B1(_08700_),
    .Y(_08711_));
 sky130_fd_sc_hd__o211ai_4 _13828_ (.A1(_06530_),
    .A2(_08656_),
    .B1(net33),
    .C1(_08700_),
    .Y(_08722_));
 sky130_fd_sc_hd__a31oi_4 _13829_ (.A1(_07242_),
    .A2(net258),
    .A3(_04484_),
    .B1(_08601_),
    .Y(_08733_));
 sky130_fd_sc_hd__nand2_2 _13830_ (.A(_08733_),
    .B(_08722_),
    .Y(_08744_));
 sky130_fd_sc_hd__a21oi_1 _13831_ (.A1(_08733_),
    .A2(_08722_),
    .B1(_08623_),
    .Y(_08754_));
 sky130_fd_sc_hd__o2bb2ai_1 _13832_ (.A1_N(_08722_),
    .A2_N(_08733_),
    .B1(_03938_),
    .B2(_08612_),
    .Y(_08765_));
 sky130_fd_sc_hd__o311a_1 _13833_ (.A1(_03938_),
    .A2(net32),
    .A3(_04331_),
    .B1(_08590_),
    .C1(_08744_),
    .X(_08776_));
 sky130_fd_sc_hd__a211oi_1 _13834_ (.A1(_08733_),
    .A2(_08722_),
    .B1(_08623_),
    .C1(_08590_),
    .Y(_08787_));
 sky130_fd_sc_hd__a211o_1 _13835_ (.A1(_08733_),
    .A2(_08722_),
    .B1(_08623_),
    .C1(_08590_),
    .X(_08798_));
 sky130_fd_sc_hd__a2bb2oi_1 _13836_ (.A1_N(_08568_),
    .A2_N(_08579_),
    .B1(_08634_),
    .B2(_08744_),
    .Y(_08809_));
 sky130_fd_sc_hd__o21ai_1 _13837_ (.A1(_08568_),
    .A2(_08579_),
    .B1(_08765_),
    .Y(_08820_));
 sky130_fd_sc_hd__o2bb2ai_1 _13838_ (.A1_N(_07329_),
    .A2_N(_07384_),
    .B1(_08590_),
    .B2(_08754_),
    .Y(_08831_));
 sky130_fd_sc_hd__o22ai_2 _13839_ (.A1(_07318_),
    .A2(_07373_),
    .B1(_08787_),
    .B2(_08809_),
    .Y(_08842_));
 sky130_fd_sc_hd__and3_1 _13840_ (.A(_08798_),
    .B(_08820_),
    .C(_08557_),
    .X(_08853_));
 sky130_fd_sc_hd__nand3_1 _13841_ (.A(_08820_),
    .B(_08557_),
    .C(_08798_),
    .Y(_08864_));
 sky130_fd_sc_hd__o221a_2 _13842_ (.A1(_08524_),
    .A2(_08535_),
    .B1(_08776_),
    .B2(_08831_),
    .C1(_08864_),
    .X(_08875_));
 sky130_fd_sc_hd__a21oi_2 _13843_ (.A1(_08842_),
    .A2(_08864_),
    .B1(_08546_),
    .Y(_08886_));
 sky130_fd_sc_hd__a2bb2o_1 _13844_ (.A1_N(_08502_),
    .A2_N(_08513_),
    .B1(_08842_),
    .B2(_08864_),
    .X(_08897_));
 sky130_fd_sc_hd__nand2_1 _13845_ (.A(_07417_),
    .B(_07603_),
    .Y(_08908_));
 sky130_fd_sc_hd__a21boi_2 _13846_ (.A1(_07406_),
    .A2(_07582_),
    .B1_N(_07417_),
    .Y(_08919_));
 sky130_fd_sc_hd__o211a_1 _13847_ (.A1(_08875_),
    .A2(_08886_),
    .B1(_07417_),
    .C1(_07603_),
    .X(_08930_));
 sky130_fd_sc_hd__o21ai_2 _13848_ (.A1(_08875_),
    .A2(_08886_),
    .B1(_08919_),
    .Y(_08941_));
 sky130_fd_sc_hd__nand3b_2 _13849_ (.A_N(_08875_),
    .B(_08908_),
    .C(_08897_),
    .Y(_08952_));
 sky130_fd_sc_hd__o2bb2a_1 _13850_ (.A1_N(net12),
    .A2_N(_07680_),
    .B1(_07669_),
    .B2(_04528_),
    .X(_08963_));
 sky130_fd_sc_hd__a22o_1 _13851_ (.A1(net12),
    .A2(_07680_),
    .B1(_04539_),
    .B2(_07658_),
    .X(_08974_));
 sky130_fd_sc_hd__a32oi_4 _13852_ (.A1(_04419_),
    .A2(_04452_),
    .A3(net292),
    .B1(_06848_),
    .B2(net23),
    .Y(_08985_));
 sky130_fd_sc_hd__nand3_1 _13853_ (.A(net314),
    .B(net267),
    .C(net299),
    .Y(_08996_));
 sky130_fd_sc_hd__nand2_1 _13854_ (.A(net26),
    .B(_05710_),
    .Y(_09007_));
 sky130_fd_sc_hd__a21oi_2 _13855_ (.A1(_08996_),
    .A2(_09007_),
    .B1(_08985_),
    .Y(_09018_));
 sky130_fd_sc_hd__o221a_1 _13856_ (.A1(_04758_),
    .A2(_05699_),
    .B1(net298),
    .B2(_03506_),
    .C1(_08985_),
    .X(_09029_));
 sky130_fd_sc_hd__o221ai_4 _13857_ (.A1(_04758_),
    .A2(_05699_),
    .B1(net298),
    .B2(_03506_),
    .C1(_08985_),
    .Y(_09040_));
 sky130_fd_sc_hd__nand3b_2 _13858_ (.A_N(_09018_),
    .B(_09040_),
    .C(_08963_),
    .Y(_09051_));
 sky130_fd_sc_hd__o21ai_2 _13859_ (.A1(_09018_),
    .A2(_09029_),
    .B1(_08974_),
    .Y(_09062_));
 sky130_fd_sc_hd__a31oi_2 _13860_ (.A1(_07439_),
    .A2(_07450_),
    .A3(_07461_),
    .B1(_07428_),
    .Y(_09073_));
 sky130_fd_sc_hd__o2bb2ai_4 _13861_ (.A1_N(_09051_),
    .A2_N(_09062_),
    .B1(_09073_),
    .B2(_07472_),
    .Y(_09084_));
 sky130_fd_sc_hd__o2111ai_2 _13862_ (.A1(_07428_),
    .A2(_07494_),
    .B1(_09051_),
    .C1(_09062_),
    .D1(_07483_),
    .Y(_09095_));
 sky130_fd_sc_hd__nand2_1 _13863_ (.A(_09084_),
    .B(_09095_),
    .Y(_09106_));
 sky130_fd_sc_hd__o31a_1 _13864_ (.A1(_03176_),
    .A2(_07702_),
    .A3(_07757_),
    .B1(_07779_),
    .X(_09117_));
 sky130_fd_sc_hd__a21oi_1 _13865_ (.A1(_09084_),
    .A2(_09095_),
    .B1(_09117_),
    .Y(_09128_));
 sky130_fd_sc_hd__and3_1 _13866_ (.A(_09084_),
    .B(_09095_),
    .C(_09117_),
    .X(_09139_));
 sky130_fd_sc_hd__o311a_1 _13867_ (.A1(_03176_),
    .A2(_07702_),
    .A3(_07757_),
    .B1(_07779_),
    .C1(_09106_),
    .X(_09150_));
 sky130_fd_sc_hd__nor2_1 _13868_ (.A(_09106_),
    .B(_09117_),
    .Y(_09161_));
 sky130_fd_sc_hd__or2_1 _13869_ (.A(_09106_),
    .B(_09117_),
    .X(_09172_));
 sky130_fd_sc_hd__nor2_1 _13870_ (.A(_09128_),
    .B(_09139_),
    .Y(_09182_));
 sky130_fd_sc_hd__o211ai_1 _13871_ (.A1(_09150_),
    .A2(_09161_),
    .B1(_08941_),
    .C1(_08952_),
    .Y(_09193_));
 sky130_fd_sc_hd__o2bb2ai_1 _13872_ (.A1_N(_08941_),
    .A2_N(_08952_),
    .B1(_09128_),
    .B2(_09139_),
    .Y(_09204_));
 sky130_fd_sc_hd__o2bb2a_1 _13873_ (.A1_N(_08941_),
    .A2_N(_08952_),
    .B1(_09150_),
    .B2(_09161_),
    .X(_09215_));
 sky130_fd_sc_hd__o2bb2ai_1 _13874_ (.A1_N(_08941_),
    .A2_N(_08952_),
    .B1(_09150_),
    .B2(_09161_),
    .Y(_09226_));
 sky130_fd_sc_hd__o211ai_1 _13875_ (.A1(_09128_),
    .A2(_09139_),
    .B1(_08941_),
    .C1(_08952_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_1 _13876_ (.A(_08381_),
    .B(_09237_),
    .Y(_09248_));
 sky130_fd_sc_hd__nand3_1 _13877_ (.A(_08381_),
    .B(_09226_),
    .C(_09237_),
    .Y(_09259_));
 sky130_fd_sc_hd__nand3_2 _13878_ (.A(_09204_),
    .B(_08370_),
    .C(_09193_),
    .Y(_09270_));
 sky130_fd_sc_hd__a21o_1 _13879_ (.A1(_09259_),
    .A2(_09270_),
    .B1(_08359_),
    .X(_09281_));
 sky130_fd_sc_hd__o211ai_2 _13880_ (.A1(_09248_),
    .A2(_09215_),
    .B1(_08359_),
    .C1(_09270_),
    .Y(_09292_));
 sky130_fd_sc_hd__nand4_2 _13881_ (.A(_08327_),
    .B(_08338_),
    .C(_09259_),
    .D(_09270_),
    .Y(_09303_));
 sky130_fd_sc_hd__a22o_1 _13882_ (.A1(_08327_),
    .A2(_08338_),
    .B1(_09259_),
    .B2(_09270_),
    .X(_09314_));
 sky130_fd_sc_hd__nand3_4 _13883_ (.A(_08239_),
    .B(_09281_),
    .C(_09292_),
    .Y(_09325_));
 sky130_fd_sc_hd__a22oi_1 _13884_ (.A1(_08031_),
    .A2(_08217_),
    .B1(_09281_),
    .B2(_09292_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand3_4 _13885_ (.A(_09314_),
    .B(_08228_),
    .C(_09303_),
    .Y(_09347_));
 sky130_fd_sc_hd__nand4_4 _13886_ (.A(_09325_),
    .B(_09347_),
    .C(_07154_),
    .D(_08086_),
    .Y(_09358_));
 sky130_fd_sc_hd__a32o_1 _13887_ (.A1(_07154_),
    .A2(_08042_),
    .A3(_08053_),
    .B1(_09325_),
    .B2(_09347_),
    .X(_09369_));
 sky130_fd_sc_hd__nand3_1 _13888_ (.A(_08097_),
    .B(_09325_),
    .C(_09347_),
    .Y(_09380_));
 sky130_fd_sc_hd__a21o_1 _13889_ (.A1(_09325_),
    .A2(_09347_),
    .B1(_08097_),
    .X(_09391_));
 sky130_fd_sc_hd__nand2_1 _13890_ (.A(_09358_),
    .B(_09369_),
    .Y(_09402_));
 sky130_fd_sc_hd__nand4_1 _13891_ (.A(_08141_),
    .B(_09358_),
    .C(_09369_),
    .D(_07045_),
    .Y(_09413_));
 sky130_fd_sc_hd__o31a_1 _13892_ (.A1(_08875_),
    .A2(_08886_),
    .A3(_08919_),
    .B1(_09182_),
    .X(_09424_));
 sky130_fd_sc_hd__o21ai_1 _13893_ (.A1(_09128_),
    .A2(_09139_),
    .B1(_08941_),
    .Y(_09435_));
 sky130_fd_sc_hd__o31ai_2 _13894_ (.A1(_08875_),
    .A2(_08886_),
    .A3(_08919_),
    .B1(_09435_),
    .Y(_09446_));
 sky130_fd_sc_hd__o22a_1 _13895_ (.A1(_08502_),
    .A2(_08513_),
    .B1(_08776_),
    .B2(_08831_),
    .X(_09457_));
 sky130_fd_sc_hd__a2bb2o_1 _13896_ (.A1_N(_08776_),
    .A2_N(_08831_),
    .B1(_08864_),
    .B2(_08546_),
    .X(_09468_));
 sky130_fd_sc_hd__a32oi_4 _13897_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net28),
    .Y(_09479_));
 sky130_fd_sc_hd__a32o_1 _13898_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net28),
    .X(_09490_));
 sky130_fd_sc_hd__a32oi_4 _13899_ (.A1(_05841_),
    .A2(_05863_),
    .A3(net305),
    .B1(_04911_),
    .B2(net29),
    .Y(_09501_));
 sky130_fd_sc_hd__o211ai_4 _13900_ (.A1(net267),
    .A2(_06508_),
    .B1(net317),
    .C1(_06486_),
    .Y(_09512_));
 sky130_fd_sc_hd__or3b_2 _13901_ (.A(net58),
    .B(_03916_),
    .C_N(net55),
    .X(_09523_));
 sky130_fd_sc_hd__a21oi_4 _13902_ (.A1(_09512_),
    .A2(_09523_),
    .B1(_09501_),
    .Y(_09534_));
 sky130_fd_sc_hd__o221a_1 _13903_ (.A1(_03916_),
    .A2(_04660_),
    .B1(_06552_),
    .B2(_04638_),
    .C1(_09501_),
    .X(_09545_));
 sky130_fd_sc_hd__o211ai_1 _13904_ (.A1(_03916_),
    .A2(_04660_),
    .B1(_09512_),
    .C1(_09501_),
    .Y(_09556_));
 sky130_fd_sc_hd__a31oi_2 _13905_ (.A1(_09501_),
    .A2(_09512_),
    .A3(_09523_),
    .B1(_09479_),
    .Y(_09567_));
 sky130_fd_sc_hd__a31o_1 _13906_ (.A1(_09501_),
    .A2(_09512_),
    .A3(_09523_),
    .B1(_09479_),
    .X(_09578_));
 sky130_fd_sc_hd__nor2_1 _13907_ (.A(_09534_),
    .B(_09578_),
    .Y(_09588_));
 sky130_fd_sc_hd__o21a_1 _13908_ (.A1(_09534_),
    .A2(_09545_),
    .B1(_09479_),
    .X(_09599_));
 sky130_fd_sc_hd__o21ai_2 _13909_ (.A1(_09534_),
    .A2(_09545_),
    .B1(_09479_),
    .Y(_09610_));
 sky130_fd_sc_hd__o21ai_1 _13910_ (.A1(_09534_),
    .A2(_09578_),
    .B1(_09610_),
    .Y(_09621_));
 sky130_fd_sc_hd__o21ai_4 _13911_ (.A1(_08590_),
    .A2(_08623_),
    .B1(_08744_),
    .Y(_09632_));
 sky130_fd_sc_hd__a32o_2 _13912_ (.A1(_07242_),
    .A2(net258),
    .A3(_04342_),
    .B1(_04364_),
    .B2(net31),
    .X(_09643_));
 sky130_fd_sc_hd__nor3_4 _13913_ (.A(net31),
    .B(net32),
    .C(net2),
    .Y(_09654_));
 sky130_fd_sc_hd__or3_4 _13914_ (.A(net31),
    .B(net32),
    .C(net2),
    .X(_09665_));
 sky130_fd_sc_hd__nand4_4 _13915_ (.A(net312),
    .B(net297),
    .C(_09654_),
    .D(_03916_),
    .Y(_09676_));
 sky130_fd_sc_hd__a41oi_4 _13916_ (.A1(net308),
    .A2(net297),
    .A3(_08645_),
    .A4(_03916_),
    .B1(_03960_),
    .Y(_09687_));
 sky130_fd_sc_hd__a41o_4 _13917_ (.A1(net309),
    .A2(net297),
    .A3(_08645_),
    .A4(_03916_),
    .B1(_03960_),
    .X(_09698_));
 sky130_fd_sc_hd__a21oi_4 _13918_ (.A1(_06519_),
    .A2(net290),
    .B1(_09687_),
    .Y(_09709_));
 sky130_fd_sc_hd__o21ai_4 _13919_ (.A1(net260),
    .A2(_09665_),
    .B1(_09698_),
    .Y(_09720_));
 sky130_fd_sc_hd__o211ai_2 _13920_ (.A1(_06530_),
    .A2(_09665_),
    .B1(net33),
    .C1(_09698_),
    .Y(_09731_));
 sky130_fd_sc_hd__nor2_2 _13921_ (.A(_03949_),
    .B(_04331_),
    .Y(_09742_));
 sky130_fd_sc_hd__or3_1 _13922_ (.A(net44),
    .B(_03949_),
    .C(_03286_),
    .X(_09753_));
 sky130_fd_sc_hd__o211ai_2 _13923_ (.A1(_06530_),
    .A2(_08656_),
    .B1(_04484_),
    .C1(_08700_),
    .Y(_09764_));
 sky130_fd_sc_hd__o211ai_4 _13924_ (.A1(_03949_),
    .A2(_04331_),
    .B1(_09731_),
    .C1(_09764_),
    .Y(_09775_));
 sky130_fd_sc_hd__nand4_4 _13925_ (.A(net255),
    .B(_09698_),
    .C(_09742_),
    .D(net33),
    .Y(_09786_));
 sky130_fd_sc_hd__o31a_1 _13926_ (.A1(_03286_),
    .A2(_09720_),
    .A3(_09753_),
    .B1(_09643_),
    .X(_09797_));
 sky130_fd_sc_hd__o311a_1 _13927_ (.A1(_03286_),
    .A2(_09720_),
    .A3(_09753_),
    .B1(_09775_),
    .C1(_09643_),
    .X(_09808_));
 sky130_fd_sc_hd__nand3_2 _13928_ (.A(_09643_),
    .B(_09775_),
    .C(_09786_),
    .Y(_09819_));
 sky130_fd_sc_hd__a21oi_2 _13929_ (.A1(_09775_),
    .A2(_09786_),
    .B1(_09643_),
    .Y(_09830_));
 sky130_fd_sc_hd__a21o_1 _13930_ (.A1(_09775_),
    .A2(_09786_),
    .B1(_09643_),
    .X(_09841_));
 sky130_fd_sc_hd__nand2_1 _13931_ (.A(_09819_),
    .B(_09841_),
    .Y(_09852_));
 sky130_fd_sc_hd__a211oi_4 _13932_ (.A1(_09797_),
    .A2(_09775_),
    .B1(_09632_),
    .C1(_09830_),
    .Y(_09863_));
 sky130_fd_sc_hd__o2111ai_4 _13933_ (.A1(_08590_),
    .A2(_08623_),
    .B1(_08744_),
    .C1(_09819_),
    .D1(_09841_),
    .Y(_09874_));
 sky130_fd_sc_hd__a21boi_2 _13934_ (.A1(_09819_),
    .A2(_09841_),
    .B1_N(_09632_),
    .Y(_09885_));
 sky130_fd_sc_hd__o21ai_2 _13935_ (.A1(_09808_),
    .A2(_09830_),
    .B1(_09632_),
    .Y(_09896_));
 sky130_fd_sc_hd__o211ai_2 _13936_ (.A1(_09588_),
    .A2(_09599_),
    .B1(_09874_),
    .C1(_09896_),
    .Y(_09907_));
 sky130_fd_sc_hd__o21bai_2 _13937_ (.A1(_09863_),
    .A2(_09885_),
    .B1_N(_09621_),
    .Y(_09918_));
 sky130_fd_sc_hd__a21oi_1 _13938_ (.A1(_09852_),
    .A2(_09632_),
    .B1(_09621_),
    .Y(_09929_));
 sky130_fd_sc_hd__o2111ai_4 _13939_ (.A1(_09534_),
    .A2(_09578_),
    .B1(_09610_),
    .C1(_09874_),
    .D1(_09896_),
    .Y(_09940_));
 sky130_fd_sc_hd__o21ai_1 _13940_ (.A1(_09863_),
    .A2(_09885_),
    .B1(_09621_),
    .Y(_09951_));
 sky130_fd_sc_hd__nand3_4 _13941_ (.A(_09951_),
    .B(_09468_),
    .C(_09940_),
    .Y(_09962_));
 sky130_fd_sc_hd__o211a_1 _13942_ (.A1(_08853_),
    .A2(_09457_),
    .B1(_09907_),
    .C1(_09918_),
    .X(_09973_));
 sky130_fd_sc_hd__o211ai_4 _13943_ (.A1(_08853_),
    .A2(_09457_),
    .B1(_09907_),
    .C1(_09918_),
    .Y(_09984_));
 sky130_fd_sc_hd__a21oi_1 _13944_ (.A1(_08425_),
    .A2(_08458_),
    .B1(_08392_),
    .Y(_09995_));
 sky130_fd_sc_hd__a21boi_1 _13945_ (.A1(_08392_),
    .A2(_08491_),
    .B1_N(_08469_),
    .Y(_10006_));
 sky130_fd_sc_hd__a32o_1 _13946_ (.A1(_07658_),
    .A2(_04452_),
    .A3(_04419_),
    .B1(net23),
    .B2(_07680_),
    .X(_10017_));
 sky130_fd_sc_hd__or3b_1 _13947_ (.A(_03616_),
    .B(net61),
    .C_N(net60),
    .X(_10027_));
 sky130_fd_sc_hd__nand3_2 _13948_ (.A(_04998_),
    .B(_05009_),
    .C(net299),
    .Y(_10038_));
 sky130_fd_sc_hd__a32oi_4 _13949_ (.A1(net314),
    .A2(net267),
    .A3(net292),
    .B1(_06848_),
    .B2(net26),
    .Y(_10049_));
 sky130_fd_sc_hd__o211a_1 _13950_ (.A1(_03616_),
    .A2(net298),
    .B1(_10038_),
    .C1(_10049_),
    .X(_10060_));
 sky130_fd_sc_hd__o211ai_2 _13951_ (.A1(_03616_),
    .A2(net298),
    .B1(_10038_),
    .C1(_10049_),
    .Y(_10071_));
 sky130_fd_sc_hd__a21oi_1 _13952_ (.A1(_10027_),
    .A2(_10038_),
    .B1(_10049_),
    .Y(_10082_));
 sky130_fd_sc_hd__a21o_1 _13953_ (.A1(_10027_),
    .A2(_10038_),
    .B1(_10049_),
    .X(_10093_));
 sky130_fd_sc_hd__a221o_1 _13954_ (.A1(_04463_),
    .A2(_07658_),
    .B1(_07680_),
    .B2(net23),
    .C1(_10082_),
    .X(_10104_));
 sky130_fd_sc_hd__a21o_1 _13955_ (.A1(_10017_),
    .A2(_10071_),
    .B1(_10082_),
    .X(_10115_));
 sky130_fd_sc_hd__nand3b_1 _13956_ (.A_N(_10017_),
    .B(_10071_),
    .C(_10093_),
    .Y(_10126_));
 sky130_fd_sc_hd__o21ai_1 _13957_ (.A1(_10060_),
    .A2(_10082_),
    .B1(_10017_),
    .Y(_10137_));
 sky130_fd_sc_hd__o211a_1 _13958_ (.A1(_08480_),
    .A2(_09995_),
    .B1(_10126_),
    .C1(_10137_),
    .X(_10148_));
 sky130_fd_sc_hd__a21oi_2 _13959_ (.A1(_10126_),
    .A2(_10137_),
    .B1(_10006_),
    .Y(_10159_));
 sky130_fd_sc_hd__a21oi_1 _13960_ (.A1(_08974_),
    .A2(_09040_),
    .B1(_09018_),
    .Y(_10170_));
 sky130_fd_sc_hd__nor3_1 _13961_ (.A(_10148_),
    .B(_10170_),
    .C(_10159_),
    .Y(_10181_));
 sky130_fd_sc_hd__o21a_1 _13962_ (.A1(_10148_),
    .A2(_10159_),
    .B1(_10170_),
    .X(_10192_));
 sky130_fd_sc_hd__o21ba_1 _13963_ (.A1(_10148_),
    .A2(_10159_),
    .B1_N(_10170_),
    .X(_10203_));
 sky130_fd_sc_hd__a2111oi_2 _13964_ (.A1(_08974_),
    .A2(_09040_),
    .B1(_10148_),
    .C1(_10159_),
    .D1(_09018_),
    .Y(_10214_));
 sky130_fd_sc_hd__nor2_1 _13965_ (.A(_10203_),
    .B(_10214_),
    .Y(_10225_));
 sky130_fd_sc_hd__o211ai_2 _13966_ (.A1(_10181_),
    .A2(_10192_),
    .B1(_09962_),
    .C1(_09984_),
    .Y(_10236_));
 sky130_fd_sc_hd__o2bb2ai_2 _13967_ (.A1_N(_09962_),
    .A2_N(_09984_),
    .B1(_10203_),
    .B2(_10214_),
    .Y(_10247_));
 sky130_fd_sc_hd__o2bb2ai_1 _13968_ (.A1_N(_09962_),
    .A2_N(_09984_),
    .B1(_10181_),
    .B2(_10192_),
    .Y(_10258_));
 sky130_fd_sc_hd__o211ai_2 _13969_ (.A1(_10203_),
    .A2(_10214_),
    .B1(_09962_),
    .C1(_09984_),
    .Y(_10269_));
 sky130_fd_sc_hd__o211a_1 _13970_ (.A1(_08930_),
    .A2(_09424_),
    .B1(_10236_),
    .C1(_10247_),
    .X(_10280_));
 sky130_fd_sc_hd__o211ai_4 _13971_ (.A1(_08930_),
    .A2(_09424_),
    .B1(_10236_),
    .C1(_10247_),
    .Y(_10291_));
 sky130_fd_sc_hd__nand3_4 _13972_ (.A(_09446_),
    .B(_10258_),
    .C(_10269_),
    .Y(_10302_));
 sky130_fd_sc_hd__and2b_4 _13973_ (.A_N(net64),
    .B(net34),
    .X(_10313_));
 sky130_fd_sc_hd__nand2b_4 _13974_ (.A_N(net64),
    .B(net34),
    .Y(_10324_));
 sky130_fd_sc_hd__and2b_4 _13975_ (.A_N(net34),
    .B(net64),
    .X(_10335_));
 sky130_fd_sc_hd__nand2_8 _13976_ (.A(_03971_),
    .B(net64),
    .Y(_10346_));
 sky130_fd_sc_hd__a21oi_1 _13977_ (.A1(_10324_),
    .A2(_10346_),
    .B1(_03176_),
    .Y(_10357_));
 sky130_fd_sc_hd__a22o_1 _13978_ (.A1(net12),
    .A2(_08272_),
    .B1(_04539_),
    .B2(_08250_),
    .X(_10368_));
 sky130_fd_sc_hd__o211a_4 _13979_ (.A1(_10313_),
    .A2(_10335_),
    .B1(net1),
    .C1(_10368_),
    .X(_10379_));
 sky130_fd_sc_hd__nor2_1 _13980_ (.A(_10357_),
    .B(_10368_),
    .Y(_10390_));
 sky130_fd_sc_hd__or2_2 _13981_ (.A(_10379_),
    .B(_10390_),
    .X(_10401_));
 sky130_fd_sc_hd__o21a_1 _13982_ (.A1(_09106_),
    .A2(_09117_),
    .B1(_09084_),
    .X(_10411_));
 sky130_fd_sc_hd__a21oi_4 _13983_ (.A1(_09084_),
    .A2(_09172_),
    .B1(_10401_),
    .Y(_10422_));
 sky130_fd_sc_hd__o221a_1 _13984_ (.A1(_10379_),
    .A2(_10390_),
    .B1(_09106_),
    .B2(_09117_),
    .C1(_09084_),
    .X(_10433_));
 sky130_fd_sc_hd__and3b_1 _13985_ (.A_N(_10401_),
    .B(_09172_),
    .C(_09084_),
    .X(_10444_));
 sky130_fd_sc_hd__o2bb2a_1 _13986_ (.A1_N(_09084_),
    .A2_N(_09172_),
    .B1(_10379_),
    .B2(_10390_),
    .X(_10455_));
 sky130_fd_sc_hd__nor2_1 _13987_ (.A(_10444_),
    .B(_10455_),
    .Y(_10466_));
 sky130_fd_sc_hd__o211ai_1 _13988_ (.A1(_10422_),
    .A2(_10433_),
    .B1(_10291_),
    .C1(_10302_),
    .Y(_10477_));
 sky130_fd_sc_hd__o2bb2ai_1 _13989_ (.A1_N(_10291_),
    .A2_N(_10302_),
    .B1(_10444_),
    .B2(_10455_),
    .Y(_10488_));
 sky130_fd_sc_hd__o2bb2ai_1 _13990_ (.A1_N(_10291_),
    .A2_N(_10302_),
    .B1(_10422_),
    .B2(_10433_),
    .Y(_10499_));
 sky130_fd_sc_hd__o211ai_2 _13991_ (.A1(_10444_),
    .A2(_10455_),
    .B1(_10291_),
    .C1(_10302_),
    .Y(_10510_));
 sky130_fd_sc_hd__o2bb2ai_1 _13992_ (.A1_N(_08349_),
    .A2_N(_09270_),
    .B1(_09248_),
    .B2(_09215_),
    .Y(_10521_));
 sky130_fd_sc_hd__a2bb2oi_1 _13993_ (.A1_N(_09215_),
    .A2_N(_09248_),
    .B1(_09270_),
    .B2(_08349_),
    .Y(_10532_));
 sky130_fd_sc_hd__nand3_2 _13994_ (.A(_10477_),
    .B(_10488_),
    .C(_10532_),
    .Y(_10543_));
 sky130_fd_sc_hd__nand3_2 _13995_ (.A(_10499_),
    .B(_10510_),
    .C(_10521_),
    .Y(_10554_));
 sky130_fd_sc_hd__a21oi_1 _13996_ (.A1(_10543_),
    .A2(_10554_),
    .B1(_08316_),
    .Y(_10565_));
 sky130_fd_sc_hd__a21o_1 _13997_ (.A1(_10543_),
    .A2(_10554_),
    .B1(_08316_),
    .X(_10576_));
 sky130_fd_sc_hd__o2111a_1 _13998_ (.A1(_07856_),
    .A2(_08305_),
    .B1(_08294_),
    .C1(_10554_),
    .D1(_10543_),
    .X(_10587_));
 sky130_fd_sc_hd__o2111ai_4 _13999_ (.A1(_07856_),
    .A2(_08305_),
    .B1(_08294_),
    .C1(_10554_),
    .D1(_10543_),
    .Y(_10598_));
 sky130_fd_sc_hd__nand2_1 _14000_ (.A(_10576_),
    .B(_10598_),
    .Y(_10609_));
 sky130_fd_sc_hd__a31o_1 _14001_ (.A1(_09325_),
    .A2(_08086_),
    .A3(_07154_),
    .B1(_09336_),
    .X(_10620_));
 sky130_fd_sc_hd__o211ai_2 _14002_ (.A1(_10565_),
    .A2(_10587_),
    .B1(_09347_),
    .C1(_09358_),
    .Y(_10631_));
 sky130_fd_sc_hd__and3_1 _14003_ (.A(_10576_),
    .B(_10598_),
    .C(_09336_),
    .X(_10642_));
 sky130_fd_sc_hd__nor2_1 _14004_ (.A(_09358_),
    .B(_10609_),
    .Y(_10653_));
 sky130_fd_sc_hd__nand3_2 _14005_ (.A(_10576_),
    .B(_10598_),
    .C(_10620_),
    .Y(_10664_));
 sky130_fd_sc_hd__nand4_1 _14006_ (.A(_09347_),
    .B(_09358_),
    .C(_10576_),
    .D(_10598_),
    .Y(_10675_));
 sky130_fd_sc_hd__o21ai_1 _14007_ (.A1(_10565_),
    .A2(_10587_),
    .B1(_10620_),
    .Y(_10686_));
 sky130_fd_sc_hd__and4_1 _14008_ (.A(_07078_),
    .B(_08119_),
    .C(_09325_),
    .D(_09347_),
    .X(_10697_));
 sky130_fd_sc_hd__and4_1 _14009_ (.A(_07078_),
    .B(_08119_),
    .C(_09325_),
    .D(_09347_),
    .X(_10708_));
 sky130_fd_sc_hd__o2111ai_4 _14010_ (.A1(_07154_),
    .A2(_08086_),
    .B1(_09325_),
    .C1(_09347_),
    .D1(_07078_),
    .Y(_10719_));
 sky130_fd_sc_hd__nand3_1 _14011_ (.A(_10675_),
    .B(_10686_),
    .C(_10719_),
    .Y(_10730_));
 sky130_fd_sc_hd__and3_1 _14012_ (.A(_10631_),
    .B(_10664_),
    .C(_10708_),
    .X(_10741_));
 sky130_fd_sc_hd__nand3_1 _14013_ (.A(_10631_),
    .B(_10664_),
    .C(_10708_),
    .Y(_10752_));
 sky130_fd_sc_hd__a31oi_1 _14014_ (.A1(_10675_),
    .A2(_10686_),
    .A3(_10719_),
    .B1(_09413_),
    .Y(_10763_));
 sky130_fd_sc_hd__o2bb2ai_1 _14015_ (.A1_N(_10730_),
    .A2_N(_10752_),
    .B1(_08163_),
    .B2(_09402_),
    .Y(_10774_));
 sky130_fd_sc_hd__nand2b_1 _14016_ (.A_N(_10763_),
    .B(_10774_),
    .Y(_10785_));
 sky130_fd_sc_hd__o211ai_1 _14017_ (.A1(_07067_),
    .A2(_08108_),
    .B1(_09380_),
    .C1(_09391_),
    .Y(_10796_));
 sky130_fd_sc_hd__nand2_1 _14018_ (.A(_10719_),
    .B(_10796_),
    .Y(_10807_));
 sky130_fd_sc_hd__nor2_1 _14019_ (.A(_08185_),
    .B(_10807_),
    .Y(_10817_));
 sky130_fd_sc_hd__or3_1 _14020_ (.A(_07133_),
    .B(_08174_),
    .C(_10807_),
    .X(_10828_));
 sky130_fd_sc_hd__xnor2_1 _14021_ (.A(_10785_),
    .B(_10817_),
    .Y(net66));
 sky130_fd_sc_hd__o21ai_2 _14022_ (.A1(_10763_),
    .A2(_10817_),
    .B1(_10774_),
    .Y(_10849_));
 sky130_fd_sc_hd__a32o_2 _14023_ (.A1(_10499_),
    .A2(_10510_),
    .A3(_10521_),
    .B1(_10543_),
    .B2(_08316_),
    .X(_10860_));
 sky130_fd_sc_hd__inv_2 _14024_ (.A(_10860_),
    .Y(_10871_));
 sky130_fd_sc_hd__o21a_1 _14025_ (.A1(_10181_),
    .A2(_10192_),
    .B1(_09962_),
    .X(_10882_));
 sky130_fd_sc_hd__a21oi_1 _14026_ (.A1(_09962_),
    .A2(_10225_),
    .B1(_09973_),
    .Y(_10893_));
 sky130_fd_sc_hd__a32o_1 _14027_ (.A1(_07658_),
    .A2(net267),
    .A3(net314),
    .B1(net26),
    .B2(_07680_),
    .X(_10904_));
 sky130_fd_sc_hd__a32oi_4 _14028_ (.A1(_04998_),
    .A2(_05009_),
    .A3(net292),
    .B1(_06848_),
    .B2(net27),
    .Y(_10915_));
 sky130_fd_sc_hd__or3b_1 _14029_ (.A(_03725_),
    .B(net61),
    .C_N(net60),
    .X(_10926_));
 sky130_fd_sc_hd__o211ai_2 _14030_ (.A1(net267),
    .A2(_05436_),
    .B1(net299),
    .C1(_05414_),
    .Y(_10937_));
 sky130_fd_sc_hd__a21oi_1 _14031_ (.A1(_10926_),
    .A2(_10937_),
    .B1(_10915_),
    .Y(_10948_));
 sky130_fd_sc_hd__a21o_1 _14032_ (.A1(_10926_),
    .A2(_10937_),
    .B1(_10915_),
    .X(_10959_));
 sky130_fd_sc_hd__o211a_1 _14033_ (.A1(_03725_),
    .A2(net298),
    .B1(_10937_),
    .C1(_10915_),
    .X(_10970_));
 sky130_fd_sc_hd__o221ai_4 _14034_ (.A1(_05457_),
    .A2(_05699_),
    .B1(net298),
    .B2(_03725_),
    .C1(_10915_),
    .Y(_10981_));
 sky130_fd_sc_hd__nand3_2 _14035_ (.A(_10904_),
    .B(_10959_),
    .C(_10981_),
    .Y(_10992_));
 sky130_fd_sc_hd__o21bai_1 _14036_ (.A1(_10948_),
    .A2(_10970_),
    .B1_N(_10904_),
    .Y(_11003_));
 sky130_fd_sc_hd__o21ai_1 _14037_ (.A1(_10948_),
    .A2(_10970_),
    .B1(_10904_),
    .Y(_11014_));
 sky130_fd_sc_hd__nand3b_1 _14038_ (.A_N(_10904_),
    .B(_10959_),
    .C(_10981_),
    .Y(_11025_));
 sky130_fd_sc_hd__a21oi_1 _14039_ (.A1(_09490_),
    .A2(_09556_),
    .B1(_09534_),
    .Y(_11036_));
 sky130_fd_sc_hd__nand3_1 _14040_ (.A(_11014_),
    .B(_11036_),
    .C(_11025_),
    .Y(_11047_));
 sky130_fd_sc_hd__o211ai_4 _14041_ (.A1(_09534_),
    .A2(_09567_),
    .B1(_10992_),
    .C1(_11003_),
    .Y(_11058_));
 sky130_fd_sc_hd__a21oi_1 _14042_ (.A1(_11047_),
    .A2(_11058_),
    .B1(_10115_),
    .Y(_11069_));
 sky130_fd_sc_hd__and3_1 _14043_ (.A(_11047_),
    .B(_11058_),
    .C(_10115_),
    .X(_11080_));
 sky130_fd_sc_hd__nand4_1 _14044_ (.A(_10071_),
    .B(_10104_),
    .C(_11047_),
    .D(_11058_),
    .Y(_11091_));
 sky130_fd_sc_hd__nand2b_1 _14045_ (.A_N(_11069_),
    .B(_11091_),
    .Y(_11102_));
 sky130_fd_sc_hd__and3_1 _14046_ (.A(_05841_),
    .B(_05863_),
    .C(_05227_),
    .X(_11113_));
 sky130_fd_sc_hd__nor2_1 _14047_ (.A(_03835_),
    .B(_05260_),
    .Y(_11124_));
 sky130_fd_sc_hd__a31o_1 _14048_ (.A1(_05841_),
    .A2(_05863_),
    .A3(_05227_),
    .B1(_11124_),
    .X(_11135_));
 sky130_fd_sc_hd__or3b_1 _14049_ (.A(net59),
    .B(_03916_),
    .C_N(net58),
    .X(_11146_));
 sky130_fd_sc_hd__o211ai_1 _14050_ (.A1(net267),
    .A2(_06508_),
    .B1(net305),
    .C1(_06486_),
    .Y(_11157_));
 sky130_fd_sc_hd__a22oi_4 _14051_ (.A1(net30),
    .A2(_04911_),
    .B1(_06541_),
    .B2(net305),
    .Y(_11168_));
 sky130_fd_sc_hd__or3b_1 _14052_ (.A(net58),
    .B(_03938_),
    .C_N(net55),
    .X(_11179_));
 sky130_fd_sc_hd__nand3_1 _14053_ (.A(_07242_),
    .B(net258),
    .C(net317),
    .Y(_11190_));
 sky130_fd_sc_hd__o221ai_4 _14054_ (.A1(_03938_),
    .A2(_04660_),
    .B1(_07263_),
    .B2(_04638_),
    .C1(_11168_),
    .Y(_11201_));
 sky130_fd_sc_hd__a21oi_2 _14055_ (.A1(_11179_),
    .A2(_11190_),
    .B1(_11168_),
    .Y(_11212_));
 sky130_fd_sc_hd__a22o_1 _14056_ (.A1(_11146_),
    .A2(_11157_),
    .B1(_11179_),
    .B2(_11190_),
    .X(_11223_));
 sky130_fd_sc_hd__a21oi_2 _14057_ (.A1(_11201_),
    .A2(_11223_),
    .B1(_11135_),
    .Y(_11233_));
 sky130_fd_sc_hd__a21o_1 _14058_ (.A1(_11201_),
    .A2(_11223_),
    .B1(_11135_),
    .X(_11244_));
 sky130_fd_sc_hd__o211a_2 _14059_ (.A1(_11113_),
    .A2(_11124_),
    .B1(_11201_),
    .C1(_11223_),
    .X(_11255_));
 sky130_fd_sc_hd__o211ai_2 _14060_ (.A1(_11113_),
    .A2(_11124_),
    .B1(_11201_),
    .C1(_11223_),
    .Y(_11266_));
 sky130_fd_sc_hd__nand2_1 _14061_ (.A(_11244_),
    .B(_11266_),
    .Y(_11277_));
 sky130_fd_sc_hd__a32oi_4 _14062_ (.A1(net33),
    .A2(_09709_),
    .A3(_09742_),
    .B1(_09775_),
    .B2(_09643_),
    .Y(_11288_));
 sky130_fd_sc_hd__o32a_2 _14063_ (.A1(_08689_),
    .A2(_04353_),
    .A3(_08667_),
    .B1(_04375_),
    .B2(_03949_),
    .X(_11299_));
 sky130_fd_sc_hd__a32o_1 _14064_ (.A1(_08700_),
    .A2(_04342_),
    .A3(net256),
    .B1(_04364_),
    .B2(net32),
    .X(_11310_));
 sky130_fd_sc_hd__o211ai_2 _14065_ (.A1(_06530_),
    .A2(_09665_),
    .B1(_04484_),
    .C1(_09698_),
    .Y(_11321_));
 sky130_fd_sc_hd__or3_4 _14066_ (.A(net44),
    .B(_03960_),
    .C(_03286_),
    .X(_11332_));
 sky130_fd_sc_hd__a31oi_4 _14067_ (.A1(net312),
    .A2(net296),
    .A3(_09654_),
    .B1(_03982_),
    .Y(_11343_));
 sky130_fd_sc_hd__a41o_4 _14068_ (.A1(net309),
    .A2(net297),
    .A3(_09654_),
    .A4(_03916_),
    .B1(_03982_),
    .X(_11354_));
 sky130_fd_sc_hd__nor2_2 _14069_ (.A(net2),
    .B(net3),
    .Y(_11365_));
 sky130_fd_sc_hd__nor4_4 _14070_ (.A(net31),
    .B(net32),
    .C(net2),
    .D(net3),
    .Y(_11376_));
 sky130_fd_sc_hd__nand2_8 _14071_ (.A(_08645_),
    .B(_11365_),
    .Y(_11387_));
 sky130_fd_sc_hd__and4_1 _14072_ (.A(net297),
    .B(_08645_),
    .C(_11365_),
    .D(_03916_),
    .X(_11398_));
 sky130_fd_sc_hd__nand4_4 _14073_ (.A(net297),
    .B(_08645_),
    .C(_11365_),
    .D(_03916_),
    .Y(_11409_));
 sky130_fd_sc_hd__nor2_8 _14074_ (.A(net267),
    .B(_11409_),
    .Y(_11420_));
 sky130_fd_sc_hd__nand4_4 _14075_ (.A(net311),
    .B(net296),
    .C(_09654_),
    .D(_03982_),
    .Y(_11431_));
 sky130_fd_sc_hd__a32oi_4 _14076_ (.A1(net312),
    .A2(net296),
    .A3(_11376_),
    .B1(_09676_),
    .B2(net3),
    .Y(_11442_));
 sky130_fd_sc_hd__o2bb2ai_4 _14077_ (.A1_N(net3),
    .A2_N(net255),
    .B1(_11387_),
    .B2(net260),
    .Y(_11453_));
 sky130_fd_sc_hd__o211ai_2 _14078_ (.A1(_06530_),
    .A2(_11387_),
    .B1(net33),
    .C1(_11354_),
    .Y(_11464_));
 sky130_fd_sc_hd__o211ai_4 _14079_ (.A1(_03960_),
    .A2(_04331_),
    .B1(_11321_),
    .C1(_11464_),
    .Y(_11475_));
 sky130_fd_sc_hd__a221o_1 _14080_ (.A1(net255),
    .A2(net3),
    .B1(_06519_),
    .B2(_11376_),
    .C1(_11332_),
    .X(_11486_));
 sky130_fd_sc_hd__a21o_2 _14081_ (.A1(_11475_),
    .A2(_11486_),
    .B1(_11299_),
    .X(_11497_));
 sky130_fd_sc_hd__o211ai_4 _14082_ (.A1(_11332_),
    .A2(net236),
    .B1(_11475_),
    .C1(_11299_),
    .Y(_11508_));
 sky130_fd_sc_hd__a21o_1 _14083_ (.A1(_11475_),
    .A2(_11486_),
    .B1(_11310_),
    .X(_11519_));
 sky130_fd_sc_hd__o211ai_2 _14084_ (.A1(_11332_),
    .A2(net236),
    .B1(_11475_),
    .C1(_11310_),
    .Y(_11530_));
 sky130_fd_sc_hd__a21boi_2 _14085_ (.A1(_11519_),
    .A2(_11530_),
    .B1_N(_11288_),
    .Y(_11541_));
 sky130_fd_sc_hd__nand4_2 _14086_ (.A(_09786_),
    .B(_09819_),
    .C(_11497_),
    .D(_11508_),
    .Y(_11552_));
 sky130_fd_sc_hd__a21oi_4 _14087_ (.A1(_11497_),
    .A2(_11508_),
    .B1(_11288_),
    .Y(_11563_));
 sky130_fd_sc_hd__nand3b_2 _14088_ (.A_N(_11288_),
    .B(_11519_),
    .C(_11530_),
    .Y(_11574_));
 sky130_fd_sc_hd__nand4_4 _14089_ (.A(_11244_),
    .B(_11266_),
    .C(_11552_),
    .D(_11574_),
    .Y(_11585_));
 sky130_fd_sc_hd__o22ai_4 _14090_ (.A1(_11233_),
    .A2(_11255_),
    .B1(_11541_),
    .B2(_11563_),
    .Y(_11596_));
 sky130_fd_sc_hd__nand2_1 _14091_ (.A(_11585_),
    .B(_11596_),
    .Y(_11606_));
 sky130_fd_sc_hd__o21ai_1 _14092_ (.A1(_09621_),
    .A2(_09885_),
    .B1(_09874_),
    .Y(_11617_));
 sky130_fd_sc_hd__o31a_1 _14093_ (.A1(_09588_),
    .A2(_09599_),
    .A3(_09885_),
    .B1(_09874_),
    .X(_11628_));
 sky130_fd_sc_hd__o211a_2 _14094_ (.A1(_09863_),
    .A2(_09929_),
    .B1(_11585_),
    .C1(_11596_),
    .X(_11639_));
 sky130_fd_sc_hd__o211ai_2 _14095_ (.A1(_09863_),
    .A2(_09929_),
    .B1(_11585_),
    .C1(_11596_),
    .Y(_11650_));
 sky130_fd_sc_hd__a21oi_2 _14096_ (.A1(_11585_),
    .A2(_11596_),
    .B1(_11617_),
    .Y(_11661_));
 sky130_fd_sc_hd__a21o_1 _14097_ (.A1(_11585_),
    .A2(_11596_),
    .B1(_11617_),
    .X(_11672_));
 sky130_fd_sc_hd__o211ai_2 _14098_ (.A1(_11069_),
    .A2(_11080_),
    .B1(_11650_),
    .C1(_11672_),
    .Y(_11683_));
 sky130_fd_sc_hd__o21bai_1 _14099_ (.A1(_11639_),
    .A2(_11661_),
    .B1_N(_11102_),
    .Y(_11694_));
 sky130_fd_sc_hd__a21oi_2 _14100_ (.A1(_11606_),
    .A2(_11628_),
    .B1(_11102_),
    .Y(_11705_));
 sky130_fd_sc_hd__nand3b_1 _14101_ (.A_N(_11102_),
    .B(_11650_),
    .C(_11672_),
    .Y(_11716_));
 sky130_fd_sc_hd__o22ai_2 _14102_ (.A1(_11069_),
    .A2(_11080_),
    .B1(_11639_),
    .B2(_11661_),
    .Y(_11727_));
 sky130_fd_sc_hd__o211a_1 _14103_ (.A1(_09973_),
    .A2(_10882_),
    .B1(_11683_),
    .C1(_11694_),
    .X(_11738_));
 sky130_fd_sc_hd__o211ai_2 _14104_ (.A1(_09973_),
    .A2(_10882_),
    .B1(_11683_),
    .C1(_11694_),
    .Y(_11749_));
 sky130_fd_sc_hd__nand3_4 _14105_ (.A(_10893_),
    .B(_11716_),
    .C(_11727_),
    .Y(_11760_));
 sky130_fd_sc_hd__nor2_4 _14106_ (.A(net34),
    .B(_03993_),
    .Y(_11771_));
 sky130_fd_sc_hd__nand2_8 _14107_ (.A(_03971_),
    .B(net35),
    .Y(_11782_));
 sky130_fd_sc_hd__nor2_8 _14108_ (.A(net35),
    .B(_03971_),
    .Y(_11793_));
 sky130_fd_sc_hd__nand2_8 _14109_ (.A(_03993_),
    .B(net34),
    .Y(_11804_));
 sky130_fd_sc_hd__a21oi_4 _14110_ (.A1(_11782_),
    .A2(_11804_),
    .B1(_03176_),
    .Y(_11815_));
 sky130_fd_sc_hd__o21ai_1 _14111_ (.A1(_04298_),
    .A2(_04506_),
    .B1(_10313_),
    .Y(_11826_));
 sky130_fd_sc_hd__nand2_1 _14112_ (.A(net12),
    .B(_10335_),
    .Y(_11837_));
 sky130_fd_sc_hd__nand3_1 _14113_ (.A(_04419_),
    .B(_04452_),
    .C(_08250_),
    .Y(_11848_));
 sky130_fd_sc_hd__nand2_1 _14114_ (.A(net23),
    .B(_08272_),
    .Y(_11859_));
 sky130_fd_sc_hd__a22oi_1 _14115_ (.A1(_11826_),
    .A2(_11837_),
    .B1(_11848_),
    .B2(_11859_),
    .Y(_11870_));
 sky130_fd_sc_hd__a22o_1 _14116_ (.A1(_11826_),
    .A2(_11837_),
    .B1(_11848_),
    .B2(_11859_),
    .X(_11881_));
 sky130_fd_sc_hd__nand4_2 _14117_ (.A(_11826_),
    .B(_11837_),
    .C(_11848_),
    .D(_11859_),
    .Y(_11892_));
 sky130_fd_sc_hd__nand2_2 _14118_ (.A(_11881_),
    .B(_11892_),
    .Y(_11903_));
 sky130_fd_sc_hd__xnor2_4 _14119_ (.A(_11815_),
    .B(_11903_),
    .Y(_11914_));
 sky130_fd_sc_hd__nand2_1 _14120_ (.A(_10379_),
    .B(_11914_),
    .Y(_11925_));
 sky130_fd_sc_hd__xnor2_4 _14121_ (.A(_10379_),
    .B(_11914_),
    .Y(_11936_));
 sky130_fd_sc_hd__o21ba_2 _14122_ (.A1(_10148_),
    .A2(_10170_),
    .B1_N(_10159_),
    .X(_11947_));
 sky130_fd_sc_hd__nor2_2 _14123_ (.A(_11936_),
    .B(_11947_),
    .Y(_11958_));
 sky130_fd_sc_hd__and2_1 _14124_ (.A(_11936_),
    .B(_11947_),
    .X(_11969_));
 sky130_fd_sc_hd__nand2_1 _14125_ (.A(_11936_),
    .B(_11947_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2b_2 _14126_ (.A_N(_11958_),
    .B(_11980_),
    .Y(_11991_));
 sky130_fd_sc_hd__o2bb2ai_2 _14127_ (.A1_N(_11749_),
    .A2_N(_11760_),
    .B1(_11958_),
    .B2(_11969_),
    .Y(_12002_));
 sky130_fd_sc_hd__nand3b_2 _14128_ (.A_N(_11991_),
    .B(_11760_),
    .C(_11749_),
    .Y(_12012_));
 sky130_fd_sc_hd__nand2_1 _14129_ (.A(_12002_),
    .B(_12012_),
    .Y(_12023_));
 sky130_fd_sc_hd__o21a_1 _14130_ (.A1(_10422_),
    .A2(_10433_),
    .B1(_10302_),
    .X(_12034_));
 sky130_fd_sc_hd__o21ai_1 _14131_ (.A1(_10466_),
    .A2(_10280_),
    .B1(_10302_),
    .Y(_12045_));
 sky130_fd_sc_hd__nand3_2 _14132_ (.A(_12002_),
    .B(_12012_),
    .C(_12045_),
    .Y(_12056_));
 sky130_fd_sc_hd__inv_2 _14133_ (.A(_12056_),
    .Y(_12067_));
 sky130_fd_sc_hd__o2bb2ai_2 _14134_ (.A1_N(_12002_),
    .A2_N(_12012_),
    .B1(_12034_),
    .B2(_10280_),
    .Y(_12078_));
 sky130_fd_sc_hd__o2bb2ai_2 _14135_ (.A1_N(_12056_),
    .A2_N(_12078_),
    .B1(_10401_),
    .B2(_10411_),
    .Y(_12089_));
 sky130_fd_sc_hd__a21boi_1 _14136_ (.A1(_10302_),
    .A2(_12023_),
    .B1_N(_10422_),
    .Y(_12100_));
 sky130_fd_sc_hd__nand3_2 _14137_ (.A(_12078_),
    .B(_10422_),
    .C(_12056_),
    .Y(_12111_));
 sky130_fd_sc_hd__nand2_1 _14138_ (.A(_12089_),
    .B(_12111_),
    .Y(_12122_));
 sky130_fd_sc_hd__a21oi_1 _14139_ (.A1(_12089_),
    .A2(_12111_),
    .B1(_10860_),
    .Y(_12133_));
 sky130_fd_sc_hd__a21o_1 _14140_ (.A1(_12089_),
    .A2(_12111_),
    .B1(_10860_),
    .X(_12144_));
 sky130_fd_sc_hd__and3_1 _14141_ (.A(_10860_),
    .B(_12089_),
    .C(_12111_),
    .X(_12155_));
 sky130_fd_sc_hd__nand3_2 _14142_ (.A(_10860_),
    .B(_12089_),
    .C(_12111_),
    .Y(_12166_));
 sky130_fd_sc_hd__nor2_1 _14143_ (.A(_12133_),
    .B(_12155_),
    .Y(_12177_));
 sky130_fd_sc_hd__nand3_1 _14144_ (.A(_10664_),
    .B(_12144_),
    .C(_12166_),
    .Y(_12188_));
 sky130_fd_sc_hd__o22ai_1 _14145_ (.A1(_10642_),
    .A2(_10653_),
    .B1(_12133_),
    .B2(_12155_),
    .Y(_12199_));
 sky130_fd_sc_hd__nand2_1 _14146_ (.A(_12188_),
    .B(_12199_),
    .Y(_12210_));
 sky130_fd_sc_hd__a31o_1 _14147_ (.A1(_10631_),
    .A2(_10664_),
    .A3(_10708_),
    .B1(_12210_),
    .X(_12221_));
 sky130_fd_sc_hd__nand4_1 _14148_ (.A(_12177_),
    .B(_10664_),
    .C(_10631_),
    .D(_10697_),
    .Y(_12232_));
 sky130_fd_sc_hd__nand2_1 _14149_ (.A(_12221_),
    .B(_12232_),
    .Y(_12243_));
 sky130_fd_sc_hd__xor2_1 _14150_ (.A(_10849_),
    .B(_12243_),
    .X(net67));
 sky130_fd_sc_hd__or3_1 _14151_ (.A(_09358_),
    .B(_10609_),
    .C(_12133_),
    .X(_12264_));
 sky130_fd_sc_hd__nor3_1 _14152_ (.A(_09347_),
    .B(_10609_),
    .C(_12133_),
    .Y(_12275_));
 sky130_fd_sc_hd__or3_1 _14153_ (.A(_09347_),
    .B(_10609_),
    .C(_12133_),
    .X(_12286_));
 sky130_fd_sc_hd__a31o_1 _14154_ (.A1(_12002_),
    .A2(_12012_),
    .A3(_12045_),
    .B1(_10422_),
    .X(_12297_));
 sky130_fd_sc_hd__a21oi_1 _14155_ (.A1(_10422_),
    .A2(_12078_),
    .B1(_12067_),
    .Y(_12308_));
 sky130_fd_sc_hd__o21ai_1 _14156_ (.A1(_11991_),
    .A2(_11738_),
    .B1(_11760_),
    .Y(_12319_));
 sky130_fd_sc_hd__and2_4 _14157_ (.A(_03993_),
    .B(net36),
    .X(_12330_));
 sky130_fd_sc_hd__nand2b_4 _14158_ (.A_N(net35),
    .B(net36),
    .Y(_12341_));
 sky130_fd_sc_hd__nor2_8 _14159_ (.A(net36),
    .B(_03993_),
    .Y(_12352_));
 sky130_fd_sc_hd__nand2b_4 _14160_ (.A_N(net36),
    .B(net35),
    .Y(_12363_));
 sky130_fd_sc_hd__a21oi_1 _14161_ (.A1(_12341_),
    .A2(_12363_),
    .B1(_03176_),
    .Y(_12374_));
 sky130_fd_sc_hd__a21oi_1 _14162_ (.A1(_11892_),
    .A2(_11815_),
    .B1(_11870_),
    .Y(_12385_));
 sky130_fd_sc_hd__a21o_1 _14163_ (.A1(_11815_),
    .A2(_11892_),
    .B1(_11870_),
    .X(_12396_));
 sky130_fd_sc_hd__a22oi_2 _14164_ (.A1(net12),
    .A2(_11793_),
    .B1(_04539_),
    .B2(_11771_),
    .Y(_12406_));
 sky130_fd_sc_hd__and3b_1 _14165_ (.A_N(net34),
    .B(net64),
    .C(net23),
    .X(_12417_));
 sky130_fd_sc_hd__nand3_1 _14166_ (.A(_04419_),
    .B(_04452_),
    .C(_10313_),
    .Y(_12428_));
 sky130_fd_sc_hd__a31oi_2 _14167_ (.A1(net318),
    .A2(_04452_),
    .A3(_10313_),
    .B1(_12417_),
    .Y(_12439_));
 sky130_fd_sc_hd__nand3_1 _14168_ (.A(_04714_),
    .B(net267),
    .C(_08250_),
    .Y(_12450_));
 sky130_fd_sc_hd__nand2_1 _14169_ (.A(net26),
    .B(_08272_),
    .Y(_12461_));
 sky130_fd_sc_hd__a32oi_2 _14170_ (.A1(net315),
    .A2(net267),
    .A3(_08250_),
    .B1(_08272_),
    .B2(net26),
    .Y(_12472_));
 sky130_fd_sc_hd__o2111a_1 _14171_ (.A1(_03396_),
    .A2(_10346_),
    .B1(_12428_),
    .C1(_12450_),
    .D1(_12461_),
    .X(_12483_));
 sky130_fd_sc_hd__nand2_1 _14172_ (.A(_12439_),
    .B(_12472_),
    .Y(_12494_));
 sky130_fd_sc_hd__a21oi_1 _14173_ (.A1(_12450_),
    .A2(_12461_),
    .B1(_12439_),
    .Y(_12505_));
 sky130_fd_sc_hd__a21o_1 _14174_ (.A1(_12450_),
    .A2(_12461_),
    .B1(_12439_),
    .X(_12516_));
 sky130_fd_sc_hd__o21bai_1 _14175_ (.A1(_12439_),
    .A2(_12472_),
    .B1_N(_12406_),
    .Y(_12527_));
 sky130_fd_sc_hd__o21ai_1 _14176_ (.A1(_12483_),
    .A2(_12505_),
    .B1(_12406_),
    .Y(_12538_));
 sky130_fd_sc_hd__nand3_1 _14177_ (.A(_12516_),
    .B(_12406_),
    .C(_12494_),
    .Y(_12549_));
 sky130_fd_sc_hd__o21bai_1 _14178_ (.A1(_12483_),
    .A2(_12505_),
    .B1_N(_12406_),
    .Y(_12560_));
 sky130_fd_sc_hd__o211a_1 _14179_ (.A1(_12527_),
    .A2(_12483_),
    .B1(_12396_),
    .C1(_12538_),
    .X(_12571_));
 sky130_fd_sc_hd__o211ai_1 _14180_ (.A1(_12527_),
    .A2(_12483_),
    .B1(_12396_),
    .C1(_12538_),
    .Y(_12582_));
 sky130_fd_sc_hd__nand3_2 _14181_ (.A(_12560_),
    .B(_12385_),
    .C(_12549_),
    .Y(_12593_));
 sky130_fd_sc_hd__o211a_1 _14182_ (.A1(_12330_),
    .A2(_12352_),
    .B1(net1),
    .C1(_12593_),
    .X(_12604_));
 sky130_fd_sc_hd__a221o_1 _14183_ (.A1(_12341_),
    .A2(_12363_),
    .B1(_12582_),
    .B2(_12593_),
    .C1(_03176_),
    .X(_12615_));
 sky130_fd_sc_hd__nand3b_1 _14184_ (.A_N(_12374_),
    .B(_12582_),
    .C(_12593_),
    .Y(_12626_));
 sky130_fd_sc_hd__a21boi_1 _14185_ (.A1(_11047_),
    .A2(_10115_),
    .B1_N(_11058_),
    .Y(_12637_));
 sky130_fd_sc_hd__and3_1 _14186_ (.A(_12637_),
    .B(_12626_),
    .C(_12615_),
    .X(_12648_));
 sky130_fd_sc_hd__nand4_1 _14187_ (.A(_11058_),
    .B(_11091_),
    .C(_12615_),
    .D(_12626_),
    .Y(_12659_));
 sky130_fd_sc_hd__a21o_1 _14188_ (.A1(_12615_),
    .A2(_12626_),
    .B1(_12637_),
    .X(_12670_));
 sky130_fd_sc_hd__a22oi_2 _14189_ (.A1(_10379_),
    .A2(_11914_),
    .B1(_12659_),
    .B2(_12670_),
    .Y(_12681_));
 sky130_fd_sc_hd__and4_1 _14190_ (.A(_12659_),
    .B(_12670_),
    .C(_10379_),
    .D(_11914_),
    .X(_12692_));
 sky130_fd_sc_hd__nand4_1 _14191_ (.A(_12659_),
    .B(_12670_),
    .C(_10379_),
    .D(_11914_),
    .Y(_12703_));
 sky130_fd_sc_hd__nand2b_1 _14192_ (.A_N(_12681_),
    .B(_12703_),
    .Y(_12714_));
 sky130_fd_sc_hd__o21ai_1 _14193_ (.A1(_11102_),
    .A2(_11661_),
    .B1(_11650_),
    .Y(_12725_));
 sky130_fd_sc_hd__a21o_1 _14194_ (.A1(_10904_),
    .A2(_10981_),
    .B1(_10948_),
    .X(_12735_));
 sky130_fd_sc_hd__a21o_1 _14195_ (.A1(_11135_),
    .A2(_11201_),
    .B1(_11212_),
    .X(_12746_));
 sky130_fd_sc_hd__a32o_1 _14196_ (.A1(_04998_),
    .A2(_05009_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net27),
    .X(_12757_));
 sky130_fd_sc_hd__a32oi_4 _14197_ (.A1(_05414_),
    .A2(_05446_),
    .A3(net292),
    .B1(_06848_),
    .B2(net28),
    .Y(_12768_));
 sky130_fd_sc_hd__or3b_1 _14198_ (.A(net61),
    .B(_03835_),
    .C_N(net60),
    .X(_12779_));
 sky130_fd_sc_hd__nand3_1 _14199_ (.A(_05841_),
    .B(_05863_),
    .C(net299),
    .Y(_12790_));
 sky130_fd_sc_hd__a32oi_4 _14200_ (.A1(_05841_),
    .A2(_05863_),
    .A3(net299),
    .B1(_05710_),
    .B2(net29),
    .Y(_12801_));
 sky130_fd_sc_hd__a21o_1 _14201_ (.A1(_12779_),
    .A2(_12790_),
    .B1(_12768_),
    .X(_12812_));
 sky130_fd_sc_hd__nand2_1 _14202_ (.A(_12768_),
    .B(_12801_),
    .Y(_12823_));
 sky130_fd_sc_hd__nand3_4 _14203_ (.A(_12757_),
    .B(_12812_),
    .C(_12823_),
    .Y(_12834_));
 sky130_fd_sc_hd__a21o_1 _14204_ (.A1(_12812_),
    .A2(_12823_),
    .B1(_12757_),
    .X(_12845_));
 sky130_fd_sc_hd__a21o_2 _14205_ (.A1(_12834_),
    .A2(_12845_),
    .B1(_12746_),
    .X(_12856_));
 sky130_fd_sc_hd__o211ai_4 _14206_ (.A1(_11212_),
    .A2(_11255_),
    .B1(_12834_),
    .C1(_12845_),
    .Y(_12867_));
 sky130_fd_sc_hd__a21oi_2 _14207_ (.A1(_12856_),
    .A2(_12867_),
    .B1(_12735_),
    .Y(_12878_));
 sky130_fd_sc_hd__and3_1 _14208_ (.A(_12735_),
    .B(_12856_),
    .C(_12867_),
    .X(_12889_));
 sky130_fd_sc_hd__a22oi_4 _14209_ (.A1(_10959_),
    .A2(_10992_),
    .B1(_12856_),
    .B2(_12867_),
    .Y(_12900_));
 sky130_fd_sc_hd__and4_1 _14210_ (.A(_10959_),
    .B(_10992_),
    .C(_12856_),
    .D(_12867_),
    .X(_12911_));
 sky130_fd_sc_hd__o2bb2ai_4 _14211_ (.A1_N(_11310_),
    .A2_N(_11475_),
    .B1(net236),
    .B2(_11332_),
    .Y(_12922_));
 sky130_fd_sc_hd__a32o_2 _14212_ (.A1(_09698_),
    .A2(_04342_),
    .A3(net255),
    .B1(_04364_),
    .B2(net2),
    .X(_12933_));
 sky130_fd_sc_hd__o211ai_2 _14213_ (.A1(_06530_),
    .A2(_11387_),
    .B1(_04484_),
    .C1(_11354_),
    .Y(_12944_));
 sky130_fd_sc_hd__nor2_1 _14214_ (.A(_03982_),
    .B(_04331_),
    .Y(_12955_));
 sky130_fd_sc_hd__or3_1 _14215_ (.A(net44),
    .B(_03982_),
    .C(_03286_),
    .X(_12966_));
 sky130_fd_sc_hd__o21bai_4 _14216_ (.A1(net267),
    .A2(_11409_),
    .B1_N(_04004_),
    .Y(_12977_));
 sky130_fd_sc_hd__nand4_4 _14217_ (.A(_04736_),
    .B(_05852_),
    .C(_03916_),
    .D(_04004_),
    .Y(_12988_));
 sky130_fd_sc_hd__nand4_4 _14218_ (.A(net312),
    .B(_06497_),
    .C(_11376_),
    .D(_04004_),
    .Y(_12999_));
 sky130_fd_sc_hd__o31a_4 _14219_ (.A1(net3),
    .A2(_09665_),
    .A3(_12988_),
    .B1(_12977_),
    .X(_13010_));
 sky130_fd_sc_hd__o21ai_4 _14220_ (.A1(_11387_),
    .A2(_12988_),
    .B1(_12977_),
    .Y(_13021_));
 sky130_fd_sc_hd__nand3_1 _14221_ (.A(_12977_),
    .B(_12999_),
    .C(net33),
    .Y(_13032_));
 sky130_fd_sc_hd__nand4_2 _14222_ (.A(_12977_),
    .B(_12999_),
    .C(net33),
    .D(_12955_),
    .Y(_13043_));
 sky130_fd_sc_hd__nand3_4 _14223_ (.A(_12944_),
    .B(_12966_),
    .C(_13032_),
    .Y(_13054_));
 sky130_fd_sc_hd__a21oi_1 _14224_ (.A1(_13043_),
    .A2(_13054_),
    .B1(_12933_),
    .Y(_13064_));
 sky130_fd_sc_hd__a21o_1 _14225_ (.A1(_13043_),
    .A2(_13054_),
    .B1(_12933_),
    .X(_13075_));
 sky130_fd_sc_hd__o311a_1 _14226_ (.A1(_03286_),
    .A2(_12966_),
    .A3(_13021_),
    .B1(_13054_),
    .C1(_12933_),
    .X(_13086_));
 sky130_fd_sc_hd__nand3_2 _14227_ (.A(_12933_),
    .B(_13043_),
    .C(_13054_),
    .Y(_13097_));
 sky130_fd_sc_hd__a21oi_4 _14228_ (.A1(_13075_),
    .A2(_13097_),
    .B1(_12922_),
    .Y(_13108_));
 sky130_fd_sc_hd__o21bai_4 _14229_ (.A1(_13064_),
    .A2(_13086_),
    .B1_N(_12922_),
    .Y(_13119_));
 sky130_fd_sc_hd__nand3_4 _14230_ (.A(_12922_),
    .B(_13075_),
    .C(_13097_),
    .Y(_13130_));
 sky130_fd_sc_hd__a22oi_2 _14231_ (.A1(net30),
    .A2(_05249_),
    .B1(_06541_),
    .B2(_05227_),
    .Y(_13141_));
 sky130_fd_sc_hd__a32o_1 _14232_ (.A1(_06486_),
    .A2(_06530_),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net30),
    .X(_13152_));
 sky130_fd_sc_hd__a32oi_4 _14233_ (.A1(_07242_),
    .A2(net258),
    .A3(net305),
    .B1(_04911_),
    .B2(net31),
    .Y(_13163_));
 sky130_fd_sc_hd__or3b_1 _14234_ (.A(net58),
    .B(_03949_),
    .C_N(net55),
    .X(_13174_));
 sky130_fd_sc_hd__o211ai_2 _14235_ (.A1(_06530_),
    .A2(_08656_),
    .B1(net317),
    .C1(_08700_),
    .Y(_13185_));
 sky130_fd_sc_hd__a21oi_2 _14236_ (.A1(_13174_),
    .A2(_13185_),
    .B1(_13163_),
    .Y(_13196_));
 sky130_fd_sc_hd__a21o_1 _14237_ (.A1(_13174_),
    .A2(_13185_),
    .B1(_13163_),
    .X(_13207_));
 sky130_fd_sc_hd__o221a_1 _14238_ (.A1(_03949_),
    .A2(_04660_),
    .B1(_08711_),
    .B2(_04638_),
    .C1(_13163_),
    .X(_13218_));
 sky130_fd_sc_hd__o221ai_4 _14239_ (.A1(_03949_),
    .A2(_04660_),
    .B1(_08711_),
    .B2(_04638_),
    .C1(_13163_),
    .Y(_13229_));
 sky130_fd_sc_hd__a21oi_1 _14240_ (.A1(_13207_),
    .A2(_13229_),
    .B1(_13152_),
    .Y(_13240_));
 sky130_fd_sc_hd__o21ai_2 _14241_ (.A1(_13196_),
    .A2(_13218_),
    .B1(_13141_),
    .Y(_13251_));
 sky130_fd_sc_hd__nand3_2 _14242_ (.A(_13152_),
    .B(_13207_),
    .C(_13229_),
    .Y(_13262_));
 sky130_fd_sc_hd__inv_2 _14243_ (.A(_13262_),
    .Y(_13273_));
 sky130_fd_sc_hd__nand2_2 _14244_ (.A(_13251_),
    .B(_13262_),
    .Y(_13284_));
 sky130_fd_sc_hd__o2bb2ai_4 _14245_ (.A1_N(_13119_),
    .A2_N(_13130_),
    .B1(_13240_),
    .B2(_13273_),
    .Y(_13295_));
 sky130_fd_sc_hd__nand4_4 _14246_ (.A(_13119_),
    .B(_13130_),
    .C(_13251_),
    .D(_13262_),
    .Y(_13306_));
 sky130_fd_sc_hd__a311oi_4 _14247_ (.A1(_11497_),
    .A2(_11508_),
    .A3(_11288_),
    .B1(_11255_),
    .C1(_11233_),
    .Y(_13317_));
 sky130_fd_sc_hd__o21ai_1 _14248_ (.A1(_11277_),
    .A2(_11541_),
    .B1(_11574_),
    .Y(_13328_));
 sky130_fd_sc_hd__o211a_2 _14249_ (.A1(_11563_),
    .A2(_13317_),
    .B1(_13306_),
    .C1(_13295_),
    .X(_13339_));
 sky130_fd_sc_hd__o211ai_4 _14250_ (.A1(_11563_),
    .A2(_13317_),
    .B1(_13306_),
    .C1(_13295_),
    .Y(_13350_));
 sky130_fd_sc_hd__a21oi_2 _14251_ (.A1(_13295_),
    .A2(_13306_),
    .B1(_13328_),
    .Y(_13361_));
 sky130_fd_sc_hd__a21o_1 _14252_ (.A1(_13295_),
    .A2(_13306_),
    .B1(_13328_),
    .X(_13371_));
 sky130_fd_sc_hd__o21ai_4 _14253_ (.A1(_12900_),
    .A2(_12911_),
    .B1(_13371_),
    .Y(_00000_));
 sky130_fd_sc_hd__o211ai_2 _14254_ (.A1(_12900_),
    .A2(_12911_),
    .B1(_13350_),
    .C1(_13371_),
    .Y(_00011_));
 sky130_fd_sc_hd__o22ai_4 _14255_ (.A1(_12878_),
    .A2(_12889_),
    .B1(_13339_),
    .B2(_13361_),
    .Y(_00022_));
 sky130_fd_sc_hd__o211a_1 _14256_ (.A1(_11639_),
    .A2(_11705_),
    .B1(_00011_),
    .C1(_00022_),
    .X(_00033_));
 sky130_fd_sc_hd__o221ai_4 _14257_ (.A1(_11639_),
    .A2(_11705_),
    .B1(_13339_),
    .B2(_00000_),
    .C1(_00022_),
    .Y(_00044_));
 sky130_fd_sc_hd__a21oi_2 _14258_ (.A1(_00011_),
    .A2(_00022_),
    .B1(_12725_),
    .Y(_00055_));
 sky130_fd_sc_hd__a21o_1 _14259_ (.A1(_00011_),
    .A2(_00022_),
    .B1(_12725_),
    .X(_00066_));
 sky130_fd_sc_hd__o211ai_2 _14260_ (.A1(_12681_),
    .A2(_12692_),
    .B1(_00044_),
    .C1(_00066_),
    .Y(_00077_));
 sky130_fd_sc_hd__o21bai_2 _14261_ (.A1(_00033_),
    .A2(_00055_),
    .B1_N(_12714_),
    .Y(_00088_));
 sky130_fd_sc_hd__nor2_1 _14262_ (.A(_12714_),
    .B(_00055_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand3b_1 _14263_ (.A_N(_12714_),
    .B(_00044_),
    .C(_00066_),
    .Y(_00110_));
 sky130_fd_sc_hd__o21ai_1 _14264_ (.A1(_00033_),
    .A2(_00055_),
    .B1(_12714_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand3_2 _14265_ (.A(_00121_),
    .B(_12319_),
    .C(_00110_),
    .Y(_00132_));
 sky130_fd_sc_hd__o2111a_1 _14266_ (.A1(_11991_),
    .A2(_11738_),
    .B1(_11760_),
    .C1(_00077_),
    .D1(_00088_),
    .X(_00143_));
 sky130_fd_sc_hd__o2111ai_4 _14267_ (.A1(_11991_),
    .A2(_11738_),
    .B1(_11760_),
    .C1(_00077_),
    .D1(_00088_),
    .Y(_00154_));
 sky130_fd_sc_hd__nand3_2 _14268_ (.A(_00132_),
    .B(_00154_),
    .C(_11958_),
    .Y(_00165_));
 sky130_fd_sc_hd__o2bb2ai_2 _14269_ (.A1_N(_00132_),
    .A2_N(_00154_),
    .B1(_11936_),
    .B2(_11947_),
    .Y(_00176_));
 sky130_fd_sc_hd__a21bo_1 _14270_ (.A1(_00132_),
    .A2(_00154_),
    .B1_N(_11958_),
    .X(_00187_));
 sky130_fd_sc_hd__o211ai_2 _14271_ (.A1(_11936_),
    .A2(_11947_),
    .B1(_00132_),
    .C1(_00154_),
    .Y(_00198_));
 sky130_fd_sc_hd__o211a_2 _14272_ (.A1(_12067_),
    .A2(_12100_),
    .B1(_00165_),
    .C1(_00176_),
    .X(_00209_));
 sky130_fd_sc_hd__o211ai_1 _14273_ (.A1(_12067_),
    .A2(_12100_),
    .B1(_00165_),
    .C1(_00176_),
    .Y(_00220_));
 sky130_fd_sc_hd__a22oi_2 _14274_ (.A1(_12078_),
    .A2(_12297_),
    .B1(_00165_),
    .B2(_00176_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand3_1 _14275_ (.A(_12308_),
    .B(_00187_),
    .C(_00198_),
    .Y(_00242_));
 sky130_fd_sc_hd__a2bb2oi_1 _14276_ (.A1_N(_10871_),
    .A2_N(_12122_),
    .B1(_00220_),
    .B2(_00242_),
    .Y(_00253_));
 sky130_fd_sc_hd__o22ai_1 _14277_ (.A1(_12122_),
    .A2(_10871_),
    .B1(_00231_),
    .B2(_00209_),
    .Y(_00264_));
 sky130_fd_sc_hd__a31oi_1 _14278_ (.A1(_12308_),
    .A2(_00187_),
    .A3(_00198_),
    .B1(_12166_),
    .Y(_00275_));
 sky130_fd_sc_hd__a31o_1 _14279_ (.A1(_12308_),
    .A2(_00187_),
    .A3(_00198_),
    .B1(_12166_),
    .X(_00286_));
 sky130_fd_sc_hd__o21ai_1 _14280_ (.A1(_12166_),
    .A2(_00231_),
    .B1(_00264_),
    .Y(_00297_));
 sky130_fd_sc_hd__and3_1 _14281_ (.A(_12275_),
    .B(_00220_),
    .C(_00242_),
    .X(_00308_));
 sky130_fd_sc_hd__nand2_1 _14282_ (.A(_00264_),
    .B(_12275_),
    .Y(_00318_));
 sky130_fd_sc_hd__o2bb2ai_1 _14283_ (.A1_N(_12144_),
    .A2_N(_10642_),
    .B1(_00275_),
    .B2(_00253_),
    .Y(_00329_));
 sky130_fd_sc_hd__a22oi_2 _14284_ (.A1(_12144_),
    .A2(_10653_),
    .B1(_00329_),
    .B2(_00318_),
    .Y(_00340_));
 sky130_fd_sc_hd__a21oi_1 _14285_ (.A1(_12286_),
    .A2(_00297_),
    .B1(_12264_),
    .Y(_00351_));
 sky130_fd_sc_hd__nor2_1 _14286_ (.A(_00340_),
    .B(_00351_),
    .Y(_00362_));
 sky130_fd_sc_hd__o2bb2ai_2 _14287_ (.A1_N(_10849_),
    .A2_N(_12232_),
    .B1(_12210_),
    .B2(_10741_),
    .Y(_00373_));
 sky130_fd_sc_hd__xnor2_1 _14288_ (.A(_00362_),
    .B(_00373_),
    .Y(net68));
 sky130_fd_sc_hd__o21bai_2 _14289_ (.A1(_00340_),
    .A2(_00373_),
    .B1_N(_00351_),
    .Y(_00394_));
 sky130_fd_sc_hd__o21ai_1 _14290_ (.A1(_11925_),
    .A2(_12648_),
    .B1(_12670_),
    .Y(_00405_));
 sky130_fd_sc_hd__o31ai_1 _14291_ (.A1(_12878_),
    .A2(_12889_),
    .A3(_13361_),
    .B1(_13350_),
    .Y(_00416_));
 sky130_fd_sc_hd__o21ai_2 _14292_ (.A1(_13108_),
    .A2(_13284_),
    .B1(_13130_),
    .Y(_00427_));
 sky130_fd_sc_hd__o21a_1 _14293_ (.A1(_13108_),
    .A2(_13284_),
    .B1(_13130_),
    .X(_00438_));
 sky130_fd_sc_hd__o22a_1 _14294_ (.A1(_03938_),
    .A2(_05260_),
    .B1(_07263_),
    .B2(_05238_),
    .X(_00449_));
 sky130_fd_sc_hd__a32o_1 _14295_ (.A1(_07242_),
    .A2(net258),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net31),
    .X(_00460_));
 sky130_fd_sc_hd__or3b_1 _14296_ (.A(net58),
    .B(_03960_),
    .C_N(net55),
    .X(_00471_));
 sky130_fd_sc_hd__o211ai_1 _14297_ (.A1(_06530_),
    .A2(_09665_),
    .B1(net317),
    .C1(_09698_),
    .Y(_00482_));
 sky130_fd_sc_hd__and3b_1 _14298_ (.A_N(net59),
    .B(net32),
    .C(net58),
    .X(_00493_));
 sky130_fd_sc_hd__o311a_1 _14299_ (.A1(net267),
    .A2(_06508_),
    .A3(_08656_),
    .B1(net305),
    .C1(_08700_),
    .X(_00504_));
 sky130_fd_sc_hd__a31oi_4 _14300_ (.A1(_08700_),
    .A2(net305),
    .A3(net256),
    .B1(_00493_),
    .Y(_00515_));
 sky130_fd_sc_hd__a21oi_1 _14301_ (.A1(_00471_),
    .A2(_00482_),
    .B1(_00515_),
    .Y(_00526_));
 sky130_fd_sc_hd__o2bb2ai_1 _14302_ (.A1_N(_00471_),
    .A2_N(_00482_),
    .B1(_00493_),
    .B2(_00504_),
    .Y(_00537_));
 sky130_fd_sc_hd__o221a_1 _14303_ (.A1(_03960_),
    .A2(_04660_),
    .B1(_09720_),
    .B2(_04638_),
    .C1(_00515_),
    .X(_00548_));
 sky130_fd_sc_hd__o221ai_4 _14304_ (.A1(_03960_),
    .A2(_04660_),
    .B1(_09720_),
    .B2(_04638_),
    .C1(_00515_),
    .Y(_00559_));
 sky130_fd_sc_hd__o21ai_2 _14305_ (.A1(_00526_),
    .A2(_00548_),
    .B1(_00460_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand3_2 _14306_ (.A(_00537_),
    .B(_00559_),
    .C(_00449_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_2 _14307_ (.A(_00570_),
    .B(_00581_),
    .Y(_00592_));
 sky130_fd_sc_hd__a32o_2 _14308_ (.A1(_11354_),
    .A2(_11431_),
    .A3(_04342_),
    .B1(_04364_),
    .B2(net3),
    .X(_00603_));
 sky130_fd_sc_hd__a41oi_4 _14309_ (.A1(net307),
    .A2(net293),
    .A3(net288),
    .A4(_04004_),
    .B1(_04015_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_8 _14310_ (.A(net251),
    .B(net5),
    .Y(_00625_));
 sky130_fd_sc_hd__nor2_4 _14311_ (.A(net4),
    .B(net5),
    .Y(_00635_));
 sky130_fd_sc_hd__or2_4 _14312_ (.A(net4),
    .B(net5),
    .X(_00646_));
 sky130_fd_sc_hd__nand4_4 _14313_ (.A(net307),
    .B(net293),
    .C(net287),
    .D(_00635_),
    .Y(_00657_));
 sky130_fd_sc_hd__o21ai_4 _14314_ (.A1(_11431_),
    .A2(_00646_),
    .B1(_00625_),
    .Y(_00668_));
 sky130_fd_sc_hd__o211ai_2 _14315_ (.A1(_11431_),
    .A2(_00646_),
    .B1(net33),
    .C1(_00625_),
    .Y(_00679_));
 sky130_fd_sc_hd__nor2_1 _14316_ (.A(_04004_),
    .B(_04331_),
    .Y(_00690_));
 sky130_fd_sc_hd__or3_2 _14317_ (.A(net44),
    .B(_04004_),
    .C(_03286_),
    .X(_00701_));
 sky130_fd_sc_hd__a31oi_4 _14318_ (.A1(_12977_),
    .A2(_12999_),
    .A3(_04484_),
    .B1(_00690_),
    .Y(_00712_));
 sky130_fd_sc_hd__o21ai_4 _14319_ (.A1(_03286_),
    .A2(_00668_),
    .B1(_00712_),
    .Y(_00723_));
 sky130_fd_sc_hd__and3_1 _14320_ (.A(net4),
    .B(_04320_),
    .C(_04015_),
    .X(_00734_));
 sky130_fd_sc_hd__o2bb2ai_2 _14321_ (.A1_N(_00712_),
    .A2_N(_00679_),
    .B1(net5),
    .B2(_00701_),
    .Y(_00745_));
 sky130_fd_sc_hd__o211ai_4 _14322_ (.A1(_00701_),
    .A2(net5),
    .B1(_00603_),
    .C1(_00723_),
    .Y(_00756_));
 sky130_fd_sc_hd__o221ai_4 _14323_ (.A1(_03982_),
    .A2(_04375_),
    .B1(net236),
    .B2(_04353_),
    .C1(_00745_),
    .Y(_00767_));
 sky130_fd_sc_hd__a211o_1 _14324_ (.A1(_00679_),
    .A2(_00712_),
    .B1(_00734_),
    .C1(_00603_),
    .X(_00778_));
 sky130_fd_sc_hd__nand2_1 _14325_ (.A(_00603_),
    .B(_00745_),
    .Y(_00789_));
 sky130_fd_sc_hd__a32oi_4 _14326_ (.A1(net33),
    .A2(_12955_),
    .A3(_13010_),
    .B1(_13054_),
    .B2(_12933_),
    .Y(_00800_));
 sky130_fd_sc_hd__a32o_2 _14327_ (.A1(net33),
    .A2(_12955_),
    .A3(_13010_),
    .B1(_13054_),
    .B2(_12933_),
    .X(_00811_));
 sky130_fd_sc_hd__nand3_4 _14328_ (.A(_00778_),
    .B(_00789_),
    .C(_00800_),
    .Y(_00822_));
 sky130_fd_sc_hd__nand3_2 _14329_ (.A(_00756_),
    .B(_00767_),
    .C(_00811_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand3_1 _14330_ (.A(_00592_),
    .B(_00822_),
    .C(_00833_),
    .Y(_00844_));
 sky130_fd_sc_hd__a21o_1 _14331_ (.A1(_00822_),
    .A2(_00833_),
    .B1(_00592_),
    .X(_00855_));
 sky130_fd_sc_hd__nand4_4 _14332_ (.A(_00570_),
    .B(_00581_),
    .C(_00822_),
    .D(_00833_),
    .Y(_00866_));
 sky130_fd_sc_hd__a22o_2 _14333_ (.A1(_00570_),
    .A2(_00581_),
    .B1(_00822_),
    .B2(_00833_),
    .X(_00877_));
 sky130_fd_sc_hd__and3_1 _14334_ (.A(_00855_),
    .B(_00427_),
    .C(_00844_),
    .X(_00888_));
 sky130_fd_sc_hd__nand3_4 _14335_ (.A(_00855_),
    .B(_00427_),
    .C(_00844_),
    .Y(_00899_));
 sky130_fd_sc_hd__o2111ai_4 _14336_ (.A1(_13284_),
    .A2(_13108_),
    .B1(_13130_),
    .C1(_00866_),
    .D1(_00877_),
    .Y(_00910_));
 sky130_fd_sc_hd__o21ai_2 _14337_ (.A1(_12768_),
    .A2(_12801_),
    .B1(_12834_),
    .Y(_00921_));
 sky130_fd_sc_hd__a32o_1 _14338_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net28),
    .X(_00931_));
 sky130_fd_sc_hd__or3b_1 _14339_ (.A(_03835_),
    .B(net62),
    .C_N(net61),
    .X(_00942_));
 sky130_fd_sc_hd__nand3_1 _14340_ (.A(_05841_),
    .B(_05863_),
    .C(net292),
    .Y(_00953_));
 sky130_fd_sc_hd__nor2_1 _14341_ (.A(_03916_),
    .B(net298),
    .Y(_00964_));
 sky130_fd_sc_hd__o311a_1 _14342_ (.A1(net26),
    .A2(_04452_),
    .A3(_06508_),
    .B1(net299),
    .C1(_06486_),
    .X(_00975_));
 sky130_fd_sc_hd__a31oi_1 _14343_ (.A1(_06486_),
    .A2(_06530_),
    .A3(net299),
    .B1(_00964_),
    .Y(_00986_));
 sky130_fd_sc_hd__o2bb2ai_2 _14344_ (.A1_N(_00942_),
    .A2_N(_00953_),
    .B1(_00964_),
    .B2(_00975_),
    .Y(_00997_));
 sky130_fd_sc_hd__o211ai_2 _14345_ (.A1(_03835_),
    .A2(_06859_),
    .B1(_00953_),
    .C1(_00986_),
    .Y(_01008_));
 sky130_fd_sc_hd__a21oi_1 _14346_ (.A1(_00997_),
    .A2(_01008_),
    .B1(_00931_),
    .Y(_01019_));
 sky130_fd_sc_hd__a21o_1 _14347_ (.A1(_00997_),
    .A2(_01008_),
    .B1(_00931_),
    .X(_01030_));
 sky130_fd_sc_hd__and3_1 _14348_ (.A(_00931_),
    .B(_00997_),
    .C(_01008_),
    .X(_01041_));
 sky130_fd_sc_hd__nand3_2 _14349_ (.A(_00931_),
    .B(_00997_),
    .C(_01008_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand2_1 _14350_ (.A(_01030_),
    .B(_01052_),
    .Y(_01063_));
 sky130_fd_sc_hd__a31oi_1 _14351_ (.A1(_13163_),
    .A2(_13174_),
    .A3(_13185_),
    .B1(_13141_),
    .Y(_01074_));
 sky130_fd_sc_hd__a21oi_2 _14352_ (.A1(_13152_),
    .A2(_13229_),
    .B1(_13196_),
    .Y(_01085_));
 sky130_fd_sc_hd__o221a_2 _14353_ (.A1(_13141_),
    .A2(_13218_),
    .B1(_01019_),
    .B2(_01041_),
    .C1(_13207_),
    .X(_01096_));
 sky130_fd_sc_hd__o21ai_1 _14354_ (.A1(_01019_),
    .A2(_01041_),
    .B1(_01085_),
    .Y(_01107_));
 sky130_fd_sc_hd__o211ai_2 _14355_ (.A1(_13196_),
    .A2(_01074_),
    .B1(_01052_),
    .C1(_01030_),
    .Y(_01118_));
 sky130_fd_sc_hd__a21oi_1 _14356_ (.A1(_01107_),
    .A2(_01118_),
    .B1(_00921_),
    .Y(_01129_));
 sky130_fd_sc_hd__a21o_1 _14357_ (.A1(_01107_),
    .A2(_01118_),
    .B1(_00921_),
    .X(_01140_));
 sky130_fd_sc_hd__o21ai_2 _14358_ (.A1(_01063_),
    .A2(_01085_),
    .B1(_00921_),
    .Y(_01151_));
 sky130_fd_sc_hd__and3_1 _14359_ (.A(_00921_),
    .B(_01107_),
    .C(_01118_),
    .X(_01162_));
 sky130_fd_sc_hd__o21a_1 _14360_ (.A1(_01096_),
    .A2(_01151_),
    .B1(_01140_),
    .X(_01173_));
 sky130_fd_sc_hd__o21ai_2 _14361_ (.A1(_01096_),
    .A2(_01151_),
    .B1(_01140_),
    .Y(_01184_));
 sky130_fd_sc_hd__a21oi_2 _14362_ (.A1(_00899_),
    .A2(_00910_),
    .B1(_01173_),
    .Y(_01195_));
 sky130_fd_sc_hd__o2bb2ai_1 _14363_ (.A1_N(_00899_),
    .A2_N(_00910_),
    .B1(_01129_),
    .B2(_01162_),
    .Y(_01206_));
 sky130_fd_sc_hd__a31oi_4 _14364_ (.A1(_00438_),
    .A2(_00866_),
    .A3(_00877_),
    .B1(_01184_),
    .Y(_01216_));
 sky130_fd_sc_hd__o2111ai_4 _14365_ (.A1(_01096_),
    .A2(_01151_),
    .B1(_01140_),
    .C1(_00899_),
    .D1(_00910_),
    .Y(_01227_));
 sky130_fd_sc_hd__a21oi_1 _14366_ (.A1(_01206_),
    .A2(_01227_),
    .B1(_00416_),
    .Y(_01238_));
 sky130_fd_sc_hd__a21o_1 _14367_ (.A1(_01206_),
    .A2(_01227_),
    .B1(_00416_),
    .X(_01249_));
 sky130_fd_sc_hd__a221oi_4 _14368_ (.A1(_01216_),
    .A2(_00899_),
    .B1(_00000_),
    .B2(_13350_),
    .C1(_01195_),
    .Y(_01260_));
 sky130_fd_sc_hd__a221o_1 _14369_ (.A1(_01216_),
    .A2(_00899_),
    .B1(_00000_),
    .B2(_13350_),
    .C1(_01195_),
    .X(_01271_));
 sky130_fd_sc_hd__a31o_1 _14370_ (.A1(_12746_),
    .A2(_12834_),
    .A3(_12845_),
    .B1(_12735_),
    .X(_01282_));
 sky130_fd_sc_hd__and2b_4 _14371_ (.A_N(net36),
    .B(net37),
    .X(_01293_));
 sky130_fd_sc_hd__nand2b_4 _14372_ (.A_N(net36),
    .B(net37),
    .Y(_01304_));
 sky130_fd_sc_hd__and2b_4 _14373_ (.A_N(net37),
    .B(net36),
    .X(_01315_));
 sky130_fd_sc_hd__nand2b_4 _14374_ (.A_N(net37),
    .B(net36),
    .Y(_01326_));
 sky130_fd_sc_hd__a21oi_2 _14375_ (.A1(_01304_),
    .A2(_01326_),
    .B1(_03176_),
    .Y(_01337_));
 sky130_fd_sc_hd__a22o_1 _14376_ (.A1(net12),
    .A2(_12352_),
    .B1(_04539_),
    .B2(_12330_),
    .X(_01348_));
 sky130_fd_sc_hd__nand2_1 _14377_ (.A(_01348_),
    .B(_01337_),
    .Y(_01359_));
 sky130_fd_sc_hd__a221o_1 _14378_ (.A1(net12),
    .A2(_12352_),
    .B1(_12330_),
    .B2(_04539_),
    .C1(_01337_),
    .X(_01370_));
 sky130_fd_sc_hd__nand2_1 _14379_ (.A(_01359_),
    .B(_01370_),
    .Y(_01381_));
 sky130_fd_sc_hd__inv_2 _14380_ (.A(_01381_),
    .Y(_01392_));
 sky130_fd_sc_hd__a32o_1 _14381_ (.A1(_11771_),
    .A2(_04452_),
    .A3(net318),
    .B1(net23),
    .B2(_11793_),
    .X(_01403_));
 sky130_fd_sc_hd__or3b_1 _14382_ (.A(_03616_),
    .B(net64),
    .C_N(net63),
    .X(_01414_));
 sky130_fd_sc_hd__nand3_1 _14383_ (.A(_04998_),
    .B(_05009_),
    .C(_08250_),
    .Y(_01425_));
 sky130_fd_sc_hd__a32oi_2 _14384_ (.A1(net315),
    .A2(net267),
    .A3(_10313_),
    .B1(_10335_),
    .B2(net26),
    .Y(_01436_));
 sky130_fd_sc_hd__a21o_1 _14385_ (.A1(_01414_),
    .A2(_01425_),
    .B1(_01436_),
    .X(_01447_));
 sky130_fd_sc_hd__o211ai_2 _14386_ (.A1(_03616_),
    .A2(_08283_),
    .B1(_01425_),
    .C1(_01436_),
    .Y(_01458_));
 sky130_fd_sc_hd__and3_1 _14387_ (.A(_01403_),
    .B(_01447_),
    .C(_01458_),
    .X(_01469_));
 sky130_fd_sc_hd__nand3_1 _14388_ (.A(_01403_),
    .B(_01447_),
    .C(_01458_),
    .Y(_01480_));
 sky130_fd_sc_hd__a21oi_2 _14389_ (.A1(_01447_),
    .A2(_01458_),
    .B1(_01403_),
    .Y(_01490_));
 sky130_fd_sc_hd__o21a_1 _14390_ (.A1(_12406_),
    .A2(_12483_),
    .B1(_12516_),
    .X(_01501_));
 sky130_fd_sc_hd__o21a_1 _14391_ (.A1(_01469_),
    .A2(_01490_),
    .B1(_01501_),
    .X(_01512_));
 sky130_fd_sc_hd__o21ai_2 _14392_ (.A1(_01469_),
    .A2(_01490_),
    .B1(_01501_),
    .Y(_01523_));
 sky130_fd_sc_hd__nor3_2 _14393_ (.A(_01501_),
    .B(_01490_),
    .C(_01469_),
    .Y(_01534_));
 sky130_fd_sc_hd__nand3b_2 _14394_ (.A_N(_01534_),
    .B(_01392_),
    .C(_01523_),
    .Y(_01545_));
 sky130_fd_sc_hd__o21ai_2 _14395_ (.A1(_01512_),
    .A2(_01534_),
    .B1(_01381_),
    .Y(_01556_));
 sky130_fd_sc_hd__a22oi_4 _14396_ (.A1(_12856_),
    .A2(_01282_),
    .B1(_01545_),
    .B2(_01556_),
    .Y(_01567_));
 sky130_fd_sc_hd__and4_1 _14397_ (.A(_12856_),
    .B(_01282_),
    .C(_01545_),
    .D(_01556_),
    .X(_01578_));
 sky130_fd_sc_hd__nand4_2 _14398_ (.A(_12856_),
    .B(_01282_),
    .C(_01545_),
    .D(_01556_),
    .Y(_01589_));
 sky130_fd_sc_hd__a21oi_2 _14399_ (.A1(_12374_),
    .A2(_12593_),
    .B1(_12571_),
    .Y(_01600_));
 sky130_fd_sc_hd__o22ai_1 _14400_ (.A1(_12571_),
    .A2(_12604_),
    .B1(_01567_),
    .B2(_01578_),
    .Y(_01611_));
 sky130_fd_sc_hd__nand3b_1 _14401_ (.A_N(_01567_),
    .B(_01589_),
    .C(_01600_),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _14402_ (.A(_01611_),
    .B(_01622_),
    .Y(_01633_));
 sky130_fd_sc_hd__o21bai_2 _14403_ (.A1(_01238_),
    .A2(_01260_),
    .B1_N(_01633_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand3_2 _14404_ (.A(_01249_),
    .B(_01271_),
    .C(_01633_),
    .Y(_01655_));
 sky130_fd_sc_hd__o21a_1 _14405_ (.A1(_12681_),
    .A2(_12692_),
    .B1(_00044_),
    .X(_01666_));
 sky130_fd_sc_hd__o2bb2ai_1 _14406_ (.A1_N(_01644_),
    .A2_N(_01655_),
    .B1(_01666_),
    .B2(_00055_),
    .Y(_01677_));
 sky130_fd_sc_hd__o211ai_4 _14407_ (.A1(_00033_),
    .A2(_00099_),
    .B1(_01644_),
    .C1(_01655_),
    .Y(_01688_));
 sky130_fd_sc_hd__nand3_2 _14408_ (.A(_01677_),
    .B(_01688_),
    .C(_00405_),
    .Y(_01699_));
 sky130_fd_sc_hd__a21o_1 _14409_ (.A1(_01677_),
    .A2(_01688_),
    .B1(_00405_),
    .X(_01710_));
 sky130_fd_sc_hd__o21a_1 _14410_ (.A1(_11936_),
    .A2(_11947_),
    .B1(_00132_),
    .X(_01721_));
 sky130_fd_sc_hd__a31o_1 _14411_ (.A1(_00121_),
    .A2(_12319_),
    .A3(_00110_),
    .B1(_11958_),
    .X(_01731_));
 sky130_fd_sc_hd__o2bb2ai_2 _14412_ (.A1_N(_01699_),
    .A2_N(_01710_),
    .B1(_01721_),
    .B2(_00143_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand4_2 _14413_ (.A(_00154_),
    .B(_01699_),
    .C(_01710_),
    .D(_01731_),
    .Y(_01753_));
 sky130_fd_sc_hd__a21oi_1 _14414_ (.A1(_01742_),
    .A2(_01753_),
    .B1(_00209_),
    .Y(_01764_));
 sky130_fd_sc_hd__a21o_1 _14415_ (.A1(_01742_),
    .A2(_01753_),
    .B1(_00209_),
    .X(_01775_));
 sky130_fd_sc_hd__and4b_1 _14416_ (.A_N(_12308_),
    .B(_00165_),
    .C(_00176_),
    .D(_01742_),
    .X(_01786_));
 sky130_fd_sc_hd__nand2_2 _14417_ (.A(_01742_),
    .B(_00209_),
    .Y(_01797_));
 sky130_fd_sc_hd__a22o_1 _14418_ (.A1(_00286_),
    .A2(_00318_),
    .B1(_01775_),
    .B2(_01797_),
    .X(_01808_));
 sky130_fd_sc_hd__nand4_1 _14419_ (.A(_00286_),
    .B(_00318_),
    .C(_01775_),
    .D(_01797_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _14420_ (.A(_01808_),
    .B(_01819_),
    .Y(_01830_));
 sky130_fd_sc_hd__xor2_1 _14421_ (.A(_00394_),
    .B(_01830_),
    .X(net69));
 sky130_fd_sc_hd__a22oi_4 _14422_ (.A1(_00308_),
    .A2(_01775_),
    .B1(_00394_),
    .B2(_01830_),
    .Y(_01851_));
 sky130_fd_sc_hd__a21oi_2 _14423_ (.A1(_01249_),
    .A2(_01633_),
    .B1(_01260_),
    .Y(_01862_));
 sky130_fd_sc_hd__a21o_1 _14424_ (.A1(_01249_),
    .A2(_01633_),
    .B1(_01260_),
    .X(_01873_));
 sky130_fd_sc_hd__a21oi_1 _14425_ (.A1(_00910_),
    .A2(_01173_),
    .B1(_00888_),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_2 _14426_ (.A(_00997_),
    .B(_01052_),
    .Y(_01895_));
 sky130_fd_sc_hd__a32o_1 _14427_ (.A1(_05841_),
    .A2(_05863_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net29),
    .X(_01906_));
 sky130_fd_sc_hd__or3b_2 _14428_ (.A(net62),
    .B(_03916_),
    .C_N(net61),
    .X(_01917_));
 sky130_fd_sc_hd__o211ai_4 _14429_ (.A1(net267),
    .A2(_06508_),
    .B1(net292),
    .C1(_06486_),
    .Y(_01928_));
 sky130_fd_sc_hd__or3b_4 _14430_ (.A(net61),
    .B(_03938_),
    .C_N(net60),
    .X(_01939_));
 sky130_fd_sc_hd__nand3_4 _14431_ (.A(_07242_),
    .B(net258),
    .C(net299),
    .Y(_01950_));
 sky130_fd_sc_hd__a22oi_4 _14432_ (.A1(_01917_),
    .A2(_01928_),
    .B1(_01939_),
    .B2(_01950_),
    .Y(_01961_));
 sky130_fd_sc_hd__a22o_1 _14433_ (.A1(_01917_),
    .A2(_01928_),
    .B1(_01939_),
    .B2(_01950_),
    .X(_01971_));
 sky130_fd_sc_hd__o2111a_1 _14434_ (.A1(_03916_),
    .A2(_06859_),
    .B1(_01928_),
    .C1(_01939_),
    .D1(_01950_),
    .X(_01982_));
 sky130_fd_sc_hd__o2111ai_4 _14435_ (.A1(_03916_),
    .A2(_06859_),
    .B1(_01928_),
    .C1(_01939_),
    .D1(_01950_),
    .Y(_01993_));
 sky130_fd_sc_hd__o21bai_4 _14436_ (.A1(_01961_),
    .A2(_01982_),
    .B1_N(_01906_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand3_2 _14437_ (.A(_01906_),
    .B(_01971_),
    .C(_01993_),
    .Y(_02015_));
 sky130_fd_sc_hd__nor2_1 _14438_ (.A(_00460_),
    .B(_00526_),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _14439_ (.A(_00537_),
    .B(_00449_),
    .Y(_02037_));
 sky130_fd_sc_hd__o2bb2ai_4 _14440_ (.A1_N(_02004_),
    .A2_N(_02015_),
    .B1(_02026_),
    .B2(_00548_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand4_4 _14441_ (.A(_00559_),
    .B(_02004_),
    .C(_02015_),
    .D(_02037_),
    .Y(_02059_));
 sky130_fd_sc_hd__a21oi_2 _14442_ (.A1(_02048_),
    .A2(_02059_),
    .B1(_01895_),
    .Y(_02070_));
 sky130_fd_sc_hd__a21o_1 _14443_ (.A1(_02048_),
    .A2(_02059_),
    .B1(_01895_),
    .X(_02081_));
 sky130_fd_sc_hd__and3_1 _14444_ (.A(_01895_),
    .B(_02048_),
    .C(_02059_),
    .X(_02092_));
 sky130_fd_sc_hd__nand3_2 _14445_ (.A(_01895_),
    .B(_02048_),
    .C(_02059_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_2 _14446_ (.A(_02081_),
    .B(_02103_),
    .Y(_02114_));
 sky130_fd_sc_hd__a32oi_4 _14447_ (.A1(_00756_),
    .A2(_00767_),
    .A3(_00811_),
    .B1(_00592_),
    .B2(_00822_),
    .Y(_02125_));
 sky130_fd_sc_hd__a32o_1 _14448_ (.A1(_00756_),
    .A2(_00767_),
    .A3(_00811_),
    .B1(_00592_),
    .B2(_00822_),
    .X(_02136_));
 sky130_fd_sc_hd__nor2_1 _14449_ (.A(_03949_),
    .B(_05260_),
    .Y(_02147_));
 sky130_fd_sc_hd__a31oi_4 _14450_ (.A1(_08700_),
    .A2(_05227_),
    .A3(net256),
    .B1(_02147_),
    .Y(_02158_));
 sky130_fd_sc_hd__a31o_1 _14451_ (.A1(_08700_),
    .A2(_05227_),
    .A3(net256),
    .B1(_02147_),
    .X(_02169_));
 sky130_fd_sc_hd__and3b_1 _14452_ (.A_N(net59),
    .B(net2),
    .C(net58),
    .X(_02180_));
 sky130_fd_sc_hd__a31oi_4 _14453_ (.A1(_09698_),
    .A2(net305),
    .A3(net255),
    .B1(_02180_),
    .Y(_02191_));
 sky130_fd_sc_hd__a31o_1 _14454_ (.A1(_09698_),
    .A2(net305),
    .A3(net255),
    .B1(_02180_),
    .X(_02202_));
 sky130_fd_sc_hd__a22oi_4 _14455_ (.A1(net3),
    .A2(_04649_),
    .B1(_11442_),
    .B2(net317),
    .Y(_02212_));
 sky130_fd_sc_hd__o22ai_1 _14456_ (.A1(_03982_),
    .A2(_04660_),
    .B1(net236),
    .B2(_04638_),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _14457_ (.A(_02191_),
    .B(_02212_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2_1 _14458_ (.A(_02202_),
    .B(_02223_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand2_2 _14459_ (.A(_02191_),
    .B(_02212_),
    .Y(_02256_));
 sky130_fd_sc_hd__a21o_1 _14460_ (.A1(_02245_),
    .A2(_02256_),
    .B1(_02158_),
    .X(_02267_));
 sky130_fd_sc_hd__nand3_1 _14461_ (.A(_02245_),
    .B(_02256_),
    .C(_02158_),
    .Y(_02278_));
 sky130_fd_sc_hd__o21ai_2 _14462_ (.A1(_02191_),
    .A2(_02212_),
    .B1(_02158_),
    .Y(_02289_));
 sky130_fd_sc_hd__a21oi_1 _14463_ (.A1(_02191_),
    .A2(_02212_),
    .B1(_02158_),
    .Y(_02300_));
 sky130_fd_sc_hd__a21o_1 _14464_ (.A1(_02245_),
    .A2(_02256_),
    .B1(_02169_),
    .X(_02311_));
 sky130_fd_sc_hd__nand3_1 _14465_ (.A(_02169_),
    .B(_02245_),
    .C(_02256_),
    .Y(_02322_));
 sky130_fd_sc_hd__nand2_2 _14466_ (.A(_02267_),
    .B(_02278_),
    .Y(_02333_));
 sky130_fd_sc_hd__a31o_1 _14467_ (.A1(net4),
    .A2(_04015_),
    .A3(_04320_),
    .B1(_00603_),
    .X(_02344_));
 sky130_fd_sc_hd__a32o_1 _14468_ (.A1(net4),
    .A2(_04320_),
    .A3(_04015_),
    .B1(_00723_),
    .B2(_00603_),
    .X(_02355_));
 sky130_fd_sc_hd__nor2_1 _14469_ (.A(_04004_),
    .B(_04375_),
    .Y(_02366_));
 sky130_fd_sc_hd__o311a_1 _14470_ (.A1(net3),
    .A2(_09665_),
    .A3(_12988_),
    .B1(net235),
    .C1(_04342_),
    .X(_02377_));
 sky130_fd_sc_hd__a31o_2 _14471_ (.A1(net235),
    .A2(_12999_),
    .A3(_04342_),
    .B1(_02366_),
    .X(_02388_));
 sky130_fd_sc_hd__nand3_1 _14472_ (.A(_00625_),
    .B(_00657_),
    .C(_04484_),
    .Y(_02399_));
 sky130_fd_sc_hd__a41oi_4 _14473_ (.A1(net307),
    .A2(net293),
    .A3(net288),
    .A4(_00635_),
    .B1(_04026_),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_8 _14474_ (.A(net250),
    .B(net6),
    .Y(_02421_));
 sky130_fd_sc_hd__nor3_4 _14475_ (.A(net4),
    .B(net5),
    .C(net6),
    .Y(_02432_));
 sky130_fd_sc_hd__or3_4 _14476_ (.A(net4),
    .B(net5),
    .C(net6),
    .X(_02442_));
 sky130_fd_sc_hd__nand4_4 _14477_ (.A(net310),
    .B(net294),
    .C(net286),
    .D(_02432_),
    .Y(_02453_));
 sky130_fd_sc_hd__o41a_4 _14478_ (.A1(_04747_),
    .A2(net264),
    .A3(_11387_),
    .A4(_02442_),
    .B1(_02421_),
    .X(_02464_));
 sky130_fd_sc_hd__o21ai_4 _14479_ (.A1(net253),
    .A2(_02442_),
    .B1(_02421_),
    .Y(_02475_));
 sky130_fd_sc_hd__o211ai_2 _14480_ (.A1(_11431_),
    .A2(_02442_),
    .B1(net33),
    .C1(_02421_),
    .Y(_02486_));
 sky130_fd_sc_hd__and4b_1 _14481_ (.A_N(net44),
    .B(_04026_),
    .C(net5),
    .D(net33),
    .X(_02497_));
 sky130_fd_sc_hd__or4_4 _14482_ (.A(net44),
    .B(net6),
    .C(_04015_),
    .D(_03286_),
    .X(_02508_));
 sky130_fd_sc_hd__o211ai_4 _14483_ (.A1(_04015_),
    .A2(_04331_),
    .B1(_02399_),
    .C1(_02486_),
    .Y(_02519_));
 sky130_fd_sc_hd__a21oi_4 _14484_ (.A1(_02508_),
    .A2(_02519_),
    .B1(_02388_),
    .Y(_02530_));
 sky130_fd_sc_hd__a21o_1 _14485_ (.A1(_02508_),
    .A2(_02519_),
    .B1(_02388_),
    .X(_02541_));
 sky130_fd_sc_hd__and3_1 _14486_ (.A(_02388_),
    .B(_02508_),
    .C(_02519_),
    .X(_02552_));
 sky130_fd_sc_hd__o211ai_4 _14487_ (.A1(_02366_),
    .A2(_02377_),
    .B1(_02508_),
    .C1(_02519_),
    .Y(_02563_));
 sky130_fd_sc_hd__a21oi_2 _14488_ (.A1(_02541_),
    .A2(_02563_),
    .B1(_02355_),
    .Y(_02574_));
 sky130_fd_sc_hd__o2bb2ai_2 _14489_ (.A1_N(_00723_),
    .A2_N(_02344_),
    .B1(_02530_),
    .B2(_02552_),
    .Y(_02585_));
 sky130_fd_sc_hd__o211ai_4 _14490_ (.A1(_00734_),
    .A2(_00603_),
    .B1(_00723_),
    .C1(_02563_),
    .Y(_02596_));
 sky130_fd_sc_hd__nor2_1 _14491_ (.A(_02530_),
    .B(_02596_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand3_1 _14492_ (.A(_02355_),
    .B(_02541_),
    .C(_02563_),
    .Y(_02618_));
 sky130_fd_sc_hd__a2bb2oi_2 _14493_ (.A1_N(_02530_),
    .A2_N(_02596_),
    .B1(_02311_),
    .B2(_02322_),
    .Y(_02629_));
 sky130_fd_sc_hd__o2bb2ai_2 _14494_ (.A1_N(_02333_),
    .A2_N(_02585_),
    .B1(_02596_),
    .B2(_02530_),
    .Y(_02640_));
 sky130_fd_sc_hd__a21oi_2 _14495_ (.A1(_02585_),
    .A2(_02618_),
    .B1(_02333_),
    .Y(_02650_));
 sky130_fd_sc_hd__o2bb2ai_2 _14496_ (.A1_N(_02311_),
    .A2_N(_02322_),
    .B1(_02574_),
    .B2(_02607_),
    .Y(_02661_));
 sky130_fd_sc_hd__o211a_4 _14497_ (.A1(_02596_),
    .A2(_02530_),
    .B1(_02333_),
    .C1(_02585_),
    .X(_02672_));
 sky130_fd_sc_hd__o211ai_1 _14498_ (.A1(_02596_),
    .A2(_02530_),
    .B1(_02333_),
    .C1(_02585_),
    .Y(_02683_));
 sky130_fd_sc_hd__a21oi_2 _14499_ (.A1(_02661_),
    .A2(_02683_),
    .B1(_02136_),
    .Y(_02694_));
 sky130_fd_sc_hd__o21ai_4 _14500_ (.A1(_02650_),
    .A2(_02672_),
    .B1(_02125_),
    .Y(_02705_));
 sky130_fd_sc_hd__nand2_4 _14501_ (.A(_02136_),
    .B(_02661_),
    .Y(_02716_));
 sky130_fd_sc_hd__nor3_1 _14502_ (.A(_02125_),
    .B(_02650_),
    .C(_02672_),
    .Y(_02727_));
 sky130_fd_sc_hd__o21ai_1 _14503_ (.A1(_02672_),
    .A2(_02716_),
    .B1(_02705_),
    .Y(_02738_));
 sky130_fd_sc_hd__o22ai_2 _14504_ (.A1(_02070_),
    .A2(_02092_),
    .B1(_02694_),
    .B2(_02727_),
    .Y(_02749_));
 sky130_fd_sc_hd__o2111ai_4 _14505_ (.A1(_02672_),
    .A2(_02716_),
    .B1(_02705_),
    .C1(_02081_),
    .D1(_02103_),
    .Y(_02760_));
 sky130_fd_sc_hd__o21bai_1 _14506_ (.A1(_02694_),
    .A2(_02727_),
    .B1_N(_02114_),
    .Y(_02771_));
 sky130_fd_sc_hd__o221ai_4 _14507_ (.A1(_02070_),
    .A2(_02092_),
    .B1(_02672_),
    .B2(_02716_),
    .C1(_02705_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand3_4 _14508_ (.A(_02771_),
    .B(_02782_),
    .C(_01884_),
    .Y(_02793_));
 sky130_fd_sc_hd__a22oi_2 _14509_ (.A1(_00899_),
    .A2(_01227_),
    .B1(_02114_),
    .B2(_02738_),
    .Y(_02804_));
 sky130_fd_sc_hd__o211ai_4 _14510_ (.A1(_00888_),
    .A2(_01216_),
    .B1(_02749_),
    .C1(_02760_),
    .Y(_02815_));
 sky130_fd_sc_hd__o211ai_1 _14511_ (.A1(_12768_),
    .A2(_12801_),
    .B1(_12834_),
    .C1(_01118_),
    .Y(_02826_));
 sky130_fd_sc_hd__a22o_1 _14512_ (.A1(_12812_),
    .A2(_12834_),
    .B1(_01063_),
    .B2(_01085_),
    .X(_02837_));
 sky130_fd_sc_hd__nand2_1 _14513_ (.A(_01107_),
    .B(_02826_),
    .Y(_02848_));
 sky130_fd_sc_hd__nor2_8 _14514_ (.A(net37),
    .B(_04037_),
    .Y(_02858_));
 sky130_fd_sc_hd__or2_4 _14515_ (.A(net37),
    .B(_04037_),
    .X(_02869_));
 sky130_fd_sc_hd__and2_4 _14516_ (.A(_04037_),
    .B(net37),
    .X(_02880_));
 sky130_fd_sc_hd__nand2_8 _14517_ (.A(_04037_),
    .B(net37),
    .Y(_02891_));
 sky130_fd_sc_hd__o21a_1 _14518_ (.A1(_02858_),
    .A2(_02880_),
    .B1(net1),
    .X(_02902_));
 sky130_fd_sc_hd__o2bb2a_1 _14519_ (.A1_N(net12),
    .A2_N(_01315_),
    .B1(_01304_),
    .B2(_04528_),
    .X(_02913_));
 sky130_fd_sc_hd__or3_1 _14520_ (.A(_12341_),
    .B(_04441_),
    .C(_04408_),
    .X(_02924_));
 sky130_fd_sc_hd__or3_1 _14521_ (.A(net36),
    .B(_03993_),
    .C(_03396_),
    .X(_02935_));
 sky130_fd_sc_hd__a21oi_2 _14522_ (.A1(_02924_),
    .A2(_02935_),
    .B1(_02913_),
    .Y(_02946_));
 sky130_fd_sc_hd__o311a_1 _14523_ (.A1(_03396_),
    .A2(_03993_),
    .A3(net36),
    .B1(_02924_),
    .C1(_02913_),
    .X(_02957_));
 sky130_fd_sc_hd__o221ai_2 _14524_ (.A1(_04474_),
    .A2(_12341_),
    .B1(_12363_),
    .B2(_03396_),
    .C1(_02913_),
    .Y(_02968_));
 sky130_fd_sc_hd__a2111oi_1 _14525_ (.A1(_02869_),
    .A2(_02891_),
    .B1(_03176_),
    .C1(_02946_),
    .D1(_02957_),
    .Y(_02979_));
 sky130_fd_sc_hd__o221a_1 _14526_ (.A1(_02858_),
    .A2(_02880_),
    .B1(_02946_),
    .B2(_02957_),
    .C1(net1),
    .X(_02990_));
 sky130_fd_sc_hd__nor3_1 _14527_ (.A(_02902_),
    .B(_02946_),
    .C(_02957_),
    .Y(_03001_));
 sky130_fd_sc_hd__nor2_1 _14528_ (.A(_02990_),
    .B(_03001_),
    .Y(_03012_));
 sky130_fd_sc_hd__a32o_1 _14529_ (.A1(_11771_),
    .A2(net267),
    .A3(net315),
    .B1(net26),
    .B2(_11793_),
    .X(_03023_));
 sky130_fd_sc_hd__or3b_1 _14530_ (.A(_03616_),
    .B(net34),
    .C_N(net64),
    .X(_03033_));
 sky130_fd_sc_hd__nand3_2 _14531_ (.A(_04998_),
    .B(net304),
    .C(_10313_),
    .Y(_03044_));
 sky130_fd_sc_hd__or3b_2 _14532_ (.A(_03725_),
    .B(net64),
    .C_N(net63),
    .X(_03055_));
 sky130_fd_sc_hd__o211ai_4 _14533_ (.A1(net267),
    .A2(_05436_),
    .B1(_08250_),
    .C1(_05414_),
    .Y(_03066_));
 sky130_fd_sc_hd__a22oi_2 _14534_ (.A1(_03033_),
    .A2(_03044_),
    .B1(_03055_),
    .B2(_03066_),
    .Y(_03077_));
 sky130_fd_sc_hd__a22o_1 _14535_ (.A1(_03033_),
    .A2(_03044_),
    .B1(_03055_),
    .B2(_03066_),
    .X(_03088_));
 sky130_fd_sc_hd__o2111a_1 _14536_ (.A1(_03616_),
    .A2(_10346_),
    .B1(_03044_),
    .C1(_03055_),
    .D1(_03066_),
    .X(_03099_));
 sky130_fd_sc_hd__o2111ai_2 _14537_ (.A1(_03616_),
    .A2(_10346_),
    .B1(_03044_),
    .C1(_03055_),
    .D1(_03066_),
    .Y(_03110_));
 sky130_fd_sc_hd__o21ai_1 _14538_ (.A1(_03077_),
    .A2(_03099_),
    .B1(_03023_),
    .Y(_03121_));
 sky130_fd_sc_hd__nand3b_1 _14539_ (.A_N(_03023_),
    .B(_03088_),
    .C(_03110_),
    .Y(_03132_));
 sky130_fd_sc_hd__a22oi_1 _14540_ (.A1(_01447_),
    .A2(_01480_),
    .B1(_03121_),
    .B2(_03132_),
    .Y(_03143_));
 sky130_fd_sc_hd__a22o_1 _14541_ (.A1(_01447_),
    .A2(_01480_),
    .B1(_03121_),
    .B2(_03132_),
    .X(_03154_));
 sky130_fd_sc_hd__and4_1 _14542_ (.A(_01447_),
    .B(_01480_),
    .C(_03121_),
    .D(_03132_),
    .X(_03165_));
 sky130_fd_sc_hd__nand4_1 _14543_ (.A(_01447_),
    .B(_01480_),
    .C(_03121_),
    .D(_03132_),
    .Y(_03177_));
 sky130_fd_sc_hd__o22ai_2 _14544_ (.A1(_02990_),
    .A2(_03001_),
    .B1(_03143_),
    .B2(_03165_),
    .Y(_03188_));
 sky130_fd_sc_hd__nand3_2 _14545_ (.A(_03012_),
    .B(_03154_),
    .C(_03177_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_4 _14546_ (.A1(_03188_),
    .A2(_03199_),
    .B1(_02848_),
    .Y(_03209_));
 sky130_fd_sc_hd__o2111a_2 _14547_ (.A1(_01063_),
    .A2(_01085_),
    .B1(_02837_),
    .C1(_03188_),
    .D1(_03199_),
    .X(_03220_));
 sky130_fd_sc_hd__a31o_1 _14548_ (.A1(_01359_),
    .A2(_01370_),
    .A3(_01523_),
    .B1(_01534_),
    .X(_03231_));
 sky130_fd_sc_hd__a21oi_1 _14549_ (.A1(_01523_),
    .A2(_01392_),
    .B1(_01534_),
    .Y(_03242_));
 sky130_fd_sc_hd__o21a_1 _14550_ (.A1(_03209_),
    .A2(_03220_),
    .B1(_03231_),
    .X(_03253_));
 sky130_fd_sc_hd__o21ai_1 _14551_ (.A1(_03209_),
    .A2(_03220_),
    .B1(_03231_),
    .Y(_03264_));
 sky130_fd_sc_hd__a2111oi_2 _14552_ (.A1(_01392_),
    .A2(_01523_),
    .B1(_01534_),
    .C1(_03209_),
    .D1(_03220_),
    .Y(_03275_));
 sky130_fd_sc_hd__or3_1 _14553_ (.A(_03209_),
    .B(_03220_),
    .C(_03231_),
    .X(_03287_));
 sky130_fd_sc_hd__o21a_1 _14554_ (.A1(_03209_),
    .A2(_03220_),
    .B1(_03242_),
    .X(_03298_));
 sky130_fd_sc_hd__nor3_2 _14555_ (.A(_03209_),
    .B(_03242_),
    .C(_03220_),
    .Y(_03309_));
 sky130_fd_sc_hd__nor2_1 _14556_ (.A(_03298_),
    .B(_03309_),
    .Y(_03320_));
 sky130_fd_sc_hd__a211o_1 _14557_ (.A1(_02793_),
    .A2(_02815_),
    .B1(_03253_),
    .C1(_03275_),
    .X(_03331_));
 sky130_fd_sc_hd__o211ai_2 _14558_ (.A1(_03253_),
    .A2(_03275_),
    .B1(_02793_),
    .C1(_02815_),
    .Y(_03342_));
 sky130_fd_sc_hd__o211a_1 _14559_ (.A1(_03298_),
    .A2(_03309_),
    .B1(_02793_),
    .C1(_02815_),
    .X(_03353_));
 sky130_fd_sc_hd__o211ai_2 _14560_ (.A1(_03298_),
    .A2(_03309_),
    .B1(_02793_),
    .C1(_02815_),
    .Y(_03363_));
 sky130_fd_sc_hd__a22oi_2 _14561_ (.A1(_02793_),
    .A2(_02815_),
    .B1(_03264_),
    .B2(_03287_),
    .Y(_03374_));
 sky130_fd_sc_hd__a22o_1 _14562_ (.A1(_02793_),
    .A2(_02815_),
    .B1(_03264_),
    .B2(_03287_),
    .X(_03385_));
 sky130_fd_sc_hd__nand3_2 _14563_ (.A(_03385_),
    .B(_01862_),
    .C(_03363_),
    .Y(_03397_));
 sky130_fd_sc_hd__o21a_1 _14564_ (.A1(_03353_),
    .A2(_03374_),
    .B1(_01873_),
    .X(_03408_));
 sky130_fd_sc_hd__o21ai_2 _14565_ (.A1(_03353_),
    .A2(_03374_),
    .B1(_01873_),
    .Y(_03419_));
 sky130_fd_sc_hd__o21ai_4 _14566_ (.A1(_01600_),
    .A2(_01567_),
    .B1(_01589_),
    .Y(_03430_));
 sky130_fd_sc_hd__inv_2 _14567_ (.A(_03430_),
    .Y(_03441_));
 sky130_fd_sc_hd__o2111ai_4 _14568_ (.A1(_01293_),
    .A2(_01315_),
    .B1(net1),
    .C1(_01348_),
    .D1(_03430_),
    .Y(_03452_));
 sky130_fd_sc_hd__a21o_1 _14569_ (.A1(_01337_),
    .A2(_01348_),
    .B1(_03430_),
    .X(_03463_));
 sky130_fd_sc_hd__and2_1 _14570_ (.A(_03452_),
    .B(_03463_),
    .X(_03474_));
 sky130_fd_sc_hd__nand2_1 _14571_ (.A(_03452_),
    .B(_03463_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand4_2 _14572_ (.A(_03397_),
    .B(_03419_),
    .C(_03452_),
    .D(_03463_),
    .Y(_03495_));
 sky130_fd_sc_hd__a22o_1 _14573_ (.A1(_03397_),
    .A2(_03419_),
    .B1(_03452_),
    .B2(_03463_),
    .X(_03507_));
 sky130_fd_sc_hd__a21o_1 _14574_ (.A1(_03397_),
    .A2(_03419_),
    .B1(_03485_),
    .X(_03518_));
 sky130_fd_sc_hd__nand3_1 _14575_ (.A(_03397_),
    .B(_03419_),
    .C(_03485_),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_1 _14576_ (.A(_01688_),
    .B(_01699_),
    .Y(_03540_));
 sky130_fd_sc_hd__nand4_2 _14577_ (.A(_01688_),
    .B(_01699_),
    .C(_03518_),
    .D(_03529_),
    .Y(_03551_));
 sky130_fd_sc_hd__nand3_2 _14578_ (.A(_03495_),
    .B(_03507_),
    .C(_03540_),
    .Y(_03562_));
 sky130_fd_sc_hd__a21bo_1 _14579_ (.A1(_03551_),
    .A2(_03562_),
    .B1_N(_01753_),
    .X(_03573_));
 sky130_fd_sc_hd__and3b_1 _14580_ (.A_N(_01753_),
    .B(_03551_),
    .C(_03562_),
    .X(_03584_));
 sky130_fd_sc_hd__nand3b_2 _14581_ (.A_N(_01753_),
    .B(_03551_),
    .C(_03562_),
    .Y(_03595_));
 sky130_fd_sc_hd__nand2_2 _14582_ (.A(_03573_),
    .B(_03595_),
    .Y(_03606_));
 sky130_fd_sc_hd__or3_1 _14583_ (.A(_12166_),
    .B(_00231_),
    .C(_01764_),
    .X(_03617_));
 sky130_fd_sc_hd__a31o_1 _14584_ (.A1(_12155_),
    .A2(_00242_),
    .A3(_01775_),
    .B1(_01786_),
    .X(_03628_));
 sky130_fd_sc_hd__o211a_1 _14585_ (.A1(_00286_),
    .A2(_01764_),
    .B1(_01797_),
    .C1(_03606_),
    .X(_03639_));
 sky130_fd_sc_hd__a31o_1 _14586_ (.A1(_03573_),
    .A2(_03595_),
    .A3(_03628_),
    .B1(_03639_),
    .X(_03650_));
 sky130_fd_sc_hd__xor2_1 _14587_ (.A(_01851_),
    .B(_03650_),
    .X(net70));
 sky130_fd_sc_hd__o22ai_4 _14588_ (.A1(_03606_),
    .A2(_03617_),
    .B1(_03650_),
    .B2(_01851_),
    .Y(_03671_));
 sky130_fd_sc_hd__a31oi_2 _14589_ (.A1(_03385_),
    .A2(_01862_),
    .A3(_03363_),
    .B1(_03485_),
    .Y(_03682_));
 sky130_fd_sc_hd__a32oi_4 _14590_ (.A1(_01873_),
    .A2(_03331_),
    .A3(_03342_),
    .B1(_03397_),
    .B2(_03474_),
    .Y(_03693_));
 sky130_fd_sc_hd__and2b_4 _14591_ (.A_N(net38),
    .B(net39),
    .X(_03704_));
 sky130_fd_sc_hd__nand2_8 _14592_ (.A(_04037_),
    .B(net39),
    .Y(_03714_));
 sky130_fd_sc_hd__nor2_4 _14593_ (.A(net39),
    .B(_04037_),
    .Y(_03726_));
 sky130_fd_sc_hd__nand2b_4 _14594_ (.A_N(net39),
    .B(net38),
    .Y(_03737_));
 sky130_fd_sc_hd__a21oi_1 _14595_ (.A1(_03714_),
    .A2(_03737_),
    .B1(_03176_),
    .Y(_03748_));
 sky130_fd_sc_hd__o221a_4 _14596_ (.A1(_02946_),
    .A2(_02979_),
    .B1(net285),
    .B2(_03726_),
    .C1(net1),
    .X(_03759_));
 sky130_fd_sc_hd__a211oi_2 _14597_ (.A1(_02968_),
    .A2(_02902_),
    .B1(_02946_),
    .C1(_03748_),
    .Y(_03770_));
 sky130_fd_sc_hd__or2_1 _14598_ (.A(_03759_),
    .B(_03770_),
    .X(_03781_));
 sky130_fd_sc_hd__o21ba_1 _14599_ (.A1(_03242_),
    .A2(_03220_),
    .B1_N(_03209_),
    .X(_03792_));
 sky130_fd_sc_hd__nor2_2 _14600_ (.A(_03781_),
    .B(_03792_),
    .Y(_03802_));
 sky130_fd_sc_hd__o21a_1 _14601_ (.A1(_03759_),
    .A2(_03770_),
    .B1(_03792_),
    .X(_03813_));
 sky130_fd_sc_hd__nor2_1 _14602_ (.A(_03802_),
    .B(_03813_),
    .Y(_03824_));
 sky130_fd_sc_hd__a21boi_2 _14603_ (.A1(_01895_),
    .A2(_02048_),
    .B1_N(_02059_),
    .Y(_03836_));
 sky130_fd_sc_hd__a21bo_2 _14604_ (.A1(_01895_),
    .A2(_02048_),
    .B1_N(_02059_),
    .X(_03847_));
 sky130_fd_sc_hd__a22o_1 _14605_ (.A1(_04539_),
    .A2(_02858_),
    .B1(_02880_),
    .B2(net12),
    .X(_03858_));
 sky130_fd_sc_hd__a32o_1 _14606_ (.A1(net318),
    .A2(_04452_),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net23),
    .X(_03869_));
 sky130_fd_sc_hd__o32a_1 _14607_ (.A1(_12341_),
    .A2(net306),
    .A3(_04703_),
    .B1(_03506_),
    .B2(_12363_),
    .X(_03879_));
 sky130_fd_sc_hd__a32o_1 _14608_ (.A1(_12330_),
    .A2(net267),
    .A3(net315),
    .B1(net26),
    .B2(_12352_),
    .X(_03890_));
 sky130_fd_sc_hd__nand2_1 _14609_ (.A(_03869_),
    .B(_03890_),
    .Y(_03901_));
 sky130_fd_sc_hd__o221ai_4 _14610_ (.A1(_04474_),
    .A2(_01304_),
    .B1(_01326_),
    .B2(_03396_),
    .C1(_03879_),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _14611_ (.A(_03901_),
    .B(_03910_),
    .Y(_03914_));
 sky130_fd_sc_hd__xnor2_1 _14612_ (.A(_03858_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__xor2_1 _14613_ (.A(_03858_),
    .B(_03914_),
    .X(_03917_));
 sky130_fd_sc_hd__a32o_1 _14614_ (.A1(_04998_),
    .A2(net304),
    .A3(_11771_),
    .B1(_11793_),
    .B2(net27),
    .X(_03918_));
 sky130_fd_sc_hd__or3b_1 _14615_ (.A(_03835_),
    .B(net64),
    .C_N(net63),
    .X(_03919_));
 sky130_fd_sc_hd__nand3_2 _14616_ (.A(_05841_),
    .B(_05863_),
    .C(_08250_),
    .Y(_03920_));
 sky130_fd_sc_hd__or3b_2 _14617_ (.A(_03725_),
    .B(net34),
    .C_N(net64),
    .X(_03921_));
 sky130_fd_sc_hd__o211ai_4 _14618_ (.A1(net267),
    .A2(_05436_),
    .B1(_10313_),
    .C1(_05414_),
    .Y(_03922_));
 sky130_fd_sc_hd__a22oi_2 _14619_ (.A1(_03919_),
    .A2(_03920_),
    .B1(_03921_),
    .B2(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__a22o_1 _14620_ (.A1(_03919_),
    .A2(_03920_),
    .B1(_03921_),
    .B2(_03922_),
    .X(_03924_));
 sky130_fd_sc_hd__and4_1 _14621_ (.A(_03919_),
    .B(_03920_),
    .C(_03921_),
    .D(_03922_),
    .X(_03925_));
 sky130_fd_sc_hd__o2111ai_2 _14622_ (.A1(_03835_),
    .A2(_08283_),
    .B1(_03920_),
    .C1(_03921_),
    .D1(_03922_),
    .Y(_03926_));
 sky130_fd_sc_hd__o21ai_2 _14623_ (.A1(_03923_),
    .A2(_03925_),
    .B1(_03918_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand3b_1 _14624_ (.A_N(_03918_),
    .B(_03924_),
    .C(_03926_),
    .Y(_03929_));
 sky130_fd_sc_hd__a21oi_2 _14625_ (.A1(_03023_),
    .A2(_03110_),
    .B1(_03077_),
    .Y(_03930_));
 sky130_fd_sc_hd__a21o_1 _14626_ (.A1(_03928_),
    .A2(_03929_),
    .B1(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__nand3_2 _14627_ (.A(_03928_),
    .B(_03929_),
    .C(_03930_),
    .Y(_03932_));
 sky130_fd_sc_hd__a21o_1 _14628_ (.A1(_03931_),
    .A2(_03932_),
    .B1(_03917_),
    .X(_03933_));
 sky130_fd_sc_hd__nand3_1 _14629_ (.A(_03917_),
    .B(_03931_),
    .C(_03932_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand3_2 _14630_ (.A(_03915_),
    .B(_03931_),
    .C(_03932_),
    .Y(_03935_));
 sky130_fd_sc_hd__a21o_1 _14631_ (.A1(_03931_),
    .A2(_03932_),
    .B1(_03915_),
    .X(_03936_));
 sky130_fd_sc_hd__a21oi_2 _14632_ (.A1(_03933_),
    .A2(_03934_),
    .B1(_03836_),
    .Y(_03937_));
 sky130_fd_sc_hd__a21oi_2 _14633_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_03847_),
    .Y(_03939_));
 sky130_fd_sc_hd__o21a_1 _14634_ (.A1(_03165_),
    .A2(_03012_),
    .B1(_03154_),
    .X(_03940_));
 sky130_fd_sc_hd__o21ai_2 _14635_ (.A1(_03937_),
    .A2(_03939_),
    .B1(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__a31o_1 _14636_ (.A1(_03847_),
    .A2(_03935_),
    .A3(_03936_),
    .B1(_03940_),
    .X(_03942_));
 sky130_fd_sc_hd__nor2_1 _14637_ (.A(_03939_),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__a31o_1 _14638_ (.A1(_03836_),
    .A2(_03933_),
    .A3(_03934_),
    .B1(_03942_),
    .X(_03944_));
 sky130_fd_sc_hd__o21ai_2 _14639_ (.A1(_03939_),
    .A2(_03942_),
    .B1(_03941_),
    .Y(_03945_));
 sky130_fd_sc_hd__nor2_1 _14640_ (.A(_04015_),
    .B(_04375_),
    .Y(_03946_));
 sky130_fd_sc_hd__a31oi_2 _14641_ (.A1(_00625_),
    .A2(_00657_),
    .A3(_04342_),
    .B1(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__a31o_1 _14642_ (.A1(_00625_),
    .A2(_00657_),
    .A3(_04342_),
    .B1(_03946_),
    .X(_03948_));
 sky130_fd_sc_hd__o211ai_2 _14643_ (.A1(_11431_),
    .A2(_02442_),
    .B1(_04484_),
    .C1(_02421_),
    .Y(_03950_));
 sky130_fd_sc_hd__a41oi_4 _14644_ (.A1(net310),
    .A2(net294),
    .A3(net286),
    .A4(_02432_),
    .B1(_04048_),
    .Y(_03951_));
 sky130_fd_sc_hd__nand2_8 _14645_ (.A(net249),
    .B(net7),
    .Y(_03952_));
 sky130_fd_sc_hd__nor4_4 _14646_ (.A(net4),
    .B(net5),
    .C(net6),
    .D(net7),
    .Y(_03953_));
 sky130_fd_sc_hd__nand3_4 _14647_ (.A(_00635_),
    .B(_04048_),
    .C(_04026_),
    .Y(_03954_));
 sky130_fd_sc_hd__nor2_8 _14648_ (.A(_11387_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__nand4_4 _14649_ (.A(net290),
    .B(_02432_),
    .C(_03982_),
    .D(_04048_),
    .Y(_03956_));
 sky130_fd_sc_hd__nor2_8 _14650_ (.A(net262),
    .B(net244),
    .Y(_03957_));
 sky130_fd_sc_hd__nand3b_4 _14651_ (.A_N(net262),
    .B(net288),
    .C(net284),
    .Y(_03958_));
 sky130_fd_sc_hd__a21oi_4 _14652_ (.A1(_11420_),
    .A2(net282),
    .B1(net247),
    .Y(_03959_));
 sky130_fd_sc_hd__o21ai_4 _14653_ (.A1(_11431_),
    .A2(_03954_),
    .B1(_03952_),
    .Y(_03961_));
 sky130_fd_sc_hd__o211ai_2 _14654_ (.A1(_11431_),
    .A2(_03954_),
    .B1(net33),
    .C1(_03952_),
    .Y(_03962_));
 sky130_fd_sc_hd__o211ai_4 _14655_ (.A1(_04026_),
    .A2(_04331_),
    .B1(_03950_),
    .C1(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__and3_1 _14656_ (.A(net6),
    .B(_04320_),
    .C(_04048_),
    .X(_03964_));
 sky130_fd_sc_hd__or4_2 _14657_ (.A(net44),
    .B(net7),
    .C(_04026_),
    .D(_03286_),
    .X(_03965_));
 sky130_fd_sc_hd__nand2_1 _14658_ (.A(_03948_),
    .B(_03963_),
    .Y(_03966_));
 sky130_fd_sc_hd__o311a_1 _14659_ (.A1(_04026_),
    .A2(net7),
    .A3(_04331_),
    .B1(_03948_),
    .C1(_03963_),
    .X(_03967_));
 sky130_fd_sc_hd__a21o_1 _14660_ (.A1(_03963_),
    .A2(_03965_),
    .B1(_03948_),
    .X(_03968_));
 sky130_fd_sc_hd__nand3_2 _14661_ (.A(_03963_),
    .B(_03965_),
    .C(_03947_),
    .Y(_03969_));
 sky130_fd_sc_hd__a21o_1 _14662_ (.A1(_03963_),
    .A2(_03965_),
    .B1(_03947_),
    .X(_03970_));
 sky130_fd_sc_hd__o31a_1 _14663_ (.A1(_02366_),
    .A2(_02377_),
    .A3(_02497_),
    .B1(_02519_),
    .X(_03972_));
 sky130_fd_sc_hd__a21oi_2 _14664_ (.A1(_02388_),
    .A2(_02519_),
    .B1(_02497_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand3_4 _14665_ (.A(_03969_),
    .B(_03970_),
    .C(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _14666_ (.A(_03968_),
    .B(_03972_),
    .Y(_03975_));
 sky130_fd_sc_hd__o211a_1 _14667_ (.A1(_03964_),
    .A2(_03966_),
    .B1(_03972_),
    .C1(_03968_),
    .X(_03976_));
 sky130_fd_sc_hd__o211ai_2 _14668_ (.A1(_03964_),
    .A2(_03966_),
    .B1(_03972_),
    .C1(_03968_),
    .Y(_03977_));
 sky130_fd_sc_hd__a32o_1 _14669_ (.A1(_09698_),
    .A2(_05227_),
    .A3(net255),
    .B1(_05249_),
    .B2(net2),
    .X(_03978_));
 sky130_fd_sc_hd__o211ai_1 _14670_ (.A1(_11387_),
    .A2(_12988_),
    .B1(net317),
    .C1(net235),
    .Y(_03979_));
 sky130_fd_sc_hd__or3b_1 _14671_ (.A(net58),
    .B(_04004_),
    .C_N(net55),
    .X(_03980_));
 sky130_fd_sc_hd__and3b_1 _14672_ (.A_N(net59),
    .B(net3),
    .C(net58),
    .X(_03981_));
 sky130_fd_sc_hd__o311a_1 _14673_ (.A1(net267),
    .A2(_06508_),
    .A3(_11387_),
    .B1(net305),
    .C1(_11354_),
    .X(_03983_));
 sky130_fd_sc_hd__a31oi_2 _14674_ (.A1(_11354_),
    .A2(_11431_),
    .A3(net305),
    .B1(_03981_),
    .Y(_03984_));
 sky130_fd_sc_hd__o221ai_4 _14675_ (.A1(_04004_),
    .A2(_04660_),
    .B1(_13021_),
    .B2(_04638_),
    .C1(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__o2bb2ai_2 _14676_ (.A1_N(_03979_),
    .A2_N(_03980_),
    .B1(_03981_),
    .B2(_03983_),
    .Y(_03986_));
 sky130_fd_sc_hd__a21boi_2 _14677_ (.A1(_03985_),
    .A2(_03986_),
    .B1_N(_03978_),
    .Y(_03987_));
 sky130_fd_sc_hd__a21bo_1 _14678_ (.A1(_03985_),
    .A2(_03986_),
    .B1_N(_03978_),
    .X(_03988_));
 sky130_fd_sc_hd__and3b_1 _14679_ (.A_N(_03978_),
    .B(_03985_),
    .C(_03986_),
    .X(_03989_));
 sky130_fd_sc_hd__nand3b_2 _14680_ (.A_N(_03978_),
    .B(_03985_),
    .C(_03986_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand2_1 _14681_ (.A(_03988_),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__a21oi_2 _14682_ (.A1(_03974_),
    .A2(_03977_),
    .B1(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__a21o_1 _14683_ (.A1(_03974_),
    .A2(_03977_),
    .B1(_03991_),
    .X(_03994_));
 sky130_fd_sc_hd__a32oi_4 _14684_ (.A1(_03969_),
    .A2(_03970_),
    .A3(_03973_),
    .B1(_03988_),
    .B2(_03990_),
    .Y(_03995_));
 sky130_fd_sc_hd__o211a_1 _14685_ (.A1(_03987_),
    .A2(_03989_),
    .B1(_03974_),
    .C1(_03977_),
    .X(_03996_));
 sky130_fd_sc_hd__o221ai_4 _14686_ (.A1(_03987_),
    .A2(_03989_),
    .B1(_03967_),
    .B2(_03975_),
    .C1(_03974_),
    .Y(_03997_));
 sky130_fd_sc_hd__and3_1 _14687_ (.A(_02640_),
    .B(_03994_),
    .C(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__nand3_4 _14688_ (.A(_02640_),
    .B(_03994_),
    .C(_03997_),
    .Y(_03999_));
 sky130_fd_sc_hd__o22a_1 _14689_ (.A1(_02574_),
    .A2(_02629_),
    .B1(_03992_),
    .B2(_03996_),
    .X(_04000_));
 sky130_fd_sc_hd__o22ai_4 _14690_ (.A1(_02574_),
    .A2(_02629_),
    .B1(_03992_),
    .B2(_03996_),
    .Y(_04001_));
 sky130_fd_sc_hd__a21oi_2 _14691_ (.A1(_01906_),
    .A2(_01993_),
    .B1(_01961_),
    .Y(_04002_));
 sky130_fd_sc_hd__a32o_1 _14692_ (.A1(_06486_),
    .A2(_06530_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net30),
    .X(_04003_));
 sky130_fd_sc_hd__and3_2 _14693_ (.A(_03927_),
    .B(net31),
    .C(net61),
    .X(_04005_));
 sky130_fd_sc_hd__nor3b_2 _14694_ (.A(_06837_),
    .B(_07231_),
    .C_N(net258),
    .Y(_04006_));
 sky130_fd_sc_hd__a31oi_4 _14695_ (.A1(_07242_),
    .A2(net258),
    .A3(net292),
    .B1(_04005_),
    .Y(_04007_));
 sky130_fd_sc_hd__nor2_2 _14696_ (.A(_03949_),
    .B(net298),
    .Y(_04008_));
 sky130_fd_sc_hd__o311a_1 _14697_ (.A1(net267),
    .A2(_06508_),
    .A3(_08656_),
    .B1(net299),
    .C1(_08700_),
    .X(_04009_));
 sky130_fd_sc_hd__a31oi_4 _14698_ (.A1(_08700_),
    .A2(net299),
    .A3(net256),
    .B1(_04008_),
    .Y(_04010_));
 sky130_fd_sc_hd__o22ai_4 _14699_ (.A1(_04005_),
    .A2(_04006_),
    .B1(_04008_),
    .B2(_04009_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand2_1 _14700_ (.A(_04007_),
    .B(_04010_),
    .Y(_04012_));
 sky130_fd_sc_hd__o21ai_1 _14701_ (.A1(_04008_),
    .A2(_04009_),
    .B1(_04007_),
    .Y(_04013_));
 sky130_fd_sc_hd__o21ai_1 _14702_ (.A1(_04005_),
    .A2(_04006_),
    .B1(_04010_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand3b_2 _14703_ (.A_N(_04003_),
    .B(_04013_),
    .C(_04014_),
    .Y(_04016_));
 sky130_fd_sc_hd__and3_1 _14704_ (.A(_04003_),
    .B(_04011_),
    .C(_04012_),
    .X(_04017_));
 sky130_fd_sc_hd__nand3_4 _14705_ (.A(_04003_),
    .B(_04011_),
    .C(_04012_),
    .Y(_04018_));
 sky130_fd_sc_hd__a22oi_4 _14706_ (.A1(_02256_),
    .A2(_02289_),
    .B1(_04016_),
    .B2(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__o21ai_2 _14707_ (.A1(_02234_),
    .A2(_02300_),
    .B1(_04016_),
    .Y(_04020_));
 sky130_fd_sc_hd__o211a_1 _14708_ (.A1(_02234_),
    .A2(_02300_),
    .B1(_04016_),
    .C1(_04018_),
    .X(_04021_));
 sky130_fd_sc_hd__a41o_1 _14709_ (.A1(_02256_),
    .A2(_02289_),
    .A3(_04016_),
    .A4(_04018_),
    .B1(_04002_),
    .X(_04022_));
 sky130_fd_sc_hd__nor2_1 _14710_ (.A(_04019_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__o21ai_2 _14711_ (.A1(_04019_),
    .A2(_04021_),
    .B1(_04002_),
    .Y(_04024_));
 sky130_fd_sc_hd__inv_2 _14712_ (.A(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__o21a_1 _14713_ (.A1(_04019_),
    .A2(_04022_),
    .B1(_04024_),
    .X(_04027_));
 sky130_fd_sc_hd__o21ai_1 _14714_ (.A1(_04019_),
    .A2(_04022_),
    .B1(_04024_),
    .Y(_04028_));
 sky130_fd_sc_hd__o2bb2ai_4 _14715_ (.A1_N(_03999_),
    .A2_N(_04001_),
    .B1(_04023_),
    .B2(_04025_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _14716_ (.A(_04027_),
    .B(_04001_),
    .Y(_04030_));
 sky130_fd_sc_hd__o2111ai_4 _14717_ (.A1(_04019_),
    .A2(_04022_),
    .B1(_04024_),
    .C1(_04001_),
    .D1(_03999_),
    .Y(_04031_));
 sky130_fd_sc_hd__o22ai_4 _14718_ (.A1(_02672_),
    .A2(_02716_),
    .B1(_02114_),
    .B2(_02694_),
    .Y(_04032_));
 sky130_fd_sc_hd__a21oi_4 _14719_ (.A1(_04029_),
    .A2(_04031_),
    .B1(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__a21o_1 _14720_ (.A1(_04029_),
    .A2(_04031_),
    .B1(_04032_),
    .X(_04034_));
 sky130_fd_sc_hd__o211a_1 _14721_ (.A1(_03998_),
    .A2(_04030_),
    .B1(_04029_),
    .C1(_04032_),
    .X(_04035_));
 sky130_fd_sc_hd__o211ai_2 _14722_ (.A1(_03998_),
    .A2(_04030_),
    .B1(_04029_),
    .C1(_04032_),
    .Y(_04036_));
 sky130_fd_sc_hd__o21bai_1 _14723_ (.A1(_04033_),
    .A2(_04035_),
    .B1_N(_03945_),
    .Y(_04038_));
 sky130_fd_sc_hd__nand3_1 _14724_ (.A(_03945_),
    .B(_04034_),
    .C(_04036_),
    .Y(_04039_));
 sky130_fd_sc_hd__o21ai_2 _14725_ (.A1(_04033_),
    .A2(_04035_),
    .B1(_03945_),
    .Y(_04040_));
 sky130_fd_sc_hd__nand3b_2 _14726_ (.A_N(_03945_),
    .B(_04034_),
    .C(_04036_),
    .Y(_04041_));
 sky130_fd_sc_hd__o21ai_2 _14727_ (.A1(_03298_),
    .A2(_03309_),
    .B1(_02815_),
    .Y(_04042_));
 sky130_fd_sc_hd__a22oi_4 _14728_ (.A1(_02804_),
    .A2(_02760_),
    .B1(_02793_),
    .B2(_03320_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand4_4 _14729_ (.A(_02793_),
    .B(_04040_),
    .C(_04041_),
    .D(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__nand3_4 _14730_ (.A(_04038_),
    .B(_04039_),
    .C(_04043_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_1 _14731_ (.A(_04045_),
    .B(_03824_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand3_1 _14732_ (.A(_04044_),
    .B(_04045_),
    .C(_03824_),
    .Y(_04047_));
 sky130_fd_sc_hd__a21o_1 _14733_ (.A1(_04044_),
    .A2(_04045_),
    .B1(_03824_),
    .X(_04049_));
 sky130_fd_sc_hd__o211ai_4 _14734_ (.A1(_03802_),
    .A2(_03813_),
    .B1(_04044_),
    .C1(_04045_),
    .Y(_04050_));
 sky130_fd_sc_hd__a21bo_1 _14735_ (.A1(_04044_),
    .A2(_04045_),
    .B1_N(_03824_),
    .X(_04051_));
 sky130_fd_sc_hd__o211ai_4 _14736_ (.A1(_03408_),
    .A2(_03682_),
    .B1(_04047_),
    .C1(_04049_),
    .Y(_04052_));
 sky130_fd_sc_hd__nand3_2 _14737_ (.A(_04051_),
    .B(_03693_),
    .C(_04050_),
    .Y(_04053_));
 sky130_fd_sc_hd__inv_2 _14738_ (.A(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__nand2_1 _14739_ (.A(_04052_),
    .B(_04053_),
    .Y(_04055_));
 sky130_fd_sc_hd__nand3b_4 _14740_ (.A_N(_03452_),
    .B(_04052_),
    .C(_04053_),
    .Y(_04056_));
 sky130_fd_sc_hd__o2bb2ai_1 _14741_ (.A1_N(_04052_),
    .A2_N(_04053_),
    .B1(_01359_),
    .B2(_03441_),
    .Y(_04057_));
 sky130_fd_sc_hd__and2_1 _14742_ (.A(_04056_),
    .B(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__a21oi_4 _14743_ (.A1(_03452_),
    .A2(_04055_),
    .B1(_03562_),
    .Y(_04060_));
 sky130_fd_sc_hd__o21ai_2 _14744_ (.A1(_03452_),
    .A2(_04055_),
    .B1(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__a32oi_2 _14745_ (.A1(_03495_),
    .A2(_03507_),
    .A3(_03540_),
    .B1(_04056_),
    .B2(_04057_),
    .Y(_04062_));
 sky130_fd_sc_hd__a21oi_2 _14746_ (.A1(_04056_),
    .A2(_04060_),
    .B1(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__a31o_1 _14747_ (.A1(_03573_),
    .A2(_00209_),
    .A3(_01742_),
    .B1(_03584_),
    .X(_04064_));
 sky130_fd_sc_hd__xor2_2 _14748_ (.A(_04063_),
    .B(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__nand2_2 _14749_ (.A(_03671_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__or2_1 _14750_ (.A(_04065_),
    .B(_03671_),
    .X(_04067_));
 sky130_fd_sc_hd__and2_1 _14751_ (.A(_04066_),
    .B(_04067_),
    .X(net71));
 sky130_fd_sc_hd__nand2_1 _14752_ (.A(_03584_),
    .B(_04058_),
    .Y(_04068_));
 sky130_fd_sc_hd__a41o_2 _14753_ (.A1(_02793_),
    .A2(_04040_),
    .A3(_04041_),
    .A4(_04042_),
    .B1(_03824_),
    .X(_04070_));
 sky130_fd_sc_hd__nand2_1 _14754_ (.A(_04044_),
    .B(_04046_),
    .Y(_04071_));
 sky130_fd_sc_hd__a32oi_4 _14755_ (.A1(_04029_),
    .A2(_04031_),
    .A3(_04032_),
    .B1(_03944_),
    .B2(_03941_),
    .Y(_04072_));
 sky130_fd_sc_hd__o21ai_2 _14756_ (.A1(_03945_),
    .A2(_04033_),
    .B1(_04036_),
    .Y(_04073_));
 sky130_fd_sc_hd__o22a_1 _14757_ (.A1(_05457_),
    .A2(_11782_),
    .B1(_11804_),
    .B2(_03725_),
    .X(_04074_));
 sky130_fd_sc_hd__a32o_1 _14758_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_11771_),
    .B1(_11793_),
    .B2(net28),
    .X(_04075_));
 sky130_fd_sc_hd__or3b_1 _14759_ (.A(_03835_),
    .B(net34),
    .C_N(net64),
    .X(_04076_));
 sky130_fd_sc_hd__nand3_2 _14760_ (.A(_05841_),
    .B(_05863_),
    .C(_10313_),
    .Y(_04077_));
 sky130_fd_sc_hd__or3b_2 _14761_ (.A(_03916_),
    .B(net64),
    .C_N(net63),
    .X(_04078_));
 sky130_fd_sc_hd__o211ai_4 _14762_ (.A1(net267),
    .A2(_06508_),
    .B1(_08250_),
    .C1(_06486_),
    .Y(_04079_));
 sky130_fd_sc_hd__a22oi_2 _14763_ (.A1(_04076_),
    .A2(_04077_),
    .B1(_04078_),
    .B2(_04079_),
    .Y(_04081_));
 sky130_fd_sc_hd__a22o_1 _14764_ (.A1(_04076_),
    .A2(_04077_),
    .B1(_04078_),
    .B2(_04079_),
    .X(_04082_));
 sky130_fd_sc_hd__o2111a_1 _14765_ (.A1(_03835_),
    .A2(_10346_),
    .B1(_04077_),
    .C1(_04078_),
    .D1(_04079_),
    .X(_04083_));
 sky130_fd_sc_hd__o2111ai_2 _14766_ (.A1(_03835_),
    .A2(_10346_),
    .B1(_04077_),
    .C1(_04078_),
    .D1(_04079_),
    .Y(_04084_));
 sky130_fd_sc_hd__o21ai_1 _14767_ (.A1(_04081_),
    .A2(_04083_),
    .B1(_04075_),
    .Y(_04085_));
 sky130_fd_sc_hd__nand3_1 _14768_ (.A(_04082_),
    .B(_04084_),
    .C(_04074_),
    .Y(_04086_));
 sky130_fd_sc_hd__o21ai_1 _14769_ (.A1(_04081_),
    .A2(_04083_),
    .B1(_04074_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand3_1 _14770_ (.A(_04075_),
    .B(_04082_),
    .C(_04084_),
    .Y(_04088_));
 sky130_fd_sc_hd__a21o_1 _14771_ (.A1(_03918_),
    .A2(_03926_),
    .B1(_03923_),
    .X(_04089_));
 sky130_fd_sc_hd__a21oi_1 _14772_ (.A1(_03918_),
    .A2(_03926_),
    .B1(_03923_),
    .Y(_04090_));
 sky130_fd_sc_hd__and3_1 _14773_ (.A(_04089_),
    .B(_04088_),
    .C(_04087_),
    .X(_04092_));
 sky130_fd_sc_hd__nand3_2 _14774_ (.A(_04089_),
    .B(_04088_),
    .C(_04087_),
    .Y(_04093_));
 sky130_fd_sc_hd__and3_1 _14775_ (.A(_04085_),
    .B(_04086_),
    .C(_04090_),
    .X(_04094_));
 sky130_fd_sc_hd__nand3_2 _14776_ (.A(_04085_),
    .B(_04086_),
    .C(_04090_),
    .Y(_04095_));
 sky130_fd_sc_hd__a32o_1 _14777_ (.A1(net318),
    .A2(_04452_),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net23),
    .X(_04096_));
 sky130_fd_sc_hd__or3_1 _14778_ (.A(net36),
    .B(_03993_),
    .C(_03616_),
    .X(_04097_));
 sky130_fd_sc_hd__nand4_1 _14779_ (.A(_03993_),
    .B(net304),
    .C(net36),
    .D(_04998_),
    .Y(_04098_));
 sky130_fd_sc_hd__o32a_1 _14780_ (.A1(_01304_),
    .A2(net306),
    .A3(_04703_),
    .B1(_03506_),
    .B2(_01326_),
    .X(_04099_));
 sky130_fd_sc_hd__a21oi_1 _14781_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__a21o_1 _14782_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_04099_),
    .X(_04101_));
 sky130_fd_sc_hd__o221ai_4 _14783_ (.A1(_05020_),
    .A2(_12341_),
    .B1(_12363_),
    .B2(_03616_),
    .C1(_04099_),
    .Y(_04103_));
 sky130_fd_sc_hd__nand3_2 _14784_ (.A(_04096_),
    .B(_04101_),
    .C(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__a21o_1 _14785_ (.A1(_04101_),
    .A2(_04103_),
    .B1(_04096_),
    .X(_04105_));
 sky130_fd_sc_hd__nand2_1 _14786_ (.A(_04104_),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a21oi_1 _14787_ (.A1(_04093_),
    .A2(_04095_),
    .B1(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__nand3_1 _14788_ (.A(_04093_),
    .B(_04095_),
    .C(_04106_),
    .Y(_04108_));
 sky130_fd_sc_hd__a22o_1 _14789_ (.A1(_04093_),
    .A2(_04095_),
    .B1(_04104_),
    .B2(_04105_),
    .X(_04109_));
 sky130_fd_sc_hd__nand4_2 _14790_ (.A(_04093_),
    .B(_04095_),
    .C(_04104_),
    .D(_04105_),
    .Y(_04110_));
 sky130_fd_sc_hd__o22a_1 _14791_ (.A1(_04020_),
    .A2(_04017_),
    .B1(_04002_),
    .B2(_04019_),
    .X(_04111_));
 sky130_fd_sc_hd__o22ai_4 _14792_ (.A1(_04020_),
    .A2(_04017_),
    .B1(_04002_),
    .B2(_04019_),
    .Y(_04112_));
 sky130_fd_sc_hd__a21oi_2 _14793_ (.A1(_04109_),
    .A2(_04110_),
    .B1(_04112_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand3b_1 _14794_ (.A_N(_04107_),
    .B(_04111_),
    .C(_04108_),
    .Y(_04115_));
 sky130_fd_sc_hd__nand3_2 _14795_ (.A(_04109_),
    .B(_04110_),
    .C(_04112_),
    .Y(_04116_));
 sky130_fd_sc_hd__a21bo_1 _14796_ (.A1(_03915_),
    .A2(_03932_),
    .B1_N(_03931_),
    .X(_04117_));
 sky130_fd_sc_hd__a32o_1 _14797_ (.A1(_03928_),
    .A2(_03929_),
    .A3(_03930_),
    .B1(_03931_),
    .B2(_03917_),
    .X(_04118_));
 sky130_fd_sc_hd__a21oi_1 _14798_ (.A1(_04115_),
    .A2(_04116_),
    .B1(_04117_),
    .Y(_04119_));
 sky130_fd_sc_hd__and3_1 _14799_ (.A(_04115_),
    .B(_04116_),
    .C(_04117_),
    .X(_04120_));
 sky130_fd_sc_hd__nor2_1 _14800_ (.A(_04119_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__a21boi_1 _14801_ (.A1(_04027_),
    .A2(_04001_),
    .B1_N(_03999_),
    .Y(_04122_));
 sky130_fd_sc_hd__o21ai_2 _14802_ (.A1(_04028_),
    .A2(_04000_),
    .B1(_03999_),
    .Y(_04123_));
 sky130_fd_sc_hd__o2bb2ai_2 _14803_ (.A1_N(_03991_),
    .A2_N(_03974_),
    .B1(_03967_),
    .B2(_03975_),
    .Y(_04125_));
 sky130_fd_sc_hd__o21ai_1 _14804_ (.A1(_03964_),
    .A2(_03948_),
    .B1(_03963_),
    .Y(_04126_));
 sky130_fd_sc_hd__o21a_1 _14805_ (.A1(_03964_),
    .A2(_03948_),
    .B1(_03963_),
    .X(_04127_));
 sky130_fd_sc_hd__a32o_1 _14806_ (.A1(_02421_),
    .A2(net249),
    .A3(_04342_),
    .B1(_04364_),
    .B2(net6),
    .X(_04128_));
 sky130_fd_sc_hd__o211ai_2 _14807_ (.A1(_11431_),
    .A2(_03954_),
    .B1(_04484_),
    .C1(_03952_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand4b_4 _14808_ (.A_N(_11409_),
    .B(_04059_),
    .C(net308),
    .D(_03953_),
    .Y(_04130_));
 sky130_fd_sc_hd__o21a_1 _14809_ (.A1(net262),
    .A2(net244),
    .B1(net8),
    .X(_04131_));
 sky130_fd_sc_hd__o21ai_4 _14810_ (.A1(net262),
    .A2(net245),
    .B1(net8),
    .Y(_04132_));
 sky130_fd_sc_hd__nand2_4 _14811_ (.A(net230),
    .B(net228),
    .Y(_04133_));
 sky130_fd_sc_hd__nand3_1 _14812_ (.A(_04132_),
    .B(net33),
    .C(_04130_),
    .Y(_04134_));
 sky130_fd_sc_hd__and4b_1 _14813_ (.A_N(net44),
    .B(_04059_),
    .C(net7),
    .D(net33),
    .X(_04136_));
 sky130_fd_sc_hd__or4_2 _14814_ (.A(net44),
    .B(net8),
    .C(_04048_),
    .D(_03286_),
    .X(_04137_));
 sky130_fd_sc_hd__o311a_2 _14815_ (.A1(_03286_),
    .A2(_04048_),
    .A3(net44),
    .B1(_04134_),
    .C1(_04129_),
    .X(_04138_));
 sky130_fd_sc_hd__o211ai_2 _14816_ (.A1(_04048_),
    .A2(_04331_),
    .B1(_04129_),
    .C1(_04134_),
    .Y(_04139_));
 sky130_fd_sc_hd__a21o_1 _14817_ (.A1(_04137_),
    .A2(_04139_),
    .B1(_04128_),
    .X(_04140_));
 sky130_fd_sc_hd__nand2_1 _14818_ (.A(_04128_),
    .B(_04137_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand3b_2 _14819_ (.A_N(_04128_),
    .B(_04137_),
    .C(_04139_),
    .Y(_04142_));
 sky130_fd_sc_hd__o21ai_2 _14820_ (.A1(_04136_),
    .A2(_04138_),
    .B1(_04128_),
    .Y(_04143_));
 sky130_fd_sc_hd__nand3_4 _14821_ (.A(_04143_),
    .B(_04126_),
    .C(_04142_),
    .Y(_04144_));
 sky130_fd_sc_hd__inv_2 _14822_ (.A(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__a22oi_1 _14823_ (.A1(_03965_),
    .A2(_03966_),
    .B1(_04142_),
    .B2(_04143_),
    .Y(_04147_));
 sky130_fd_sc_hd__o211ai_4 _14824_ (.A1(_04141_),
    .A2(_04138_),
    .B1(_04127_),
    .C1(_04140_),
    .Y(_04148_));
 sky130_fd_sc_hd__o32a_1 _14825_ (.A1(_11420_),
    .A2(_05238_),
    .A3(_11343_),
    .B1(_05260_),
    .B2(_03982_),
    .X(_04149_));
 sky130_fd_sc_hd__a32o_1 _14826_ (.A1(_11354_),
    .A2(_11431_),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net3),
    .X(_04150_));
 sky130_fd_sc_hd__o211ai_4 _14827_ (.A1(_11431_),
    .A2(_00646_),
    .B1(net317),
    .C1(_00625_),
    .Y(_04151_));
 sky130_fd_sc_hd__or3b_2 _14828_ (.A(net58),
    .B(_04015_),
    .C_N(net55),
    .X(_04152_));
 sky130_fd_sc_hd__and3b_1 _14829_ (.A_N(net59),
    .B(net4),
    .C(net58),
    .X(_04153_));
 sky130_fd_sc_hd__a31oi_4 _14830_ (.A1(net235),
    .A2(_12999_),
    .A3(net305),
    .B1(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__o221ai_4 _14831_ (.A1(_04015_),
    .A2(_04660_),
    .B1(_00668_),
    .B2(_04638_),
    .C1(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__a21o_2 _14832_ (.A1(_04151_),
    .A2(_04152_),
    .B1(_04154_),
    .X(_04156_));
 sky130_fd_sc_hd__a21oi_2 _14833_ (.A1(_04155_),
    .A2(_04156_),
    .B1(_04150_),
    .Y(_04158_));
 sky130_fd_sc_hd__a21o_1 _14834_ (.A1(_04155_),
    .A2(_04156_),
    .B1(_04150_),
    .X(_04159_));
 sky130_fd_sc_hd__and3_1 _14835_ (.A(_04150_),
    .B(_04155_),
    .C(_04156_),
    .X(_04160_));
 sky130_fd_sc_hd__nand3_1 _14836_ (.A(_04150_),
    .B(_04155_),
    .C(_04156_),
    .Y(_04161_));
 sky130_fd_sc_hd__o2bb2ai_4 _14837_ (.A1_N(_04144_),
    .A2_N(_04148_),
    .B1(_04158_),
    .B2(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__nand4_4 _14838_ (.A(_04144_),
    .B(_04148_),
    .C(_04159_),
    .D(_04161_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_2 _14839_ (.A1(_04162_),
    .A2(_04163_),
    .B1(_04125_),
    .Y(_04164_));
 sky130_fd_sc_hd__a21o_2 _14840_ (.A1(_04162_),
    .A2(_04163_),
    .B1(_04125_),
    .X(_04165_));
 sky130_fd_sc_hd__o211a_1 _14841_ (.A1(_03976_),
    .A2(_03995_),
    .B1(_04162_),
    .C1(_04163_),
    .X(_04166_));
 sky130_fd_sc_hd__o211ai_4 _14842_ (.A1(_03976_),
    .A2(_03995_),
    .B1(_04162_),
    .C1(_04163_),
    .Y(_04167_));
 sky130_fd_sc_hd__o21ai_2 _14843_ (.A1(_04007_),
    .A2(_04010_),
    .B1(_04018_),
    .Y(_04169_));
 sky130_fd_sc_hd__nand2_1 _14844_ (.A(_03978_),
    .B(_03985_),
    .Y(_04170_));
 sky130_fd_sc_hd__a21boi_2 _14845_ (.A1(_03978_),
    .A2(_03985_),
    .B1_N(_03986_),
    .Y(_04171_));
 sky130_fd_sc_hd__and3_1 _14846_ (.A(_07242_),
    .B(_07253_),
    .C(_07658_),
    .X(_04172_));
 sky130_fd_sc_hd__nor2_1 _14847_ (.A(_03938_),
    .B(_07691_),
    .Y(_04173_));
 sky130_fd_sc_hd__a31o_1 _14848_ (.A1(_07242_),
    .A2(_07253_),
    .A3(_07658_),
    .B1(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__or3b_1 _14849_ (.A(net61),
    .B(_03960_),
    .C_N(net60),
    .X(_04175_));
 sky130_fd_sc_hd__o211ai_4 _14850_ (.A1(_06530_),
    .A2(_09665_),
    .B1(net299),
    .C1(_09698_),
    .Y(_04176_));
 sky130_fd_sc_hd__and3_1 _14851_ (.A(_03927_),
    .B(net32),
    .C(net61),
    .X(_04177_));
 sky130_fd_sc_hd__o311a_1 _14852_ (.A1(net267),
    .A2(_06508_),
    .A3(_08656_),
    .B1(net292),
    .C1(_08700_),
    .X(_04178_));
 sky130_fd_sc_hd__a31oi_2 _14853_ (.A1(_08700_),
    .A2(net292),
    .A3(net256),
    .B1(_04177_),
    .Y(_04180_));
 sky130_fd_sc_hd__o211ai_4 _14854_ (.A1(_03960_),
    .A2(net298),
    .B1(_04176_),
    .C1(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__o2bb2ai_2 _14855_ (.A1_N(_04175_),
    .A2_N(_04176_),
    .B1(_04177_),
    .B2(_04178_),
    .Y(_04182_));
 sky130_fd_sc_hd__o211a_1 _14856_ (.A1(_04172_),
    .A2(_04173_),
    .B1(_04181_),
    .C1(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__o211ai_2 _14857_ (.A1(_04172_),
    .A2(_04173_),
    .B1(_04181_),
    .C1(_04182_),
    .Y(_04184_));
 sky130_fd_sc_hd__a21oi_2 _14858_ (.A1(_04181_),
    .A2(_04182_),
    .B1(_04174_),
    .Y(_04185_));
 sky130_fd_sc_hd__a21o_1 _14859_ (.A1(_04181_),
    .A2(_04182_),
    .B1(_04174_),
    .X(_04186_));
 sky130_fd_sc_hd__a21o_1 _14860_ (.A1(_03986_),
    .A2(_04170_),
    .B1(_04185_),
    .X(_04187_));
 sky130_fd_sc_hd__nand3b_4 _14861_ (.A_N(_04171_),
    .B(_04184_),
    .C(_04186_),
    .Y(_04188_));
 sky130_fd_sc_hd__o21ai_4 _14862_ (.A1(_04183_),
    .A2(_04185_),
    .B1(_04171_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand3_2 _14863_ (.A(_04169_),
    .B(_04188_),
    .C(_04189_),
    .Y(_04191_));
 sky130_fd_sc_hd__a21o_1 _14864_ (.A1(_04188_),
    .A2(_04189_),
    .B1(_04169_),
    .X(_04192_));
 sky130_fd_sc_hd__a22o_1 _14865_ (.A1(_04011_),
    .A2(_04018_),
    .B1(_04188_),
    .B2(_04189_),
    .X(_04193_));
 sky130_fd_sc_hd__o2111ai_4 _14866_ (.A1(_04007_),
    .A2(_04010_),
    .B1(_04018_),
    .C1(_04188_),
    .D1(_04189_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _14867_ (.A(_04193_),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _14868_ (.A(_04191_),
    .B(_04192_),
    .Y(_04196_));
 sky130_fd_sc_hd__o21ai_2 _14869_ (.A1(_04164_),
    .A2(_04166_),
    .B1(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__a21o_1 _14870_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04164_),
    .X(_04198_));
 sky130_fd_sc_hd__nand4_4 _14871_ (.A(_04165_),
    .B(_04167_),
    .C(_04191_),
    .D(_04192_),
    .Y(_04199_));
 sky130_fd_sc_hd__o21ai_1 _14872_ (.A1(_04164_),
    .A2(_04166_),
    .B1(_04195_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand4_2 _14873_ (.A(_04165_),
    .B(_04167_),
    .C(_04193_),
    .D(_04194_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21oi_4 _14874_ (.A1(_04197_),
    .A2(_04199_),
    .B1(_04123_),
    .Y(_04203_));
 sky130_fd_sc_hd__nand3_2 _14875_ (.A(_04122_),
    .B(_04200_),
    .C(_04202_),
    .Y(_04204_));
 sky130_fd_sc_hd__a21oi_2 _14876_ (.A1(_04200_),
    .A2(_04202_),
    .B1(_04122_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand3_4 _14877_ (.A(_04123_),
    .B(_04197_),
    .C(_04199_),
    .Y(_04206_));
 sky130_fd_sc_hd__o211ai_2 _14878_ (.A1(_04119_),
    .A2(_04120_),
    .B1(_04204_),
    .C1(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__o21ai_2 _14879_ (.A1(_04203_),
    .A2(_04205_),
    .B1(_04121_),
    .Y(_04208_));
 sky130_fd_sc_hd__a21o_1 _14880_ (.A1(_04204_),
    .A2(_04206_),
    .B1(_04121_),
    .X(_04209_));
 sky130_fd_sc_hd__nand2_2 _14881_ (.A(_04204_),
    .B(_04121_),
    .Y(_04210_));
 sky130_fd_sc_hd__o211ai_4 _14882_ (.A1(_04033_),
    .A2(_04072_),
    .B1(_04207_),
    .C1(_04208_),
    .Y(_04211_));
 sky130_fd_sc_hd__o211ai_4 _14883_ (.A1(_04205_),
    .A2(_04210_),
    .B1(_04073_),
    .C1(_04209_),
    .Y(_04213_));
 sky130_fd_sc_hd__o21ba_1 _14884_ (.A1(_03940_),
    .A2(_03939_),
    .B1_N(_03937_),
    .X(_04214_));
 sky130_fd_sc_hd__and2b_4 _14885_ (.A_N(net39),
    .B(net40),
    .X(_04215_));
 sky130_fd_sc_hd__nand2b_4 _14886_ (.A_N(net39),
    .B(net40),
    .Y(_04216_));
 sky130_fd_sc_hd__and2b_4 _14887_ (.A_N(net40),
    .B(net39),
    .X(_04217_));
 sky130_fd_sc_hd__nand2b_4 _14888_ (.A_N(net40),
    .B(net39),
    .Y(_04218_));
 sky130_fd_sc_hd__a21oi_1 _14889_ (.A1(_04216_),
    .A2(_04218_),
    .B1(_03176_),
    .Y(_04219_));
 sky130_fd_sc_hd__a22o_1 _14890_ (.A1(net12),
    .A2(_03726_),
    .B1(_04539_),
    .B2(net285),
    .X(_04220_));
 sky130_fd_sc_hd__nand2_1 _14891_ (.A(_04220_),
    .B(_04219_),
    .Y(_04221_));
 sky130_fd_sc_hd__a221o_1 _14892_ (.A1(_04539_),
    .A2(net285),
    .B1(_03726_),
    .B2(net12),
    .C1(_04219_),
    .X(_04222_));
 sky130_fd_sc_hd__nand2_1 _14893_ (.A(_04221_),
    .B(_04222_),
    .Y(_04224_));
 sky130_fd_sc_hd__a21boi_2 _14894_ (.A1(_03858_),
    .A2(_03910_),
    .B1_N(_03901_),
    .Y(_04225_));
 sky130_fd_sc_hd__nor2_2 _14895_ (.A(_04224_),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__and2_1 _14896_ (.A(_04225_),
    .B(_04224_),
    .X(_04227_));
 sky130_fd_sc_hd__nor2_4 _14897_ (.A(_04226_),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__xnor2_4 _14898_ (.A(_03759_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nor2_2 _14899_ (.A(_04229_),
    .B(_04214_),
    .Y(_04230_));
 sky130_fd_sc_hd__inv_2 _14900_ (.A(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__and3b_1 _14901_ (.A_N(_03937_),
    .B(_03944_),
    .C(_04229_),
    .X(_04232_));
 sky130_fd_sc_hd__o21a_1 _14902_ (.A1(_03937_),
    .A2(_03943_),
    .B1(_04229_),
    .X(_04233_));
 sky130_fd_sc_hd__a311oi_4 _14903_ (.A1(_03847_),
    .A2(_03935_),
    .A3(_03936_),
    .B1(_04229_),
    .C1(_03943_),
    .Y(_04235_));
 sky130_fd_sc_hd__nor2_1 _14904_ (.A(_04230_),
    .B(_04232_),
    .Y(_04236_));
 sky130_fd_sc_hd__o211a_1 _14905_ (.A1(_04233_),
    .A2(_04235_),
    .B1(_04211_),
    .C1(_04213_),
    .X(_04237_));
 sky130_fd_sc_hd__o211ai_4 _14906_ (.A1(_04233_),
    .A2(_04235_),
    .B1(_04211_),
    .C1(_04213_),
    .Y(_04238_));
 sky130_fd_sc_hd__a21oi_1 _14907_ (.A1(_04211_),
    .A2(_04213_),
    .B1(_04236_),
    .Y(_04239_));
 sky130_fd_sc_hd__o2bb2ai_2 _14908_ (.A1_N(_04211_),
    .A2_N(_04213_),
    .B1(_04230_),
    .B2(_04232_),
    .Y(_04240_));
 sky130_fd_sc_hd__and3_1 _14909_ (.A(_04071_),
    .B(_04238_),
    .C(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__nand4_4 _14910_ (.A(_04045_),
    .B(_04070_),
    .C(_04238_),
    .D(_04240_),
    .Y(_04242_));
 sky130_fd_sc_hd__o2bb2ai_4 _14911_ (.A1_N(_04045_),
    .A2_N(_04070_),
    .B1(_04237_),
    .B2(_04239_),
    .Y(_04243_));
 sky130_fd_sc_hd__o2bb2ai_4 _14912_ (.A1_N(_04242_),
    .A2_N(_04243_),
    .B1(_03781_),
    .B2(_03792_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_1 _14913_ (.A(_04243_),
    .B(_03802_),
    .Y(_04246_));
 sky130_fd_sc_hd__nand3_2 _14914_ (.A(_04243_),
    .B(_03802_),
    .C(_04242_),
    .Y(_04247_));
 sky130_fd_sc_hd__o21a_1 _14915_ (.A1(_01359_),
    .A2(_03441_),
    .B1(_04052_),
    .X(_04248_));
 sky130_fd_sc_hd__a32oi_4 _14916_ (.A1(_03693_),
    .A2(_04050_),
    .A3(_04051_),
    .B1(_04052_),
    .B2(_03452_),
    .Y(_04249_));
 sky130_fd_sc_hd__o2bb2a_1 _14917_ (.A1_N(_04244_),
    .A2_N(_04247_),
    .B1(_04248_),
    .B2(_04054_),
    .X(_04250_));
 sky130_fd_sc_hd__o2bb2ai_2 _14918_ (.A1_N(_04244_),
    .A2_N(_04247_),
    .B1(_04248_),
    .B2(_04054_),
    .Y(_04251_));
 sky130_fd_sc_hd__o211ai_4 _14919_ (.A1(_04241_),
    .A2(_04246_),
    .B1(_04249_),
    .C1(_04244_),
    .Y(_04252_));
 sky130_fd_sc_hd__a22oi_4 _14920_ (.A1(_04056_),
    .A2(_04060_),
    .B1(_04251_),
    .B2(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__and3_1 _14921_ (.A(_04056_),
    .B(_04251_),
    .C(_04060_),
    .X(_04254_));
 sky130_fd_sc_hd__a2bb2o_2 _14922_ (.A1_N(_04253_),
    .A2_N(_04254_),
    .B1(_03584_),
    .B2(_04058_),
    .X(_04255_));
 sky130_fd_sc_hd__or3b_2 _14923_ (.A(_03595_),
    .B(_04253_),
    .C_N(_04058_),
    .X(_04257_));
 sky130_fd_sc_hd__o21a_1 _14924_ (.A1(_04068_),
    .A2(_04253_),
    .B1(_04255_),
    .X(_04258_));
 sky130_fd_sc_hd__or4b_4 _14925_ (.A(_01797_),
    .B(_04062_),
    .C(_03606_),
    .D_N(_04061_),
    .X(_04259_));
 sky130_fd_sc_hd__a32o_2 _14926_ (.A1(_01786_),
    .A2(_03573_),
    .A3(_04063_),
    .B1(_03671_),
    .B2(_04065_),
    .X(_04260_));
 sky130_fd_sc_hd__a21oi_1 _14927_ (.A1(_04255_),
    .A2(_04257_),
    .B1(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__a21oi_1 _14928_ (.A1(_04255_),
    .A2(_04260_),
    .B1(_04261_),
    .Y(net72));
 sky130_fd_sc_hd__a21oi_1 _14929_ (.A1(_03802_),
    .A2(_04243_),
    .B1(_04241_),
    .Y(_04262_));
 sky130_fd_sc_hd__a32o_1 _14930_ (.A1(_04071_),
    .A2(_04238_),
    .A3(_04240_),
    .B1(_04243_),
    .B2(_03802_),
    .X(_04263_));
 sky130_fd_sc_hd__o21ai_1 _14931_ (.A1(_04118_),
    .A2(_04114_),
    .B1(_04116_),
    .Y(_04264_));
 sky130_fd_sc_hd__a21o_1 _14932_ (.A1(_04096_),
    .A2(_04103_),
    .B1(_04100_),
    .X(_04265_));
 sky130_fd_sc_hd__and2b_4 _14933_ (.A_N(net40),
    .B(net41),
    .X(_04267_));
 sky130_fd_sc_hd__nand2b_4 _14934_ (.A_N(net40),
    .B(net41),
    .Y(_04268_));
 sky130_fd_sc_hd__and2b_4 _14935_ (.A_N(net41),
    .B(net40),
    .X(_04269_));
 sky130_fd_sc_hd__nand2b_4 _14936_ (.A_N(net41),
    .B(net40),
    .Y(_04270_));
 sky130_fd_sc_hd__nand2_1 _14937_ (.A(_04268_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__a22oi_2 _14938_ (.A1(net12),
    .A2(_04217_),
    .B1(_04539_),
    .B2(_04215_),
    .Y(_04272_));
 sky130_fd_sc_hd__a22o_1 _14939_ (.A1(net12),
    .A2(_04217_),
    .B1(_04539_),
    .B2(_04215_),
    .X(_04273_));
 sky130_fd_sc_hd__a32o_1 _14940_ (.A1(net318),
    .A2(_04452_),
    .A3(net285),
    .B1(_03726_),
    .B2(net23),
    .X(_04274_));
 sky130_fd_sc_hd__nand2_1 _14941_ (.A(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__o221ai_4 _14942_ (.A1(_04474_),
    .A2(_03714_),
    .B1(_03737_),
    .B2(_03396_),
    .C1(_04272_),
    .Y(_04276_));
 sky130_fd_sc_hd__o2111ai_4 _14943_ (.A1(net280),
    .A2(_04269_),
    .B1(_04276_),
    .C1(net1),
    .D1(_04275_),
    .Y(_04278_));
 sky130_fd_sc_hd__a22o_1 _14944_ (.A1(net1),
    .A2(_04271_),
    .B1(_04275_),
    .B2(_04276_),
    .X(_04279_));
 sky130_fd_sc_hd__a21oi_1 _14945_ (.A1(_04278_),
    .A2(_04279_),
    .B1(_04265_),
    .Y(_04280_));
 sky130_fd_sc_hd__a221o_1 _14946_ (.A1(_04096_),
    .A2(_04103_),
    .B1(_04278_),
    .B2(_04279_),
    .C1(_04100_),
    .X(_04281_));
 sky130_fd_sc_hd__nand3_1 _14947_ (.A(_04265_),
    .B(_04278_),
    .C(_04279_),
    .Y(_04282_));
 sky130_fd_sc_hd__and2_1 _14948_ (.A(_04281_),
    .B(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__o21a_1 _14949_ (.A1(_04224_),
    .A2(_04225_),
    .B1(_04221_),
    .X(_04284_));
 sky130_fd_sc_hd__a21oi_2 _14950_ (.A1(_04281_),
    .A2(_04282_),
    .B1(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__o2111a_1 _14951_ (.A1(_04225_),
    .A2(_04224_),
    .B1(_04221_),
    .C1(_04282_),
    .D1(_04281_),
    .X(_04286_));
 sky130_fd_sc_hd__nor2_1 _14952_ (.A(_04285_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__o21a_1 _14953_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04264_),
    .X(_04288_));
 sky130_fd_sc_hd__o21ai_2 _14954_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04264_),
    .Y(_04289_));
 sky130_fd_sc_hd__a311o_1 _14955_ (.A1(_04109_),
    .A2(_04110_),
    .A3(_04112_),
    .B1(_04285_),
    .C1(_04286_),
    .X(_04290_));
 sky130_fd_sc_hd__o211ai_4 _14956_ (.A1(_04118_),
    .A2(_04114_),
    .B1(_04116_),
    .C1(_04287_),
    .Y(_04291_));
 sky130_fd_sc_hd__a22oi_4 _14957_ (.A1(_03759_),
    .A2(_04228_),
    .B1(_04289_),
    .B2(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__o2111a_1 _14958_ (.A1(_04290_),
    .A2(_04120_),
    .B1(_03759_),
    .C1(_04228_),
    .D1(_04289_),
    .X(_04293_));
 sky130_fd_sc_hd__or2_1 _14959_ (.A(_04292_),
    .B(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__o21a_1 _14960_ (.A1(_04119_),
    .A2(_04120_),
    .B1(_04206_),
    .X(_04295_));
 sky130_fd_sc_hd__a21o_1 _14961_ (.A1(_04121_),
    .A2(_04204_),
    .B1(_04205_),
    .X(_04296_));
 sky130_fd_sc_hd__o2bb2ai_1 _14962_ (.A1_N(_04169_),
    .A2_N(_04189_),
    .B1(_04183_),
    .B2(_04187_),
    .Y(_04297_));
 sky130_fd_sc_hd__a22oi_2 _14963_ (.A1(_05874_),
    .A2(_11771_),
    .B1(_11793_),
    .B2(net29),
    .Y(_04299_));
 sky130_fd_sc_hd__or3b_1 _14964_ (.A(_03916_),
    .B(net34),
    .C_N(net64),
    .X(_04300_));
 sky130_fd_sc_hd__o211ai_4 _14965_ (.A1(net267),
    .A2(_06508_),
    .B1(net289),
    .C1(_06486_),
    .Y(_04301_));
 sky130_fd_sc_hd__or3b_2 _14966_ (.A(_03938_),
    .B(net64),
    .C_N(net63),
    .X(_04302_));
 sky130_fd_sc_hd__nand3_2 _14967_ (.A(_07242_),
    .B(_07253_),
    .C(_08250_),
    .Y(_04303_));
 sky130_fd_sc_hd__o2111a_1 _14968_ (.A1(_03916_),
    .A2(_10346_),
    .B1(_04301_),
    .C1(_04302_),
    .D1(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__o2111ai_4 _14969_ (.A1(_03916_),
    .A2(_10346_),
    .B1(_04301_),
    .C1(_04302_),
    .D1(_04303_),
    .Y(_04305_));
 sky130_fd_sc_hd__a22oi_1 _14970_ (.A1(_04300_),
    .A2(_04301_),
    .B1(_04302_),
    .B2(_04303_),
    .Y(_04306_));
 sky130_fd_sc_hd__a22o_2 _14971_ (.A1(_04300_),
    .A2(_04301_),
    .B1(_04302_),
    .B2(_04303_),
    .X(_04307_));
 sky130_fd_sc_hd__o21ai_1 _14972_ (.A1(_04304_),
    .A2(_04306_),
    .B1(_04299_),
    .Y(_04308_));
 sky130_fd_sc_hd__nand3b_4 _14973_ (.A_N(_04299_),
    .B(_04305_),
    .C(_04307_),
    .Y(_04310_));
 sky130_fd_sc_hd__a21o_1 _14974_ (.A1(_04075_),
    .A2(_04084_),
    .B1(_04081_),
    .X(_04311_));
 sky130_fd_sc_hd__a21oi_2 _14975_ (.A1(_04308_),
    .A2(_04310_),
    .B1(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__and3_1 _14976_ (.A(_04308_),
    .B(_04310_),
    .C(_04311_),
    .X(_04313_));
 sky130_fd_sc_hd__nand3_1 _14977_ (.A(_04308_),
    .B(_04310_),
    .C(_04311_),
    .Y(_04314_));
 sky130_fd_sc_hd__a32o_1 _14978_ (.A1(net315),
    .A2(net267),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net26),
    .X(_04315_));
 sky130_fd_sc_hd__or3b_1 _14979_ (.A(_03616_),
    .B(net37),
    .C_N(net36),
    .X(_04316_));
 sky130_fd_sc_hd__nand3_1 _14980_ (.A(_04998_),
    .B(net304),
    .C(_01293_),
    .Y(_04317_));
 sky130_fd_sc_hd__or3_1 _14981_ (.A(net36),
    .B(_03993_),
    .C(_03725_),
    .X(_04318_));
 sky130_fd_sc_hd__o211ai_2 _14982_ (.A1(net267),
    .A2(_05436_),
    .B1(_12330_),
    .C1(_05414_),
    .Y(_04319_));
 sky130_fd_sc_hd__a22oi_1 _14983_ (.A1(_04316_),
    .A2(_04317_),
    .B1(_04318_),
    .B2(_04319_),
    .Y(_04321_));
 sky130_fd_sc_hd__a22o_1 _14984_ (.A1(_04316_),
    .A2(_04317_),
    .B1(_04318_),
    .B2(_04319_),
    .X(_04322_));
 sky130_fd_sc_hd__o2111ai_1 _14985_ (.A1(_03616_),
    .A2(_01326_),
    .B1(_04317_),
    .C1(_04318_),
    .D1(_04319_),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2_1 _14986_ (.A(_04322_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__xnor2_1 _14987_ (.A(_04315_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__xor2_1 _14988_ (.A(_04315_),
    .B(_04324_),
    .X(_04326_));
 sky130_fd_sc_hd__o21ai_1 _14989_ (.A1(_04312_),
    .A2(_04313_),
    .B1(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand3b_1 _14990_ (.A_N(_04312_),
    .B(_04314_),
    .C(_04325_),
    .Y(_04328_));
 sky130_fd_sc_hd__o21ai_1 _14991_ (.A1(_04312_),
    .A2(_04313_),
    .B1(_04325_),
    .Y(_04329_));
 sky130_fd_sc_hd__nand3b_1 _14992_ (.A_N(_04312_),
    .B(_04314_),
    .C(_04326_),
    .Y(_04330_));
 sky130_fd_sc_hd__nand3_2 _14993_ (.A(_04297_),
    .B(_04327_),
    .C(_04328_),
    .Y(_04332_));
 sky130_fd_sc_hd__a21oi_1 _14994_ (.A1(_04327_),
    .A2(_04328_),
    .B1(_04297_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand4_2 _14995_ (.A(_04188_),
    .B(_04191_),
    .C(_04329_),
    .D(_04330_),
    .Y(_04334_));
 sky130_fd_sc_hd__a21oi_1 _14996_ (.A1(_04104_),
    .A2(_04105_),
    .B1(_04092_),
    .Y(_04335_));
 sky130_fd_sc_hd__a31o_1 _14997_ (.A1(_04095_),
    .A2(_04104_),
    .A3(_04105_),
    .B1(_04092_),
    .X(_04336_));
 sky130_fd_sc_hd__inv_2 _14998_ (.A(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__o2bb2a_1 _14999_ (.A1_N(_04332_),
    .A2_N(_04334_),
    .B1(_04335_),
    .B2(_04094_),
    .X(_04338_));
 sky130_fd_sc_hd__o2bb2ai_2 _15000_ (.A1_N(_04332_),
    .A2_N(_04334_),
    .B1(_04335_),
    .B2(_04094_),
    .Y(_04339_));
 sky130_fd_sc_hd__and3_1 _15001_ (.A(_04332_),
    .B(_04334_),
    .C(_04336_),
    .X(_04340_));
 sky130_fd_sc_hd__nand3_2 _15002_ (.A(_04332_),
    .B(_04334_),
    .C(_04336_),
    .Y(_04341_));
 sky130_fd_sc_hd__nand2_1 _15003_ (.A(_04339_),
    .B(_04341_),
    .Y(_04343_));
 sky130_fd_sc_hd__a32o_1 _15004_ (.A1(_04125_),
    .A2(_04162_),
    .A3(_04163_),
    .B1(_04191_),
    .B2(_04192_),
    .X(_04344_));
 sky130_fd_sc_hd__o21ai_2 _15005_ (.A1(_04164_),
    .A2(_04196_),
    .B1(_04167_),
    .Y(_04345_));
 sky130_fd_sc_hd__a31o_2 _15006_ (.A1(_04167_),
    .A2(_04193_),
    .A3(_04194_),
    .B1(_04164_),
    .X(_04346_));
 sky130_fd_sc_hd__a21bo_1 _15007_ (.A1(_04174_),
    .A2(_04181_),
    .B1_N(_04182_),
    .X(_04347_));
 sky130_fd_sc_hd__a32oi_4 _15008_ (.A1(_04151_),
    .A2(_04152_),
    .A3(_04154_),
    .B1(_04156_),
    .B2(_04149_),
    .Y(_04348_));
 sky130_fd_sc_hd__a32o_1 _15009_ (.A1(_04151_),
    .A2(_04152_),
    .A3(_04154_),
    .B1(_04156_),
    .B2(_04149_),
    .X(_04349_));
 sky130_fd_sc_hd__a32o_1 _15010_ (.A1(_08700_),
    .A2(_07658_),
    .A3(net256),
    .B1(_07680_),
    .B2(net32),
    .X(_04350_));
 sky130_fd_sc_hd__and3_1 _15011_ (.A(_03927_),
    .B(net2),
    .C(net61),
    .X(_04351_));
 sky130_fd_sc_hd__a31oi_2 _15012_ (.A1(_09698_),
    .A2(net292),
    .A3(net255),
    .B1(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__a31o_1 _15013_ (.A1(_09698_),
    .A2(net292),
    .A3(net255),
    .B1(_04351_),
    .X(_04354_));
 sky130_fd_sc_hd__nor2_1 _15014_ (.A(_03982_),
    .B(net298),
    .Y(_04355_));
 sky130_fd_sc_hd__or3b_1 _15015_ (.A(net61),
    .B(_03982_),
    .C_N(net60),
    .X(_04356_));
 sky130_fd_sc_hd__a221oi_2 _15016_ (.A1(_09676_),
    .A2(net3),
    .B1(_06519_),
    .B2(_11376_),
    .C1(_05699_),
    .Y(_04357_));
 sky130_fd_sc_hd__o211ai_4 _15017_ (.A1(_05699_),
    .A2(net236),
    .B1(_04356_),
    .C1(_04352_),
    .Y(_04358_));
 sky130_fd_sc_hd__o21ai_2 _15018_ (.A1(_04355_),
    .A2(_04357_),
    .B1(_04354_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand3b_1 _15019_ (.A_N(_04350_),
    .B(_04358_),
    .C(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__a21bo_1 _15020_ (.A1(_04358_),
    .A2(_04359_),
    .B1_N(_04350_),
    .X(_04361_));
 sky130_fd_sc_hd__a21boi_2 _15021_ (.A1(_04350_),
    .A2(_04358_),
    .B1_N(_04359_),
    .Y(_04362_));
 sky130_fd_sc_hd__and3_1 _15022_ (.A(_04350_),
    .B(_04358_),
    .C(_04359_),
    .X(_04363_));
 sky130_fd_sc_hd__nand3_1 _15023_ (.A(_04350_),
    .B(_04358_),
    .C(_04359_),
    .Y(_04365_));
 sky130_fd_sc_hd__a21o_1 _15024_ (.A1(_04358_),
    .A2(_04359_),
    .B1(_04350_),
    .X(_04366_));
 sky130_fd_sc_hd__nand2_1 _15025_ (.A(_04366_),
    .B(_04348_),
    .Y(_04367_));
 sky130_fd_sc_hd__and3_2 _15026_ (.A(_04366_),
    .B(_04348_),
    .C(_04365_),
    .X(_04368_));
 sky130_fd_sc_hd__nand3_1 _15027_ (.A(_04366_),
    .B(_04348_),
    .C(_04365_),
    .Y(_04369_));
 sky130_fd_sc_hd__nand3_2 _15028_ (.A(_04349_),
    .B(_04360_),
    .C(_04361_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_2 _15029_ (.A(_04370_),
    .B(_04347_),
    .Y(_04371_));
 sky130_fd_sc_hd__a31o_1 _15030_ (.A1(_04348_),
    .A2(_04365_),
    .A3(_04366_),
    .B1(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__a21o_2 _15031_ (.A1(_04369_),
    .A2(_04370_),
    .B1(_04347_),
    .X(_04373_));
 sky130_fd_sc_hd__o21ai_4 _15032_ (.A1(_04368_),
    .A2(_04371_),
    .B1(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__o21a_1 _15033_ (.A1(_04158_),
    .A2(_04160_),
    .B1(_04148_),
    .X(_04376_));
 sky130_fd_sc_hd__a31o_1 _15034_ (.A1(_04144_),
    .A2(_04159_),
    .A3(_04161_),
    .B1(_04147_),
    .X(_04377_));
 sky130_fd_sc_hd__a32o_1 _15035_ (.A1(net235),
    .A2(_12999_),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net4),
    .X(_04378_));
 sky130_fd_sc_hd__nand3_2 _15036_ (.A(_02421_),
    .B(net249),
    .C(net317),
    .Y(_04379_));
 sky130_fd_sc_hd__or3b_1 _15037_ (.A(net58),
    .B(_04026_),
    .C_N(net55),
    .X(_04380_));
 sky130_fd_sc_hd__and3b_1 _15038_ (.A_N(net59),
    .B(net5),
    .C(net58),
    .X(_04381_));
 sky130_fd_sc_hd__or3b_2 _15039_ (.A(net59),
    .B(_04015_),
    .C_N(net58),
    .X(_04382_));
 sky130_fd_sc_hd__o311a_1 _15040_ (.A1(net263),
    .A2(_11387_),
    .A3(_00646_),
    .B1(net305),
    .C1(_00625_),
    .X(_04383_));
 sky130_fd_sc_hd__o211ai_4 _15041_ (.A1(_11431_),
    .A2(_00646_),
    .B1(net305),
    .C1(_00625_),
    .Y(_04384_));
 sky130_fd_sc_hd__a22oi_2 _15042_ (.A1(_04379_),
    .A2(_04380_),
    .B1(_04382_),
    .B2(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__o2bb2ai_1 _15043_ (.A1_N(_04379_),
    .A2_N(_04380_),
    .B1(_04381_),
    .B2(_04383_),
    .Y(_04387_));
 sky130_fd_sc_hd__o2111ai_4 _15044_ (.A1(_04026_),
    .A2(net316),
    .B1(_04379_),
    .C1(_04382_),
    .D1(_04384_),
    .Y(_04388_));
 sky130_fd_sc_hd__a21boi_1 _15045_ (.A1(_04387_),
    .A2(_04388_),
    .B1_N(_04378_),
    .Y(_04389_));
 sky130_fd_sc_hd__a21bo_1 _15046_ (.A1(_04387_),
    .A2(_04388_),
    .B1_N(_04378_),
    .X(_04390_));
 sky130_fd_sc_hd__nor3b_1 _15047_ (.A(_04378_),
    .B(_04385_),
    .C_N(_04388_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand3b_1 _15048_ (.A_N(_04378_),
    .B(_04387_),
    .C(_04388_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2_1 _15049_ (.A(_04390_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__o221a_1 _15050_ (.A1(_04026_),
    .A2(_04375_),
    .B1(_02475_),
    .B2(_04353_),
    .C1(_04137_),
    .X(_04394_));
 sky130_fd_sc_hd__nand2_1 _15051_ (.A(_04128_),
    .B(_04139_),
    .Y(_04395_));
 sky130_fd_sc_hd__a21o_1 _15052_ (.A1(_04128_),
    .A2(_04139_),
    .B1(_04136_),
    .X(_04396_));
 sky130_fd_sc_hd__nor2_1 _15053_ (.A(_04048_),
    .B(_04375_),
    .Y(_04398_));
 sky130_fd_sc_hd__o311a_1 _15054_ (.A1(net263),
    .A2(_11387_),
    .A3(_03954_),
    .B1(_04342_),
    .C1(_03952_),
    .X(_04399_));
 sky130_fd_sc_hd__o32a_1 _15055_ (.A1(_04353_),
    .A2(net247),
    .A3(_03957_),
    .B1(_04375_),
    .B2(_04048_),
    .X(_04400_));
 sky130_fd_sc_hd__a31o_1 _15056_ (.A1(_03952_),
    .A2(net232),
    .A3(_04342_),
    .B1(_04398_),
    .X(_04401_));
 sky130_fd_sc_hd__nor2_1 _15057_ (.A(_04059_),
    .B(_04331_),
    .Y(_04402_));
 sky130_fd_sc_hd__or3_1 _15058_ (.A(net44),
    .B(net9),
    .C(_03286_),
    .X(_04403_));
 sky130_fd_sc_hd__and3_1 _15059_ (.A(net8),
    .B(_04320_),
    .C(_04069_),
    .X(_04404_));
 sky130_fd_sc_hd__or4_1 _15060_ (.A(net44),
    .B(net9),
    .C(_04059_),
    .D(_03286_),
    .X(_04405_));
 sky130_fd_sc_hd__nor2_4 _15061_ (.A(net8),
    .B(net9),
    .Y(_04406_));
 sky130_fd_sc_hd__or2_4 _15062_ (.A(net8),
    .B(net9),
    .X(_04407_));
 sky130_fd_sc_hd__nand4_4 _15063_ (.A(_06519_),
    .B(net287),
    .C(_03953_),
    .D(_04406_),
    .Y(_04409_));
 sky130_fd_sc_hd__a41oi_4 _15064_ (.A1(_11398_),
    .A2(_04059_),
    .A3(net308),
    .A4(net284),
    .B1(_04069_),
    .Y(_04410_));
 sky130_fd_sc_hd__o41ai_4 _15065_ (.A1(net8),
    .A2(net267),
    .A3(_06508_),
    .A4(net245),
    .B1(net9),
    .Y(_04411_));
 sky130_fd_sc_hd__o31ai_4 _15066_ (.A1(net7),
    .A2(net249),
    .A3(_04407_),
    .B1(net226),
    .Y(_04412_));
 sky130_fd_sc_hd__nand3_1 _15067_ (.A(net226),
    .B(net33),
    .C(net188),
    .Y(_04413_));
 sky130_fd_sc_hd__a31oi_2 _15068_ (.A1(_04132_),
    .A2(_04484_),
    .A3(_04130_),
    .B1(_04402_),
    .Y(_04414_));
 sky130_fd_sc_hd__nand2_1 _15069_ (.A(_04414_),
    .B(_04413_),
    .Y(_04415_));
 sky130_fd_sc_hd__o2bb2ai_1 _15070_ (.A1_N(_04413_),
    .A2_N(_04414_),
    .B1(_04059_),
    .B2(_04403_),
    .Y(_04416_));
 sky130_fd_sc_hd__o21ai_1 _15071_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__a211o_1 _15072_ (.A1(_04414_),
    .A2(_04413_),
    .B1(_04404_),
    .C1(_04401_),
    .X(_04418_));
 sky130_fd_sc_hd__o2bb2ai_1 _15073_ (.A1_N(_04413_),
    .A2_N(_04414_),
    .B1(_04398_),
    .B2(_04399_),
    .Y(_04420_));
 sky130_fd_sc_hd__a21oi_1 _15074_ (.A1(_04405_),
    .A2(_04415_),
    .B1(_04401_),
    .Y(_04421_));
 sky130_fd_sc_hd__nand2_1 _15075_ (.A(_04416_),
    .B(_04400_),
    .Y(_04422_));
 sky130_fd_sc_hd__o211ai_4 _15076_ (.A1(_04138_),
    .A2(_04394_),
    .B1(_04417_),
    .C1(_04418_),
    .Y(_04423_));
 sky130_fd_sc_hd__o2bb2ai_1 _15077_ (.A1_N(_04137_),
    .A2_N(_04395_),
    .B1(_04404_),
    .B2(_04420_),
    .Y(_04424_));
 sky130_fd_sc_hd__o211ai_2 _15078_ (.A1(_04404_),
    .A2(_04420_),
    .B1(_04396_),
    .C1(_04422_),
    .Y(_04425_));
 sky130_fd_sc_hd__o221a_2 _15079_ (.A1(_04389_),
    .A2(_04391_),
    .B1(_04421_),
    .B2(_04424_),
    .C1(_04423_),
    .X(_04426_));
 sky130_fd_sc_hd__a21oi_2 _15080_ (.A1(_04423_),
    .A2(_04425_),
    .B1(_04393_),
    .Y(_04427_));
 sky130_fd_sc_hd__a21o_1 _15081_ (.A1(_04423_),
    .A2(_04425_),
    .B1(_04393_),
    .X(_04428_));
 sky130_fd_sc_hd__nand3b_4 _15082_ (.A_N(_04426_),
    .B(_04428_),
    .C(_04377_),
    .Y(_04429_));
 sky130_fd_sc_hd__o22a_1 _15083_ (.A1(_04145_),
    .A2(_04376_),
    .B1(_04426_),
    .B2(_04427_),
    .X(_04431_));
 sky130_fd_sc_hd__o22ai_4 _15084_ (.A1(_04145_),
    .A2(_04376_),
    .B1(_04426_),
    .B2(_04427_),
    .Y(_04432_));
 sky130_fd_sc_hd__a21o_2 _15085_ (.A1(_04429_),
    .A2(_04432_),
    .B1(_04374_),
    .X(_04433_));
 sky130_fd_sc_hd__nand3_4 _15086_ (.A(_04374_),
    .B(_04429_),
    .C(_04432_),
    .Y(_04434_));
 sky130_fd_sc_hd__o2111ai_4 _15087_ (.A1(_04368_),
    .A2(_04371_),
    .B1(_04373_),
    .C1(_04429_),
    .D1(_04432_),
    .Y(_04435_));
 sky130_fd_sc_hd__a22o_2 _15088_ (.A1(_04372_),
    .A2(_04373_),
    .B1(_04429_),
    .B2(_04432_),
    .X(_04436_));
 sky130_fd_sc_hd__a22oi_4 _15089_ (.A1(_04167_),
    .A2(_04198_),
    .B1(_04433_),
    .B2(_04434_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand3_4 _15090_ (.A(_04436_),
    .B(_04345_),
    .C(_04435_),
    .Y(_04438_));
 sky130_fd_sc_hd__a22oi_4 _15091_ (.A1(_04165_),
    .A2(_04344_),
    .B1(_04435_),
    .B2(_04436_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand3_4 _15092_ (.A(_04346_),
    .B(_04433_),
    .C(_04434_),
    .Y(_04440_));
 sky130_fd_sc_hd__a31oi_4 _15093_ (.A1(_04346_),
    .A2(_04433_),
    .A3(_04434_),
    .B1(_04343_),
    .Y(_04442_));
 sky130_fd_sc_hd__nand4_4 _15094_ (.A(_04339_),
    .B(_04341_),
    .C(_04438_),
    .D(_04440_),
    .Y(_04443_));
 sky130_fd_sc_hd__a2bb2oi_1 _15095_ (.A1_N(_04338_),
    .A2_N(_04340_),
    .B1(_04438_),
    .B2(_04440_),
    .Y(_04444_));
 sky130_fd_sc_hd__o22ai_4 _15096_ (.A1(_04338_),
    .A2(_04340_),
    .B1(_04437_),
    .B2(_04439_),
    .Y(_04445_));
 sky130_fd_sc_hd__o211ai_1 _15097_ (.A1(_04338_),
    .A2(_04340_),
    .B1(_04438_),
    .C1(_04440_),
    .Y(_04446_));
 sky130_fd_sc_hd__a21o_1 _15098_ (.A1(_04438_),
    .A2(_04440_),
    .B1(_04343_),
    .X(_04447_));
 sky130_fd_sc_hd__a221oi_4 _15099_ (.A1(_04206_),
    .A2(_04210_),
    .B1(_04438_),
    .B2(_04442_),
    .C1(_04444_),
    .Y(_04448_));
 sky130_fd_sc_hd__nand3_2 _15100_ (.A(_04445_),
    .B(_04296_),
    .C(_04443_),
    .Y(_04449_));
 sky130_fd_sc_hd__a2bb2oi_4 _15101_ (.A1_N(_04203_),
    .A2_N(_04295_),
    .B1(_04443_),
    .B2(_04445_),
    .Y(_04450_));
 sky130_fd_sc_hd__o211ai_2 _15102_ (.A1(_04203_),
    .A2(_04295_),
    .B1(_04446_),
    .C1(_04447_),
    .Y(_04451_));
 sky130_fd_sc_hd__nand3b_2 _15103_ (.A_N(_04294_),
    .B(_04449_),
    .C(_04451_),
    .Y(_04453_));
 sky130_fd_sc_hd__a21boi_1 _15104_ (.A1(_04449_),
    .A2(_04451_),
    .B1_N(_04294_),
    .Y(_04454_));
 sky130_fd_sc_hd__o22ai_4 _15105_ (.A1(_04292_),
    .A2(_04293_),
    .B1(_04448_),
    .B2(_04450_),
    .Y(_04455_));
 sky130_fd_sc_hd__a21boi_1 _15106_ (.A1(_04211_),
    .A2(_04236_),
    .B1_N(_04213_),
    .Y(_04456_));
 sky130_fd_sc_hd__a21boi_2 _15107_ (.A1(_04453_),
    .A2(_04455_),
    .B1_N(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__a21bo_1 _15108_ (.A1(_04453_),
    .A2(_04455_),
    .B1_N(_04456_),
    .X(_04458_));
 sky130_fd_sc_hd__nor3b_1 _15109_ (.A(_04456_),
    .B(_04454_),
    .C_N(_04453_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand3b_2 _15110_ (.A_N(_04456_),
    .B(_04455_),
    .C(_04453_),
    .Y(_04460_));
 sky130_fd_sc_hd__o21ai_1 _15111_ (.A1(_04457_),
    .A2(_04459_),
    .B1(_04230_),
    .Y(_04461_));
 sky130_fd_sc_hd__o211ai_2 _15112_ (.A1(_04229_),
    .A2(_04214_),
    .B1(_04460_),
    .C1(_04458_),
    .Y(_04462_));
 sky130_fd_sc_hd__o22ai_2 _15113_ (.A1(_04214_),
    .A2(_04229_),
    .B1(_04457_),
    .B2(_04459_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand3_1 _15114_ (.A(_04458_),
    .B(_04460_),
    .C(_04230_),
    .Y(_04465_));
 sky130_fd_sc_hd__and3_1 _15115_ (.A(_04461_),
    .B(_04462_),
    .C(_04262_),
    .X(_04466_));
 sky130_fd_sc_hd__nand3_1 _15116_ (.A(_04461_),
    .B(_04462_),
    .C(_04262_),
    .Y(_04467_));
 sky130_fd_sc_hd__a32oi_1 _15117_ (.A1(_04458_),
    .A2(_04460_),
    .A3(_04230_),
    .B1(_04242_),
    .B2(_04246_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand3_2 _15118_ (.A(_04263_),
    .B(_04464_),
    .C(_04465_),
    .Y(_04469_));
 sky130_fd_sc_hd__a31oi_1 _15119_ (.A1(_04262_),
    .A2(_04461_),
    .A3(_04462_),
    .B1(_04252_),
    .Y(_04470_));
 sky130_fd_sc_hd__a31o_1 _15120_ (.A1(_04262_),
    .A2(_04461_),
    .A3(_04462_),
    .B1(_04252_),
    .X(_04471_));
 sky130_fd_sc_hd__a32oi_4 _15121_ (.A1(_04244_),
    .A2(_04249_),
    .A3(_04247_),
    .B1(_04469_),
    .B2(_04467_),
    .Y(_04472_));
 sky130_fd_sc_hd__nor2_1 _15122_ (.A(_04470_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__o22ai_1 _15123_ (.A1(_04061_),
    .A2(_04250_),
    .B1(_04470_),
    .B2(_04472_),
    .Y(_04475_));
 sky130_fd_sc_hd__o31a_2 _15124_ (.A1(_04061_),
    .A2(_04250_),
    .A3(_04472_),
    .B1(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__a2bb2o_1 _15125_ (.A1_N(_04068_),
    .A2_N(_04253_),
    .B1(_04258_),
    .B2(_04260_),
    .X(_04477_));
 sky130_fd_sc_hd__xor2_1 _15126_ (.A(_04476_),
    .B(_04477_),
    .X(net73));
 sky130_fd_sc_hd__o21a_1 _15127_ (.A1(_04292_),
    .A2(_04293_),
    .B1(_04449_),
    .X(_04478_));
 sky130_fd_sc_hd__o21ai_1 _15128_ (.A1(_04294_),
    .A2(_04450_),
    .B1(_04449_),
    .Y(_04479_));
 sky130_fd_sc_hd__and2b_4 _15129_ (.A_N(net41),
    .B(net42),
    .X(_04480_));
 sky130_fd_sc_hd__nand2b_4 _15130_ (.A_N(net41),
    .B(net42),
    .Y(_04481_));
 sky130_fd_sc_hd__and2b_4 _15131_ (.A_N(net42),
    .B(net41),
    .X(_04482_));
 sky130_fd_sc_hd__nand2b_4 _15132_ (.A_N(net42),
    .B(net41),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _15133_ (.A(_04481_),
    .B(_04483_),
    .Y(_04485_));
 sky130_fd_sc_hd__a21o_1 _15134_ (.A1(_04315_),
    .A2(_04323_),
    .B1(_04321_),
    .X(_04486_));
 sky130_fd_sc_hd__o2bb2a_1 _15135_ (.A1_N(net12),
    .A2_N(_04269_),
    .B1(_04268_),
    .B2(_04528_),
    .X(_04487_));
 sky130_fd_sc_hd__a22o_1 _15136_ (.A1(net12),
    .A2(_04269_),
    .B1(_04539_),
    .B2(net280),
    .X(_04488_));
 sky130_fd_sc_hd__nand2_1 _15137_ (.A(net23),
    .B(_04217_),
    .Y(_04489_));
 sky130_fd_sc_hd__nand3_2 _15138_ (.A(net318),
    .B(_04452_),
    .C(_04215_),
    .Y(_04490_));
 sky130_fd_sc_hd__nand3_2 _15139_ (.A(net315),
    .B(net267),
    .C(net285),
    .Y(_04491_));
 sky130_fd_sc_hd__nand2_1 _15140_ (.A(net26),
    .B(_03726_),
    .Y(_04492_));
 sky130_fd_sc_hd__and4_1 _15141_ (.A(_04489_),
    .B(_04490_),
    .C(_04491_),
    .D(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__o2111ai_1 _15142_ (.A1(_03396_),
    .A2(_04218_),
    .B1(_04490_),
    .C1(_04491_),
    .D1(_04492_),
    .Y(_04494_));
 sky130_fd_sc_hd__a22oi_4 _15143_ (.A1(_04489_),
    .A2(_04490_),
    .B1(_04491_),
    .B2(_04492_),
    .Y(_04496_));
 sky130_fd_sc_hd__a22o_1 _15144_ (.A1(_04489_),
    .A2(_04490_),
    .B1(_04491_),
    .B2(_04492_),
    .X(_04497_));
 sky130_fd_sc_hd__o21ai_1 _15145_ (.A1(_04493_),
    .A2(_04496_),
    .B1(_04487_),
    .Y(_04498_));
 sky130_fd_sc_hd__and3_1 _15146_ (.A(_04488_),
    .B(_04494_),
    .C(_04497_),
    .X(_04499_));
 sky130_fd_sc_hd__nand3_1 _15147_ (.A(_04488_),
    .B(_04494_),
    .C(_04497_),
    .Y(_04500_));
 sky130_fd_sc_hd__a21oi_1 _15148_ (.A1(_04498_),
    .A2(_04500_),
    .B1(_04486_),
    .Y(_04501_));
 sky130_fd_sc_hd__a21o_1 _15149_ (.A1(_04498_),
    .A2(_04500_),
    .B1(_04486_),
    .X(_04502_));
 sky130_fd_sc_hd__nand3_1 _15150_ (.A(_04486_),
    .B(_04498_),
    .C(_04500_),
    .Y(_04503_));
 sky130_fd_sc_hd__o221a_1 _15151_ (.A1(net280),
    .A2(_04269_),
    .B1(_04273_),
    .B2(_04274_),
    .C1(net1),
    .X(_04504_));
 sky130_fd_sc_hd__a21oi_1 _15152_ (.A1(_04273_),
    .A2(_04274_),
    .B1(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__a21bo_1 _15153_ (.A1(_04502_),
    .A2(_04503_),
    .B1_N(_04505_),
    .X(_04507_));
 sky130_fd_sc_hd__nand3b_1 _15154_ (.A_N(_04505_),
    .B(_04503_),
    .C(_04502_),
    .Y(_04508_));
 sky130_fd_sc_hd__o21ai_1 _15155_ (.A1(_04221_),
    .A2(_04280_),
    .B1(_04282_),
    .Y(_04509_));
 sky130_fd_sc_hd__a21o_1 _15156_ (.A1(_04507_),
    .A2(_04508_),
    .B1(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__nand3_2 _15157_ (.A(_04507_),
    .B(_04508_),
    .C(_04509_),
    .Y(_04511_));
 sky130_fd_sc_hd__a22o_1 _15158_ (.A1(net1),
    .A2(_04485_),
    .B1(_04510_),
    .B2(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__o2111ai_4 _15159_ (.A1(_04480_),
    .A2(_04482_),
    .B1(_04511_),
    .C1(net1),
    .D1(_04510_),
    .Y(_04513_));
 sky130_fd_sc_hd__o21ai_2 _15160_ (.A1(_04337_),
    .A2(_04333_),
    .B1(_04332_),
    .Y(_04514_));
 sky130_fd_sc_hd__and3_1 _15161_ (.A(_04512_),
    .B(_04513_),
    .C(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__nand3_2 _15162_ (.A(_04512_),
    .B(_04513_),
    .C(_04514_),
    .Y(_04516_));
 sky130_fd_sc_hd__a21o_1 _15163_ (.A1(_04512_),
    .A2(_04513_),
    .B1(_04514_),
    .X(_04518_));
 sky130_fd_sc_hd__a22oi_4 _15164_ (.A1(_04226_),
    .A2(_04283_),
    .B1(_04516_),
    .B2(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__and3_1 _15165_ (.A(_04516_),
    .B(_04283_),
    .C(_04226_),
    .X(_04520_));
 sky130_fd_sc_hd__and4_2 _15166_ (.A(_04518_),
    .B(_04283_),
    .C(_04226_),
    .D(_04516_),
    .X(_04521_));
 sky130_fd_sc_hd__a21oi_1 _15167_ (.A1(_04520_),
    .A2(_04518_),
    .B1(_04519_),
    .Y(_04522_));
 sky130_fd_sc_hd__a32o_1 _15168_ (.A1(_04436_),
    .A2(_04345_),
    .A3(_04435_),
    .B1(_04341_),
    .B2(_04339_),
    .X(_04523_));
 sky130_fd_sc_hd__a31o_1 _15169_ (.A1(_04345_),
    .A2(_04435_),
    .A3(_04436_),
    .B1(_04442_),
    .X(_04524_));
 sky130_fd_sc_hd__o41a_1 _15170_ (.A1(_04145_),
    .A2(_04376_),
    .A3(_04426_),
    .A4(_04427_),
    .B1(_04374_),
    .X(_04525_));
 sky130_fd_sc_hd__o21ai_2 _15171_ (.A1(_04374_),
    .A2(_04431_),
    .B1(_04429_),
    .Y(_04526_));
 sky130_fd_sc_hd__a32o_1 _15172_ (.A1(_09698_),
    .A2(_07658_),
    .A3(net255),
    .B1(_07680_),
    .B2(net2),
    .X(_04527_));
 sky130_fd_sc_hd__o211ai_4 _15173_ (.A1(net263),
    .A2(_11387_),
    .B1(net292),
    .C1(_11354_),
    .Y(_04529_));
 sky130_fd_sc_hd__or3b_1 _15174_ (.A(net62),
    .B(_03982_),
    .C_N(net61),
    .X(_04530_));
 sky130_fd_sc_hd__o211ai_4 _15175_ (.A1(_11387_),
    .A2(_12988_),
    .B1(net299),
    .C1(net235),
    .Y(_04531_));
 sky130_fd_sc_hd__or3b_2 _15176_ (.A(net61),
    .B(_04004_),
    .C_N(net60),
    .X(_04532_));
 sky130_fd_sc_hd__a22oi_2 _15177_ (.A1(_04529_),
    .A2(_04530_),
    .B1(_04531_),
    .B2(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__a22o_1 _15178_ (.A1(_04529_),
    .A2(_04530_),
    .B1(_04531_),
    .B2(_04532_),
    .X(_04534_));
 sky130_fd_sc_hd__and4_1 _15179_ (.A(_04529_),
    .B(_04530_),
    .C(_04531_),
    .D(_04532_),
    .X(_04535_));
 sky130_fd_sc_hd__o2111ai_4 _15180_ (.A1(_03982_),
    .A2(_06859_),
    .B1(_04529_),
    .C1(_04531_),
    .D1(_04532_),
    .Y(_04536_));
 sky130_fd_sc_hd__o21bai_1 _15181_ (.A1(_04533_),
    .A2(_04535_),
    .B1_N(_04527_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand3_1 _15182_ (.A(_04527_),
    .B(_04534_),
    .C(_04536_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand3b_1 _15183_ (.A_N(_04527_),
    .B(_04534_),
    .C(_04536_),
    .Y(_04540_));
 sky130_fd_sc_hd__o21ai_1 _15184_ (.A1(_04533_),
    .A2(_04535_),
    .B1(_04527_),
    .Y(_04541_));
 sky130_fd_sc_hd__a21o_1 _15185_ (.A1(_04378_),
    .A2(_04388_),
    .B1(_04385_),
    .X(_04542_));
 sky130_fd_sc_hd__a21oi_1 _15186_ (.A1(_04378_),
    .A2(_04388_),
    .B1(_04385_),
    .Y(_04543_));
 sky130_fd_sc_hd__a21oi_2 _15187_ (.A1(_04537_),
    .A2(_04538_),
    .B1(_04542_),
    .Y(_04544_));
 sky130_fd_sc_hd__a21o_1 _15188_ (.A1(_04537_),
    .A2(_04538_),
    .B1(_04542_),
    .X(_04545_));
 sky130_fd_sc_hd__a21oi_1 _15189_ (.A1(_04540_),
    .A2(_04541_),
    .B1(_04543_),
    .Y(_04546_));
 sky130_fd_sc_hd__a21o_1 _15190_ (.A1(_04540_),
    .A2(_04541_),
    .B1(_04543_),
    .X(_04547_));
 sky130_fd_sc_hd__nand3b_2 _15191_ (.A_N(_04362_),
    .B(_04545_),
    .C(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__o21ai_2 _15192_ (.A1(_04544_),
    .A2(_04546_),
    .B1(_04362_),
    .Y(_04549_));
 sky130_fd_sc_hd__nand2_2 _15193_ (.A(_04548_),
    .B(_04549_),
    .Y(_04551_));
 sky130_fd_sc_hd__a22o_2 _15194_ (.A1(_04069_),
    .A2(_04402_),
    .B1(_04415_),
    .B2(_04401_),
    .X(_04552_));
 sky130_fd_sc_hd__a32o_2 _15195_ (.A1(_04132_),
    .A2(_04342_),
    .A3(_04130_),
    .B1(_04364_),
    .B2(net8),
    .X(_04553_));
 sky130_fd_sc_hd__a41oi_4 _15196_ (.A1(_06519_),
    .A2(net287),
    .A3(net283),
    .A4(_04406_),
    .B1(_04080_),
    .Y(_04554_));
 sky130_fd_sc_hd__o31ai_4 _15197_ (.A1(net262),
    .A2(net245),
    .A3(_04407_),
    .B1(net10),
    .Y(_04555_));
 sky130_fd_sc_hd__and3_4 _15198_ (.A(_04059_),
    .B(_04069_),
    .C(_04080_),
    .X(_04556_));
 sky130_fd_sc_hd__or3_4 _15199_ (.A(net8),
    .B(net9),
    .C(net10),
    .X(_04557_));
 sky130_fd_sc_hd__nor3_4 _15200_ (.A(net260),
    .B(_03956_),
    .C(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__nand3_4 _15201_ (.A(_06519_),
    .B(_03955_),
    .C(_04556_),
    .Y(_04559_));
 sky130_fd_sc_hd__o31a_2 _15202_ (.A1(net7),
    .A2(net249),
    .A3(_04557_),
    .B1(_04555_),
    .X(_04560_));
 sky130_fd_sc_hd__o21ai_4 _15203_ (.A1(_03958_),
    .A2(_04557_),
    .B1(_04555_),
    .Y(_04562_));
 sky130_fd_sc_hd__nand3_1 _15204_ (.A(_04555_),
    .B(_04559_),
    .C(net33),
    .Y(_04563_));
 sky130_fd_sc_hd__nand3_1 _15205_ (.A(net226),
    .B(_04484_),
    .C(net188),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_1 _15206_ (.A(_04069_),
    .B(_04331_),
    .Y(_04565_));
 sky130_fd_sc_hd__or3_2 _15207_ (.A(net44),
    .B(_04069_),
    .C(_03286_),
    .X(_04566_));
 sky130_fd_sc_hd__or4_1 _15208_ (.A(net44),
    .B(net10),
    .C(_04069_),
    .D(_03286_),
    .X(_04567_));
 sky130_fd_sc_hd__nand3_4 _15209_ (.A(_04563_),
    .B(_04564_),
    .C(_04566_),
    .Y(_04568_));
 sky130_fd_sc_hd__a21oi_1 _15210_ (.A1(_04567_),
    .A2(_04568_),
    .B1(_04553_),
    .Y(_04569_));
 sky130_fd_sc_hd__a21o_1 _15211_ (.A1(_04567_),
    .A2(_04568_),
    .B1(_04553_),
    .X(_04570_));
 sky130_fd_sc_hd__o311a_1 _15212_ (.A1(_03286_),
    .A2(_04562_),
    .A3(_04566_),
    .B1(_04568_),
    .C1(_04553_),
    .X(_04571_));
 sky130_fd_sc_hd__nand3_2 _15213_ (.A(_04553_),
    .B(_04567_),
    .C(_04568_),
    .Y(_04573_));
 sky130_fd_sc_hd__a21oi_2 _15214_ (.A1(_04570_),
    .A2(_04573_),
    .B1(_04552_),
    .Y(_04574_));
 sky130_fd_sc_hd__o21bai_4 _15215_ (.A1(_04569_),
    .A2(_04571_),
    .B1_N(_04552_),
    .Y(_04575_));
 sky130_fd_sc_hd__and3_1 _15216_ (.A(_04552_),
    .B(_04570_),
    .C(_04573_),
    .X(_04576_));
 sky130_fd_sc_hd__nand3_4 _15217_ (.A(_04552_),
    .B(_04570_),
    .C(_04573_),
    .Y(_04577_));
 sky130_fd_sc_hd__o22a_1 _15218_ (.A1(_04015_),
    .A2(_05260_),
    .B1(_00668_),
    .B2(_05238_),
    .X(_04578_));
 sky130_fd_sc_hd__a32o_1 _15219_ (.A1(_00625_),
    .A2(_00657_),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net5),
    .X(_04579_));
 sky130_fd_sc_hd__and3b_1 _15220_ (.A_N(net59),
    .B(net6),
    .C(net58),
    .X(_04580_));
 sky130_fd_sc_hd__or3b_2 _15221_ (.A(net59),
    .B(_04026_),
    .C_N(net58),
    .X(_04581_));
 sky130_fd_sc_hd__a31o_1 _15222_ (.A1(_02421_),
    .A2(net249),
    .A3(net305),
    .B1(_04580_),
    .X(_04582_));
 sky130_fd_sc_hd__o21a_1 _15223_ (.A1(net263),
    .A2(net245),
    .B1(net317),
    .X(_04584_));
 sky130_fd_sc_hd__a22oi_2 _15224_ (.A1(net7),
    .A2(_04649_),
    .B1(_04584_),
    .B2(_03952_),
    .Y(_04585_));
 sky130_fd_sc_hd__o2bb2ai_1 _15225_ (.A1_N(_03952_),
    .A2_N(_04584_),
    .B1(_04048_),
    .B2(net316),
    .Y(_04586_));
 sky130_fd_sc_hd__nand2_2 _15226_ (.A(_04582_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__o211a_1 _15227_ (.A1(_04900_),
    .A2(_02475_),
    .B1(_04581_),
    .C1(_04585_),
    .X(_04588_));
 sky130_fd_sc_hd__o211ai_4 _15228_ (.A1(_04900_),
    .A2(_02475_),
    .B1(_04581_),
    .C1(_04585_),
    .Y(_04589_));
 sky130_fd_sc_hd__a21oi_2 _15229_ (.A1(_04587_),
    .A2(_04589_),
    .B1(_04579_),
    .Y(_04590_));
 sky130_fd_sc_hd__and3_1 _15230_ (.A(_04579_),
    .B(_04587_),
    .C(_04589_),
    .X(_04591_));
 sky130_fd_sc_hd__a21oi_2 _15231_ (.A1(_04587_),
    .A2(_04589_),
    .B1(_04578_),
    .Y(_04592_));
 sky130_fd_sc_hd__and3_1 _15232_ (.A(_04578_),
    .B(_04587_),
    .C(_04589_),
    .X(_04593_));
 sky130_fd_sc_hd__nor2_1 _15233_ (.A(_04592_),
    .B(_04593_),
    .Y(_04595_));
 sky130_fd_sc_hd__o21ai_2 _15234_ (.A1(_04592_),
    .A2(_04593_),
    .B1(_04575_),
    .Y(_04596_));
 sky130_fd_sc_hd__o2bb2ai_2 _15235_ (.A1_N(_04575_),
    .A2_N(_04577_),
    .B1(_04590_),
    .B2(_04591_),
    .Y(_04597_));
 sky130_fd_sc_hd__o211ai_4 _15236_ (.A1(_04590_),
    .A2(_04591_),
    .B1(_04575_),
    .C1(_04577_),
    .Y(_04598_));
 sky130_fd_sc_hd__o2bb2ai_2 _15237_ (.A1_N(_04575_),
    .A2_N(_04577_),
    .B1(_04592_),
    .B2(_04593_),
    .Y(_04599_));
 sky130_fd_sc_hd__a2bb2o_1 _15238_ (.A1_N(_04421_),
    .A2_N(_04424_),
    .B1(_04423_),
    .B2(_04393_),
    .X(_04600_));
 sky130_fd_sc_hd__a21boi_2 _15239_ (.A1(_04393_),
    .A2(_04423_),
    .B1_N(_04425_),
    .Y(_04601_));
 sky130_fd_sc_hd__nand3_4 _15240_ (.A(_04598_),
    .B(_04599_),
    .C(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__o211a_1 _15241_ (.A1(_04576_),
    .A2(_04596_),
    .B1(_04600_),
    .C1(_04597_),
    .X(_04603_));
 sky130_fd_sc_hd__o211ai_4 _15242_ (.A1(_04576_),
    .A2(_04596_),
    .B1(_04600_),
    .C1(_04597_),
    .Y(_04604_));
 sky130_fd_sc_hd__nand3_1 _15243_ (.A(_04551_),
    .B(_04602_),
    .C(_04604_),
    .Y(_04606_));
 sky130_fd_sc_hd__a21o_1 _15244_ (.A1(_04602_),
    .A2(_04604_),
    .B1(_04551_),
    .X(_04607_));
 sky130_fd_sc_hd__a22o_1 _15245_ (.A1(_04548_),
    .A2(_04549_),
    .B1(_04602_),
    .B2(_04604_),
    .X(_04608_));
 sky130_fd_sc_hd__a31oi_4 _15246_ (.A1(_04598_),
    .A2(_04599_),
    .A3(_04601_),
    .B1(_04551_),
    .Y(_04609_));
 sky130_fd_sc_hd__nand4_2 _15247_ (.A(_04548_),
    .B(_04549_),
    .C(_04602_),
    .D(_04604_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand3_4 _15248_ (.A(_04608_),
    .B(_04610_),
    .C(_04526_),
    .Y(_04611_));
 sky130_fd_sc_hd__o211ai_4 _15249_ (.A1(_04431_),
    .A2(_04525_),
    .B1(_04606_),
    .C1(_04607_),
    .Y(_04612_));
 sky130_fd_sc_hd__o2bb2ai_2 _15250_ (.A1_N(_04347_),
    .A2_N(_04370_),
    .B1(_04367_),
    .B2(_04363_),
    .Y(_04613_));
 sky130_fd_sc_hd__o21ai_1 _15251_ (.A1(_04299_),
    .A2(_04304_),
    .B1(_04307_),
    .Y(_04614_));
 sky130_fd_sc_hd__a22oi_4 _15252_ (.A1(_06541_),
    .A2(net252),
    .B1(_11793_),
    .B2(net30),
    .Y(_04615_));
 sky130_fd_sc_hd__a32o_1 _15253_ (.A1(_06486_),
    .A2(net263),
    .A3(_11771_),
    .B1(_11793_),
    .B2(net30),
    .X(_04617_));
 sky130_fd_sc_hd__or3b_2 _15254_ (.A(net64),
    .B(_03949_),
    .C_N(net63),
    .X(_04618_));
 sky130_fd_sc_hd__o211ai_4 _15255_ (.A1(net263),
    .A2(_08656_),
    .B1(_08250_),
    .C1(_08700_),
    .Y(_04619_));
 sky130_fd_sc_hd__and3_1 _15256_ (.A(_03971_),
    .B(net64),
    .C(net31),
    .X(_04620_));
 sky130_fd_sc_hd__and3_1 _15257_ (.A(_07242_),
    .B(_07253_),
    .C(net289),
    .X(_04621_));
 sky130_fd_sc_hd__a31oi_2 _15258_ (.A1(_07242_),
    .A2(_07253_),
    .A3(net289),
    .B1(_04620_),
    .Y(_04622_));
 sky130_fd_sc_hd__o221ai_2 _15259_ (.A1(_03949_),
    .A2(_08283_),
    .B1(_08711_),
    .B2(_08261_),
    .C1(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__o2bb2ai_4 _15260_ (.A1_N(_04618_),
    .A2_N(_04619_),
    .B1(_04620_),
    .B2(_04621_),
    .Y(_04624_));
 sky130_fd_sc_hd__o2111ai_1 _15261_ (.A1(_03949_),
    .A2(_08283_),
    .B1(_04619_),
    .C1(_04622_),
    .D1(_04615_),
    .Y(_04625_));
 sky130_fd_sc_hd__a31o_2 _15262_ (.A1(_04622_),
    .A2(_04619_),
    .A3(_04618_),
    .B1(_04615_),
    .X(_04626_));
 sky130_fd_sc_hd__nand3_1 _15263_ (.A(_04624_),
    .B(_04625_),
    .C(_04626_),
    .Y(_04628_));
 sky130_fd_sc_hd__a21o_1 _15264_ (.A1(_04623_),
    .A2(_04624_),
    .B1(_04617_),
    .X(_04629_));
 sky130_fd_sc_hd__nand3_1 _15265_ (.A(_04617_),
    .B(_04623_),
    .C(_04624_),
    .Y(_04630_));
 sky130_fd_sc_hd__o2111a_1 _15266_ (.A1(_04624_),
    .A2(_04615_),
    .B1(_04310_),
    .C1(_04307_),
    .D1(_04628_),
    .X(_04631_));
 sky130_fd_sc_hd__o2111ai_4 _15267_ (.A1(_04624_),
    .A2(_04615_),
    .B1(_04310_),
    .C1(_04307_),
    .D1(_04628_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand3_2 _15268_ (.A(_04614_),
    .B(_04629_),
    .C(_04630_),
    .Y(_04633_));
 sky130_fd_sc_hd__a32o_1 _15269_ (.A1(_04998_),
    .A2(net304),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net27),
    .X(_04634_));
 sky130_fd_sc_hd__nor2_1 _15270_ (.A(_03725_),
    .B(_01326_),
    .Y(_04635_));
 sky130_fd_sc_hd__a31oi_1 _15271_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_01293_),
    .B1(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__nor2_1 _15272_ (.A(_03835_),
    .B(_12363_),
    .Y(_04637_));
 sky130_fd_sc_hd__a31oi_1 _15273_ (.A1(_05841_),
    .A2(_05863_),
    .A3(_12330_),
    .B1(_04637_),
    .Y(_04639_));
 sky130_fd_sc_hd__nor2_1 _15274_ (.A(_04636_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__or2_1 _15275_ (.A(_04636_),
    .B(_04639_),
    .X(_04641_));
 sky130_fd_sc_hd__nand2_1 _15276_ (.A(_04636_),
    .B(_04639_),
    .Y(_04642_));
 sky130_fd_sc_hd__and3_1 _15277_ (.A(_04634_),
    .B(_04641_),
    .C(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__nand3_1 _15278_ (.A(_04634_),
    .B(_04641_),
    .C(_04642_),
    .Y(_04644_));
 sky130_fd_sc_hd__a21oi_1 _15279_ (.A1(_04641_),
    .A2(_04642_),
    .B1(_04634_),
    .Y(_04645_));
 sky130_fd_sc_hd__a21o_1 _15280_ (.A1(_04641_),
    .A2(_04642_),
    .B1(_04634_),
    .X(_04646_));
 sky130_fd_sc_hd__nand2_1 _15281_ (.A(_04644_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__o2bb2ai_2 _15282_ (.A1_N(_04632_),
    .A2_N(_04633_),
    .B1(_04643_),
    .B2(_04645_),
    .Y(_04648_));
 sky130_fd_sc_hd__nand4_2 _15283_ (.A(_04632_),
    .B(_04633_),
    .C(_04644_),
    .D(_04646_),
    .Y(_04650_));
 sky130_fd_sc_hd__a21oi_1 _15284_ (.A1(_04648_),
    .A2(_04650_),
    .B1(_04613_),
    .Y(_04651_));
 sky130_fd_sc_hd__a21o_1 _15285_ (.A1(_04648_),
    .A2(_04650_),
    .B1(_04613_),
    .X(_04652_));
 sky130_fd_sc_hd__nand3_2 _15286_ (.A(_04613_),
    .B(_04648_),
    .C(_04650_),
    .Y(_04653_));
 sky130_fd_sc_hd__o21ai_2 _15287_ (.A1(_04312_),
    .A2(_04326_),
    .B1(_04314_),
    .Y(_04654_));
 sky130_fd_sc_hd__inv_2 _15288_ (.A(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__nor2_1 _15289_ (.A(_04655_),
    .B(_04651_),
    .Y(_04656_));
 sky130_fd_sc_hd__and3_1 _15290_ (.A(_04652_),
    .B(_04653_),
    .C(_04654_),
    .X(_04657_));
 sky130_fd_sc_hd__a21oi_2 _15291_ (.A1(_04652_),
    .A2(_04653_),
    .B1(_04654_),
    .Y(_04658_));
 sky130_fd_sc_hd__a21oi_2 _15292_ (.A1(_04652_),
    .A2(_04653_),
    .B1(_04655_),
    .Y(_04659_));
 sky130_fd_sc_hd__and3_1 _15293_ (.A(_04652_),
    .B(_04653_),
    .C(_04655_),
    .X(_04661_));
 sky130_fd_sc_hd__a21oi_1 _15294_ (.A1(_04653_),
    .A2(_04656_),
    .B1(_04658_),
    .Y(_04662_));
 sky130_fd_sc_hd__a21o_1 _15295_ (.A1(_04653_),
    .A2(_04656_),
    .B1(_04658_),
    .X(_04663_));
 sky130_fd_sc_hd__o211ai_2 _15296_ (.A1(_04657_),
    .A2(_04658_),
    .B1(_04611_),
    .C1(_04612_),
    .Y(_04664_));
 sky130_fd_sc_hd__o2bb2ai_1 _15297_ (.A1_N(_04611_),
    .A2_N(_04612_),
    .B1(_04659_),
    .B2(_04661_),
    .Y(_04665_));
 sky130_fd_sc_hd__o2bb2ai_2 _15298_ (.A1_N(_04611_),
    .A2_N(_04612_),
    .B1(_04657_),
    .B2(_04658_),
    .Y(_04666_));
 sky130_fd_sc_hd__o211ai_4 _15299_ (.A1(_04659_),
    .A2(_04661_),
    .B1(_04611_),
    .C1(_04612_),
    .Y(_04667_));
 sky130_fd_sc_hd__a22oi_4 _15300_ (.A1(_04440_),
    .A2(_04523_),
    .B1(_04666_),
    .B2(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__nand4_2 _15301_ (.A(_04438_),
    .B(_04443_),
    .C(_04664_),
    .D(_04665_),
    .Y(_04669_));
 sky130_fd_sc_hd__a22oi_2 _15302_ (.A1(_04438_),
    .A2(_04443_),
    .B1(_04664_),
    .B2(_04665_),
    .Y(_04670_));
 sky130_fd_sc_hd__o211ai_2 _15303_ (.A1(_04437_),
    .A2(_04442_),
    .B1(_04666_),
    .C1(_04667_),
    .Y(_04672_));
 sky130_fd_sc_hd__nand3_1 _15304_ (.A(_04669_),
    .B(_04672_),
    .C(_04522_),
    .Y(_04673_));
 sky130_fd_sc_hd__o22ai_2 _15305_ (.A1(_04519_),
    .A2(_04521_),
    .B1(_04668_),
    .B2(_04670_),
    .Y(_04674_));
 sky130_fd_sc_hd__o211ai_2 _15306_ (.A1(_04519_),
    .A2(_04521_),
    .B1(_04669_),
    .C1(_04672_),
    .Y(_04675_));
 sky130_fd_sc_hd__o21ai_1 _15307_ (.A1(_04668_),
    .A2(_04670_),
    .B1(_04522_),
    .Y(_04676_));
 sky130_fd_sc_hd__o211ai_4 _15308_ (.A1(_04450_),
    .A2(_04478_),
    .B1(_04675_),
    .C1(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__and3_1 _15309_ (.A(_04674_),
    .B(_04479_),
    .C(_04673_),
    .X(_04678_));
 sky130_fd_sc_hd__nand3_1 _15310_ (.A(_04674_),
    .B(_04479_),
    .C(_04673_),
    .Y(_04679_));
 sky130_fd_sc_hd__and3_1 _15311_ (.A(_04291_),
    .B(_04228_),
    .C(_03759_),
    .X(_04680_));
 sky130_fd_sc_hd__a31o_1 _15312_ (.A1(_03759_),
    .A2(_04228_),
    .A3(_04291_),
    .B1(_04288_),
    .X(_04681_));
 sky130_fd_sc_hd__a21oi_1 _15313_ (.A1(_04677_),
    .A2(_04679_),
    .B1(_04681_),
    .Y(_04683_));
 sky130_fd_sc_hd__a21o_1 _15314_ (.A1(_04677_),
    .A2(_04679_),
    .B1(_04681_),
    .X(_04684_));
 sky130_fd_sc_hd__o21ai_2 _15315_ (.A1(_04288_),
    .A2(_04680_),
    .B1(_04677_),
    .Y(_04685_));
 sky130_fd_sc_hd__o211a_1 _15316_ (.A1(_04288_),
    .A2(_04680_),
    .B1(_04679_),
    .C1(_04677_),
    .X(_04686_));
 sky130_fd_sc_hd__o21ai_1 _15317_ (.A1(_04678_),
    .A2(_04685_),
    .B1(_04684_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21a_1 _15318_ (.A1(_04231_),
    .A2(_04457_),
    .B1(_04460_),
    .X(_04688_));
 sky130_fd_sc_hd__o21ai_1 _15319_ (.A1(_04231_),
    .A2(_04457_),
    .B1(_04460_),
    .Y(_04689_));
 sky130_fd_sc_hd__o21ai_1 _15320_ (.A1(_04683_),
    .A2(_04686_),
    .B1(_04688_),
    .Y(_04690_));
 sky130_fd_sc_hd__o211a_1 _15321_ (.A1(_04685_),
    .A2(_04678_),
    .B1(_04684_),
    .C1(_04689_),
    .X(_04691_));
 sky130_fd_sc_hd__o211ai_2 _15322_ (.A1(_04685_),
    .A2(_04678_),
    .B1(_04684_),
    .C1(_04689_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand2_2 _15323_ (.A(_04690_),
    .B(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__a22oi_1 _15324_ (.A1(_04464_),
    .A2(_04468_),
    .B1(_04690_),
    .B2(_04692_),
    .Y(_04695_));
 sky130_fd_sc_hd__a21oi_1 _15325_ (.A1(_04687_),
    .A2(_04688_),
    .B1(_04469_),
    .Y(_04696_));
 sky130_fd_sc_hd__o22ai_2 _15326_ (.A1(_04466_),
    .A2(_04252_),
    .B1(_04696_),
    .B2(_04695_),
    .Y(_04697_));
 sky130_fd_sc_hd__o21ai_1 _15327_ (.A1(_04471_),
    .A2(_04694_),
    .B1(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__o22ai_2 _15328_ (.A1(_04061_),
    .A2(_04250_),
    .B1(_04068_),
    .B2(_04253_),
    .Y(_04699_));
 sky130_fd_sc_hd__a32oi_4 _15329_ (.A1(_04260_),
    .A2(_04476_),
    .A3(_04258_),
    .B1(_04699_),
    .B2(_04473_),
    .Y(_04700_));
 sky130_fd_sc_hd__xor2_1 _15330_ (.A(_04698_),
    .B(_04700_),
    .X(net74));
 sky130_fd_sc_hd__a32oi_2 _15331_ (.A1(_04526_),
    .A2(_04608_),
    .A3(_04610_),
    .B1(_04612_),
    .B2(_04662_),
    .Y(_04701_));
 sky130_fd_sc_hd__a21boi_1 _15332_ (.A1(_04611_),
    .A2(_04663_),
    .B1_N(_04612_),
    .Y(_04702_));
 sky130_fd_sc_hd__o21ai_4 _15333_ (.A1(_04362_),
    .A2(_04544_),
    .B1(_04547_),
    .Y(_04704_));
 sky130_fd_sc_hd__o22a_2 _15334_ (.A1(_05457_),
    .A2(_02869_),
    .B1(_02891_),
    .B2(_03725_),
    .X(_04705_));
 sky130_fd_sc_hd__a32o_1 _15335_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net28),
    .X(_04706_));
 sky130_fd_sc_hd__a32oi_2 _15336_ (.A1(_05841_),
    .A2(_05863_),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net29),
    .Y(_04707_));
 sky130_fd_sc_hd__or3_1 _15337_ (.A(net36),
    .B(_03993_),
    .C(_03916_),
    .X(_04708_));
 sky130_fd_sc_hd__a221o_1 _15338_ (.A1(net306),
    .A2(_06497_),
    .B1(_05863_),
    .B2(net30),
    .C1(_12341_),
    .X(_04709_));
 sky130_fd_sc_hd__a21oi_1 _15339_ (.A1(_04708_),
    .A2(_04709_),
    .B1(_04707_),
    .Y(_04710_));
 sky130_fd_sc_hd__a21o_1 _15340_ (.A1(_04708_),
    .A2(_04709_),
    .B1(_04707_),
    .X(_04711_));
 sky130_fd_sc_hd__o311a_2 _15341_ (.A1(_03916_),
    .A2(_03993_),
    .A3(net36),
    .B1(_04709_),
    .C1(_04707_),
    .X(_04712_));
 sky130_fd_sc_hd__o21a_1 _15342_ (.A1(_04710_),
    .A2(_04712_),
    .B1(_04705_),
    .X(_04713_));
 sky130_fd_sc_hd__nor3_1 _15343_ (.A(_04705_),
    .B(_04710_),
    .C(_04712_),
    .Y(_04715_));
 sky130_fd_sc_hd__o21a_1 _15344_ (.A1(_04710_),
    .A2(_04712_),
    .B1(_04706_),
    .X(_04716_));
 sky130_fd_sc_hd__nor3_1 _15345_ (.A(_04706_),
    .B(_04710_),
    .C(_04712_),
    .Y(_04717_));
 sky130_fd_sc_hd__nor2_1 _15346_ (.A(_04716_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__and3_2 _15347_ (.A(_03993_),
    .B(net34),
    .C(net31),
    .X(_04719_));
 sky130_fd_sc_hd__and3_1 _15348_ (.A(_07242_),
    .B(_07253_),
    .C(net252),
    .X(_04720_));
 sky130_fd_sc_hd__a31oi_4 _15349_ (.A1(_07242_),
    .A2(_07253_),
    .A3(net252),
    .B1(_04719_),
    .Y(_04721_));
 sky130_fd_sc_hd__a32oi_4 _15350_ (.A1(_09698_),
    .A2(net291),
    .A3(net255),
    .B1(_08272_),
    .B2(net2),
    .Y(_04722_));
 sky130_fd_sc_hd__and3_1 _15351_ (.A(_03971_),
    .B(net64),
    .C(net32),
    .X(_04723_));
 sky130_fd_sc_hd__or3b_1 _15352_ (.A(_03949_),
    .B(net34),
    .C_N(net64),
    .X(_04724_));
 sky130_fd_sc_hd__a211o_2 _15353_ (.A1(_06519_),
    .A2(_08645_),
    .B1(_10324_),
    .C1(_08689_),
    .X(_04726_));
 sky130_fd_sc_hd__a31oi_4 _15354_ (.A1(net256),
    .A2(_08700_),
    .A3(net289),
    .B1(_04723_),
    .Y(_04727_));
 sky130_fd_sc_hd__o2111ai_4 _15355_ (.A1(_03949_),
    .A2(_10346_),
    .B1(_04721_),
    .C1(_04726_),
    .D1(_04722_),
    .Y(_04728_));
 sky130_fd_sc_hd__a21o_1 _15356_ (.A1(_04724_),
    .A2(_04726_),
    .B1(_04722_),
    .X(_04729_));
 sky130_fd_sc_hd__o2bb2ai_4 _15357_ (.A1_N(_04722_),
    .A2_N(_04727_),
    .B1(_04719_),
    .B2(_04720_),
    .Y(_04730_));
 sky130_fd_sc_hd__o21ai_2 _15358_ (.A1(_04722_),
    .A2(_04727_),
    .B1(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__o211ai_4 _15359_ (.A1(_04722_),
    .A2(_04727_),
    .B1(_04728_),
    .C1(_04730_),
    .Y(_04732_));
 sky130_fd_sc_hd__a211o_1 _15360_ (.A1(_04724_),
    .A2(_04726_),
    .B1(_04721_),
    .C1(_04722_),
    .X(_04733_));
 sky130_fd_sc_hd__a22oi_4 _15361_ (.A1(_04624_),
    .A2(_04626_),
    .B1(_04732_),
    .B2(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__a22o_1 _15362_ (.A1(_04624_),
    .A2(_04626_),
    .B1(_04732_),
    .B2(_04733_),
    .X(_04735_));
 sky130_fd_sc_hd__o2111a_1 _15363_ (.A1(_04729_),
    .A2(_04721_),
    .B1(_04626_),
    .C1(_04624_),
    .D1(_04732_),
    .X(_04737_));
 sky130_fd_sc_hd__o2111ai_1 _15364_ (.A1(_04729_),
    .A2(_04721_),
    .B1(_04626_),
    .C1(_04624_),
    .D1(_04732_),
    .Y(_04738_));
 sky130_fd_sc_hd__a41o_2 _15365_ (.A1(_04624_),
    .A2(_04626_),
    .A3(_04732_),
    .A4(_04733_),
    .B1(_04718_),
    .X(_04739_));
 sky130_fd_sc_hd__o211ai_2 _15366_ (.A1(_04716_),
    .A2(_04717_),
    .B1(_04735_),
    .C1(_04738_),
    .Y(_04740_));
 sky130_fd_sc_hd__o22ai_4 _15367_ (.A1(_04713_),
    .A2(_04715_),
    .B1(_04734_),
    .B2(_04737_),
    .Y(_04741_));
 sky130_fd_sc_hd__a21oi_2 _15368_ (.A1(_04740_),
    .A2(_04741_),
    .B1(_04704_),
    .Y(_04742_));
 sky130_fd_sc_hd__a21o_1 _15369_ (.A1(_04740_),
    .A2(_04741_),
    .B1(_04704_),
    .X(_04743_));
 sky130_fd_sc_hd__and3_2 _15370_ (.A(_04704_),
    .B(_04740_),
    .C(_04741_),
    .X(_04744_));
 sky130_fd_sc_hd__o211ai_4 _15371_ (.A1(_04734_),
    .A2(_04739_),
    .B1(_04741_),
    .C1(_04704_),
    .Y(_04745_));
 sky130_fd_sc_hd__o21ai_1 _15372_ (.A1(_04647_),
    .A2(_04631_),
    .B1(_04633_),
    .Y(_04746_));
 sky130_fd_sc_hd__o31a_2 _15373_ (.A1(_04631_),
    .A2(_04643_),
    .A3(_04645_),
    .B1(_04633_),
    .X(_04748_));
 sky130_fd_sc_hd__o221a_1 _15374_ (.A1(_04631_),
    .A2(_04647_),
    .B1(_04742_),
    .B2(_04744_),
    .C1(_04633_),
    .X(_04749_));
 sky130_fd_sc_hd__o21ai_1 _15375_ (.A1(_04742_),
    .A2(_04744_),
    .B1(_04748_),
    .Y(_04750_));
 sky130_fd_sc_hd__nor2_1 _15376_ (.A(_04748_),
    .B(_04742_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand2_1 _15377_ (.A(_04743_),
    .B(_04746_),
    .Y(_04752_));
 sky130_fd_sc_hd__and3_1 _15378_ (.A(_04743_),
    .B(_04745_),
    .C(_04746_),
    .X(_04753_));
 sky130_fd_sc_hd__o21a_1 _15379_ (.A1(_04744_),
    .A2(_04752_),
    .B1(_04750_),
    .X(_04754_));
 sky130_fd_sc_hd__o21ai_2 _15380_ (.A1(_04744_),
    .A2(_04752_),
    .B1(_04750_),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _15381_ (.A(_04551_),
    .B(_04604_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_1 _15382_ (.A(_04602_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__o21a_1 _15383_ (.A1(_04590_),
    .A2(_04591_),
    .B1(_04577_),
    .X(_04759_));
 sky130_fd_sc_hd__o21ai_1 _15384_ (.A1(_04595_),
    .A2(_04574_),
    .B1(_04577_),
    .Y(_04760_));
 sky130_fd_sc_hd__or3b_4 _15385_ (.A(net58),
    .B(_04059_),
    .C_N(net55),
    .X(_04761_));
 sky130_fd_sc_hd__nand3_4 _15386_ (.A(_04132_),
    .B(net317),
    .C(_04130_),
    .Y(_04762_));
 sky130_fd_sc_hd__o211ai_4 _15387_ (.A1(_11431_),
    .A2(_03954_),
    .B1(net305),
    .C1(_03952_),
    .Y(_04763_));
 sky130_fd_sc_hd__or3b_4 _15388_ (.A(net59),
    .B(_04048_),
    .C_N(net58),
    .X(_04764_));
 sky130_fd_sc_hd__and4_1 _15389_ (.A(_04761_),
    .B(_04762_),
    .C(_04763_),
    .D(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__o2111ai_4 _15390_ (.A1(_04059_),
    .A2(net316),
    .B1(_04762_),
    .C1(_04763_),
    .D1(_04764_),
    .Y(_04766_));
 sky130_fd_sc_hd__a22oi_4 _15391_ (.A1(net6),
    .A2(_05249_),
    .B1(_02464_),
    .B2(_05227_),
    .Y(_04767_));
 sky130_fd_sc_hd__a32o_1 _15392_ (.A1(_02421_),
    .A2(net249),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net6),
    .X(_04768_));
 sky130_fd_sc_hd__a22oi_4 _15393_ (.A1(_04761_),
    .A2(_04762_),
    .B1(_04763_),
    .B2(_04764_),
    .Y(_04770_));
 sky130_fd_sc_hd__a22o_1 _15394_ (.A1(_04761_),
    .A2(_04762_),
    .B1(_04763_),
    .B2(_04764_),
    .X(_04771_));
 sky130_fd_sc_hd__nor2_1 _15395_ (.A(_04768_),
    .B(_04770_),
    .Y(_04772_));
 sky130_fd_sc_hd__a41oi_4 _15396_ (.A1(_04761_),
    .A2(_04762_),
    .A3(_04763_),
    .A4(_04764_),
    .B1(_04767_),
    .Y(_04773_));
 sky130_fd_sc_hd__a21o_1 _15397_ (.A1(_04766_),
    .A2(_04768_),
    .B1(_04770_),
    .X(_04774_));
 sky130_fd_sc_hd__a221o_1 _15398_ (.A1(_04761_),
    .A2(_04762_),
    .B1(_04763_),
    .B2(_04764_),
    .C1(_04767_),
    .X(_04775_));
 sky130_fd_sc_hd__a21oi_2 _15399_ (.A1(_04766_),
    .A2(_04771_),
    .B1(_04767_),
    .Y(_04776_));
 sky130_fd_sc_hd__and3_1 _15400_ (.A(_04766_),
    .B(_04771_),
    .C(_04767_),
    .X(_04777_));
 sky130_fd_sc_hd__a22oi_4 _15401_ (.A1(_04765_),
    .A2(_04767_),
    .B1(_04775_),
    .B2(_04774_),
    .Y(_04778_));
 sky130_fd_sc_hd__a32oi_4 _15402_ (.A1(net33),
    .A2(_04560_),
    .A3(_04565_),
    .B1(_04568_),
    .B2(_04553_),
    .Y(_04779_));
 sky130_fd_sc_hd__a32o_1 _15403_ (.A1(net33),
    .A2(_04560_),
    .A3(_04565_),
    .B1(_04568_),
    .B2(_04553_),
    .X(_04781_));
 sky130_fd_sc_hd__nor2_1 _15404_ (.A(_04069_),
    .B(_04375_),
    .Y(_04782_));
 sky130_fd_sc_hd__o311a_1 _15405_ (.A1(net7),
    .A2(net249),
    .A3(_04407_),
    .B1(_04342_),
    .C1(net226),
    .X(_04783_));
 sky130_fd_sc_hd__a31oi_4 _15406_ (.A1(net226),
    .A2(_04342_),
    .A3(_04409_),
    .B1(_04782_),
    .Y(_04784_));
 sky130_fd_sc_hd__nor2_2 _15407_ (.A(net10),
    .B(net11),
    .Y(_04785_));
 sky130_fd_sc_hd__nor4_2 _15408_ (.A(net8),
    .B(net9),
    .C(net10),
    .D(net11),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2_8 _15409_ (.A(_04406_),
    .B(_04785_),
    .Y(_04787_));
 sky130_fd_sc_hd__nor3_4 _15410_ (.A(net259),
    .B(net246),
    .C(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand4_4 _15411_ (.A(_06519_),
    .B(net286),
    .C(net283),
    .D(net278),
    .Y(_04789_));
 sky130_fd_sc_hd__o31ai_4 _15412_ (.A1(net263),
    .A2(net245),
    .A3(_04557_),
    .B1(net11),
    .Y(_04790_));
 sky130_fd_sc_hd__a21oi_4 _15413_ (.A1(net186),
    .A2(net11),
    .B1(_04788_),
    .Y(_04792_));
 sky130_fd_sc_hd__o21ai_4 _15414_ (.A1(net232),
    .A2(_04787_),
    .B1(net215),
    .Y(_04793_));
 sky130_fd_sc_hd__nand3_2 _15415_ (.A(_04790_),
    .B(net33),
    .C(net185),
    .Y(_04794_));
 sky130_fd_sc_hd__nand3_2 _15416_ (.A(_04555_),
    .B(_04559_),
    .C(_04484_),
    .Y(_04795_));
 sky130_fd_sc_hd__nor2_2 _15417_ (.A(_04080_),
    .B(_04331_),
    .Y(_04796_));
 sky130_fd_sc_hd__or3_1 _15418_ (.A(net44),
    .B(_04080_),
    .C(_03286_),
    .X(_04797_));
 sky130_fd_sc_hd__and4_1 _15419_ (.A(net185),
    .B(_04790_),
    .C(_04796_),
    .D(net33),
    .X(_04798_));
 sky130_fd_sc_hd__nand4_4 _15420_ (.A(net185),
    .B(_04790_),
    .C(_04796_),
    .D(net33),
    .Y(_04799_));
 sky130_fd_sc_hd__nand2_1 _15421_ (.A(_04794_),
    .B(_04795_),
    .Y(_04800_));
 sky130_fd_sc_hd__o311a_2 _15422_ (.A1(_03286_),
    .A2(net44),
    .A3(_04080_),
    .B1(_04794_),
    .C1(_04795_),
    .X(_04801_));
 sky130_fd_sc_hd__o21ai_2 _15423_ (.A1(_04798_),
    .A2(_04801_),
    .B1(_04784_),
    .Y(_04803_));
 sky130_fd_sc_hd__a31o_1 _15424_ (.A1(net33),
    .A2(_04792_),
    .A3(_04796_),
    .B1(_04784_),
    .X(_04804_));
 sky130_fd_sc_hd__o211ai_2 _15425_ (.A1(_04796_),
    .A2(_04800_),
    .B1(_04799_),
    .C1(_04784_),
    .Y(_04805_));
 sky130_fd_sc_hd__o22ai_2 _15426_ (.A1(_04782_),
    .A2(_04783_),
    .B1(_04798_),
    .B2(_04801_),
    .Y(_04806_));
 sky130_fd_sc_hd__nand3_4 _15427_ (.A(_04806_),
    .B(_04779_),
    .C(_04805_),
    .Y(_04807_));
 sky130_fd_sc_hd__o211a_2 _15428_ (.A1(_04804_),
    .A2(_04801_),
    .B1(_04781_),
    .C1(_04803_),
    .X(_04808_));
 sky130_fd_sc_hd__o211ai_4 _15429_ (.A1(_04804_),
    .A2(_04801_),
    .B1(_04781_),
    .C1(_04803_),
    .Y(_04809_));
 sky130_fd_sc_hd__o211a_4 _15430_ (.A1(_04776_),
    .A2(_04777_),
    .B1(_04807_),
    .C1(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__o211ai_4 _15431_ (.A1(_04776_),
    .A2(_04777_),
    .B1(_04807_),
    .C1(_04809_),
    .Y(_04811_));
 sky130_fd_sc_hd__a21oi_2 _15432_ (.A1(_04807_),
    .A2(_04809_),
    .B1(_04778_),
    .Y(_04812_));
 sky130_fd_sc_hd__a21o_1 _15433_ (.A1(_04807_),
    .A2(_04809_),
    .B1(_04778_),
    .X(_04814_));
 sky130_fd_sc_hd__nand2_1 _15434_ (.A(_04814_),
    .B(_04760_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand3_2 _15435_ (.A(_04814_),
    .B(_04760_),
    .C(_04811_),
    .Y(_04816_));
 sky130_fd_sc_hd__o221a_1 _15436_ (.A1(_04574_),
    .A2(_04595_),
    .B1(_04810_),
    .B2(_04812_),
    .C1(_04577_),
    .X(_04817_));
 sky130_fd_sc_hd__o22ai_4 _15437_ (.A1(_04574_),
    .A2(_04759_),
    .B1(_04810_),
    .B2(_04812_),
    .Y(_04818_));
 sky130_fd_sc_hd__a221o_1 _15438_ (.A1(net2),
    .A2(_07680_),
    .B1(_09709_),
    .B2(_07658_),
    .C1(_04533_),
    .X(_04819_));
 sky130_fd_sc_hd__a21oi_1 _15439_ (.A1(_04527_),
    .A2(_04536_),
    .B1(_04533_),
    .Y(_04820_));
 sky130_fd_sc_hd__o221a_1 _15440_ (.A1(_04015_),
    .A2(_05260_),
    .B1(_00668_),
    .B2(_05238_),
    .C1(_04587_),
    .X(_04821_));
 sky130_fd_sc_hd__o21ai_1 _15441_ (.A1(_04578_),
    .A2(_04588_),
    .B1(_04587_),
    .Y(_04822_));
 sky130_fd_sc_hd__o32a_2 _15442_ (.A1(_11420_),
    .A2(_07669_),
    .A3(_11343_),
    .B1(_07691_),
    .B2(_03982_),
    .X(_04823_));
 sky130_fd_sc_hd__a32o_1 _15443_ (.A1(_11354_),
    .A2(_11431_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net3),
    .X(_04825_));
 sky130_fd_sc_hd__o211ai_2 _15444_ (.A1(_11431_),
    .A2(_00646_),
    .B1(net299),
    .C1(_00625_),
    .Y(_04826_));
 sky130_fd_sc_hd__or3b_1 _15445_ (.A(net61),
    .B(_04015_),
    .C_N(net60),
    .X(_04827_));
 sky130_fd_sc_hd__a32oi_4 _15446_ (.A1(net235),
    .A2(_12999_),
    .A3(net292),
    .B1(_06848_),
    .B2(net4),
    .Y(_04828_));
 sky130_fd_sc_hd__a21oi_2 _15447_ (.A1(_04826_),
    .A2(_04827_),
    .B1(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__a21o_1 _15448_ (.A1(_04826_),
    .A2(_04827_),
    .B1(_04828_),
    .X(_04830_));
 sky130_fd_sc_hd__o211a_1 _15449_ (.A1(_04015_),
    .A2(net298),
    .B1(_04826_),
    .C1(_04828_),
    .X(_04831_));
 sky130_fd_sc_hd__o221ai_4 _15450_ (.A1(_04015_),
    .A2(net298),
    .B1(_00668_),
    .B2(_05699_),
    .C1(_04828_),
    .Y(_04832_));
 sky130_fd_sc_hd__a21oi_1 _15451_ (.A1(_04830_),
    .A2(_04832_),
    .B1(_04825_),
    .Y(_04833_));
 sky130_fd_sc_hd__o21ai_1 _15452_ (.A1(_04829_),
    .A2(_04831_),
    .B1(_04823_),
    .Y(_04834_));
 sky130_fd_sc_hd__nor3_1 _15453_ (.A(_04823_),
    .B(_04829_),
    .C(_04831_),
    .Y(_04836_));
 sky130_fd_sc_hd__nand3_1 _15454_ (.A(_04825_),
    .B(_04830_),
    .C(_04832_),
    .Y(_04837_));
 sky130_fd_sc_hd__nand3_2 _15455_ (.A(_04822_),
    .B(_04834_),
    .C(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21oi_1 _15456_ (.A1(_04834_),
    .A2(_04837_),
    .B1(_04822_),
    .Y(_04839_));
 sky130_fd_sc_hd__o22ai_2 _15457_ (.A1(_04588_),
    .A2(_04821_),
    .B1(_04833_),
    .B2(_04836_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_1 _15458_ (.A(_04820_),
    .B(_04839_),
    .Y(_04841_));
 sky130_fd_sc_hd__nand4_1 _15459_ (.A(_04536_),
    .B(_04819_),
    .C(_04838_),
    .D(_04840_),
    .Y(_04842_));
 sky130_fd_sc_hd__inv_2 _15460_ (.A(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__a22oi_4 _15461_ (.A1(_04536_),
    .A2(_04819_),
    .B1(_04838_),
    .B2(_04840_),
    .Y(_04844_));
 sky130_fd_sc_hd__a21oi_2 _15462_ (.A1(_04841_),
    .A2(_04838_),
    .B1(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__a21bo_1 _15463_ (.A1(_04816_),
    .A2(_04818_),
    .B1_N(_04845_),
    .X(_04847_));
 sky130_fd_sc_hd__o221ai_4 _15464_ (.A1(_04810_),
    .A2(_04815_),
    .B1(_04843_),
    .B2(_04844_),
    .C1(_04818_),
    .Y(_04848_));
 sky130_fd_sc_hd__o2bb2ai_4 _15465_ (.A1_N(_04816_),
    .A2_N(_04818_),
    .B1(_04843_),
    .B2(_04844_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_1 _15466_ (.A(_04816_),
    .B(_04845_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand3_1 _15467_ (.A(_04816_),
    .B(_04818_),
    .C(_04845_),
    .Y(_04851_));
 sky130_fd_sc_hd__a22oi_4 _15468_ (.A1(_04602_),
    .A2(_04756_),
    .B1(_04849_),
    .B2(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__nand3_1 _15469_ (.A(_04757_),
    .B(_04847_),
    .C(_04848_),
    .Y(_04853_));
 sky130_fd_sc_hd__o221a_2 _15470_ (.A1(_04603_),
    .A2(_04609_),
    .B1(_04817_),
    .B2(_04850_),
    .C1(_04849_),
    .X(_04854_));
 sky130_fd_sc_hd__o221ai_4 _15471_ (.A1(_04603_),
    .A2(_04609_),
    .B1(_04817_),
    .B2(_04850_),
    .C1(_04849_),
    .Y(_04855_));
 sky130_fd_sc_hd__o211ai_1 _15472_ (.A1(_04749_),
    .A2(_04753_),
    .B1(_04853_),
    .C1(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__o21ai_1 _15473_ (.A1(_04852_),
    .A2(_04854_),
    .B1(_04754_),
    .Y(_04858_));
 sky130_fd_sc_hd__o22ai_1 _15474_ (.A1(_04749_),
    .A2(_04753_),
    .B1(_04852_),
    .B2(_04854_),
    .Y(_04859_));
 sky130_fd_sc_hd__a31oi_2 _15475_ (.A1(_04757_),
    .A2(_04847_),
    .A3(_04848_),
    .B1(_04755_),
    .Y(_04860_));
 sky130_fd_sc_hd__nand3_1 _15476_ (.A(_04853_),
    .B(_04855_),
    .C(_04754_),
    .Y(_04861_));
 sky130_fd_sc_hd__nand3_2 _15477_ (.A(_04858_),
    .B(_04701_),
    .C(_04856_),
    .Y(_04862_));
 sky130_fd_sc_hd__nand3_2 _15478_ (.A(_04702_),
    .B(_04859_),
    .C(_04861_),
    .Y(_04863_));
 sky130_fd_sc_hd__nand2_1 _15479_ (.A(_04511_),
    .B(_04513_),
    .Y(_04864_));
 sky130_fd_sc_hd__a31o_1 _15480_ (.A1(_04613_),
    .A2(_04648_),
    .A3(_04650_),
    .B1(_04654_),
    .X(_04865_));
 sky130_fd_sc_hd__o21ai_1 _15481_ (.A1(_04487_),
    .A2(_04493_),
    .B1(_04497_),
    .Y(_04866_));
 sky130_fd_sc_hd__a21oi_1 _15482_ (.A1(_04634_),
    .A2(_04642_),
    .B1(_04640_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21o_1 _15483_ (.A1(_04634_),
    .A2(_04642_),
    .B1(_04640_),
    .X(_04869_));
 sky130_fd_sc_hd__nor2_1 _15484_ (.A(_03396_),
    .B(_04270_),
    .Y(_04870_));
 sky130_fd_sc_hd__and3_1 _15485_ (.A(net318),
    .B(_04452_),
    .C(net280),
    .X(_04871_));
 sky130_fd_sc_hd__a31o_1 _15486_ (.A1(net318),
    .A2(_04452_),
    .A3(net280),
    .B1(_04870_),
    .X(_04872_));
 sky130_fd_sc_hd__or3_1 _15487_ (.A(net39),
    .B(_04037_),
    .C(_03616_),
    .X(_04873_));
 sky130_fd_sc_hd__nand4_4 _15488_ (.A(_04037_),
    .B(net304),
    .C(net39),
    .D(_04998_),
    .Y(_04874_));
 sky130_fd_sc_hd__a211oi_2 _15489_ (.A1(_04397_),
    .A2(_04725_),
    .B1(_04216_),
    .C1(_04703_),
    .Y(_04875_));
 sky130_fd_sc_hd__nor2_1 _15490_ (.A(_03506_),
    .B(_04218_),
    .Y(_04876_));
 sky130_fd_sc_hd__a31oi_2 _15491_ (.A1(net315),
    .A2(net267),
    .A3(_04215_),
    .B1(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__o2bb2a_1 _15492_ (.A1_N(_04873_),
    .A2_N(_04874_),
    .B1(_04875_),
    .B2(_04876_),
    .X(_04878_));
 sky130_fd_sc_hd__o2bb2ai_4 _15493_ (.A1_N(_04873_),
    .A2_N(_04874_),
    .B1(_04875_),
    .B2(_04876_),
    .Y(_04879_));
 sky130_fd_sc_hd__o211ai_4 _15494_ (.A1(_03616_),
    .A2(_03737_),
    .B1(_04874_),
    .C1(_04877_),
    .Y(_04880_));
 sky130_fd_sc_hd__a21oi_1 _15495_ (.A1(_04879_),
    .A2(_04880_),
    .B1(_04872_),
    .Y(_04881_));
 sky130_fd_sc_hd__a21o_1 _15496_ (.A1(_04879_),
    .A2(_04880_),
    .B1(_04872_),
    .X(_04882_));
 sky130_fd_sc_hd__o211a_1 _15497_ (.A1(_04870_),
    .A2(_04871_),
    .B1(_04879_),
    .C1(_04880_),
    .X(_04883_));
 sky130_fd_sc_hd__o211ai_4 _15498_ (.A1(_04870_),
    .A2(_04871_),
    .B1(_04879_),
    .C1(_04880_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand3_4 _15499_ (.A(_04869_),
    .B(_04882_),
    .C(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21ai_2 _15500_ (.A1(_04881_),
    .A2(_04883_),
    .B1(_04867_),
    .Y(_04886_));
 sky130_fd_sc_hd__a21oi_1 _15501_ (.A1(_04885_),
    .A2(_04886_),
    .B1(_04866_),
    .Y(_04887_));
 sky130_fd_sc_hd__a21o_1 _15502_ (.A1(_04885_),
    .A2(_04886_),
    .B1(_04866_),
    .X(_04888_));
 sky130_fd_sc_hd__o211a_1 _15503_ (.A1(_04496_),
    .A2(_04499_),
    .B1(_04885_),
    .C1(_04886_),
    .X(_04890_));
 sky130_fd_sc_hd__o211ai_1 _15504_ (.A1(_04496_),
    .A2(_04499_),
    .B1(_04885_),
    .C1(_04886_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_1 _15505_ (.A1(_04505_),
    .A2(_04501_),
    .B1(_04503_),
    .Y(_04892_));
 sky130_fd_sc_hd__o21bai_2 _15506_ (.A1(_04887_),
    .A2(_04890_),
    .B1_N(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand3_1 _15507_ (.A(_04888_),
    .B(_04891_),
    .C(_04892_),
    .Y(_04894_));
 sky130_fd_sc_hd__nor2_8 _15508_ (.A(net42),
    .B(_04102_),
    .Y(_04895_));
 sky130_fd_sc_hd__nand2b_4 _15509_ (.A_N(net42),
    .B(net43),
    .Y(_04896_));
 sky130_fd_sc_hd__and2b_4 _15510_ (.A_N(net43),
    .B(net42),
    .X(_04897_));
 sky130_fd_sc_hd__nand2_8 _15511_ (.A(_04102_),
    .B(net42),
    .Y(_04898_));
 sky130_fd_sc_hd__a21oi_1 _15512_ (.A1(_04896_),
    .A2(_04898_),
    .B1(_03176_),
    .Y(_04899_));
 sky130_fd_sc_hd__a22o_1 _15513_ (.A1(net12),
    .A2(_04482_),
    .B1(_04539_),
    .B2(net279),
    .X(_04901_));
 sky130_fd_sc_hd__o211a_1 _15514_ (.A1(net243),
    .A2(_04897_),
    .B1(net1),
    .C1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__nor2_1 _15515_ (.A(_04899_),
    .B(_04901_),
    .Y(_04903_));
 sky130_fd_sc_hd__nor2_1 _15516_ (.A(_04902_),
    .B(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__a21oi_1 _15517_ (.A1(_04893_),
    .A2(_04894_),
    .B1(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21o_1 _15518_ (.A1(_04893_),
    .A2(_04894_),
    .B1(_04904_),
    .X(_04906_));
 sky130_fd_sc_hd__and3_1 _15519_ (.A(_04893_),
    .B(_04894_),
    .C(_04904_),
    .X(_04907_));
 sky130_fd_sc_hd__nand3_1 _15520_ (.A(_04893_),
    .B(_04894_),
    .C(_04904_),
    .Y(_04908_));
 sky130_fd_sc_hd__o2bb2ai_1 _15521_ (.A1_N(_04652_),
    .A2_N(_04865_),
    .B1(_04905_),
    .B2(_04907_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand4_1 _15522_ (.A(_04652_),
    .B(_04865_),
    .C(_04906_),
    .D(_04908_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand2_1 _15523_ (.A(_04909_),
    .B(_04910_),
    .Y(_04912_));
 sky130_fd_sc_hd__and3_1 _15524_ (.A(_04511_),
    .B(_04513_),
    .C(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__and3_1 _15525_ (.A(_04864_),
    .B(_04909_),
    .C(_04910_),
    .X(_04914_));
 sky130_fd_sc_hd__xnor2_1 _15526_ (.A(_04864_),
    .B(_04912_),
    .Y(_04915_));
 sky130_fd_sc_hd__o2bb2ai_1 _15527_ (.A1_N(_04862_),
    .A2_N(_04863_),
    .B1(_04913_),
    .B2(_04914_),
    .Y(_04916_));
 sky130_fd_sc_hd__nand3_2 _15528_ (.A(_04862_),
    .B(_04915_),
    .C(_04863_),
    .Y(_04917_));
 sky130_fd_sc_hd__o21a_1 _15529_ (.A1(_04519_),
    .A2(_04521_),
    .B1(_04672_),
    .X(_04918_));
 sky130_fd_sc_hd__a31o_1 _15530_ (.A1(_04524_),
    .A2(_04666_),
    .A3(_04667_),
    .B1(_04522_),
    .X(_04919_));
 sky130_fd_sc_hd__o2bb2ai_2 _15531_ (.A1_N(_04916_),
    .A2_N(_04917_),
    .B1(_04918_),
    .B2(_04668_),
    .Y(_04920_));
 sky130_fd_sc_hd__nand4_2 _15532_ (.A(_04669_),
    .B(_04916_),
    .C(_04917_),
    .D(_04919_),
    .Y(_04921_));
 sky130_fd_sc_hd__a31o_1 _15533_ (.A1(_04226_),
    .A2(_04518_),
    .A3(_04283_),
    .B1(_04515_),
    .X(_04923_));
 sky130_fd_sc_hd__a21oi_1 _15534_ (.A1(_04920_),
    .A2(_04921_),
    .B1(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__o211a_1 _15535_ (.A1(_04515_),
    .A2(_04521_),
    .B1(_04920_),
    .C1(_04921_),
    .X(_04925_));
 sky130_fd_sc_hd__o211ai_2 _15536_ (.A1(_04515_),
    .A2(_04521_),
    .B1(_04920_),
    .C1(_04921_),
    .Y(_04926_));
 sky130_fd_sc_hd__a32o_1 _15537_ (.A1(_04479_),
    .A2(_04673_),
    .A3(_04674_),
    .B1(_04677_),
    .B2(_04681_),
    .X(_04927_));
 sky130_fd_sc_hd__o21bai_2 _15538_ (.A1(_04924_),
    .A2(_04925_),
    .B1_N(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__a211oi_1 _15539_ (.A1(_04679_),
    .A2(_04685_),
    .B1(_04924_),
    .C1(_04925_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand3b_2 _15540_ (.A_N(_04924_),
    .B(_04926_),
    .C(_04927_),
    .Y(_04930_));
 sky130_fd_sc_hd__o2bb2ai_2 _15541_ (.A1_N(_04928_),
    .A2_N(_04930_),
    .B1(_04687_),
    .B2(_04688_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand3_2 _15542_ (.A(_04928_),
    .B(_04930_),
    .C(_04691_),
    .Y(_04932_));
 sky130_fd_sc_hd__o2bb2ai_2 _15543_ (.A1_N(_04931_),
    .A2_N(_04932_),
    .B1(_04469_),
    .B2(_04694_),
    .Y(_04934_));
 sky130_fd_sc_hd__a21bo_1 _15544_ (.A1(_04696_),
    .A2(_04931_),
    .B1_N(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__o22a_1 _15545_ (.A1(_04471_),
    .A2(_04694_),
    .B1(_04698_),
    .B2(_04700_),
    .X(_04936_));
 sky130_fd_sc_hd__xor2_1 _15546_ (.A(_04935_),
    .B(_04936_),
    .X(net75));
 sky130_fd_sc_hd__o311a_1 _15547_ (.A1(_04252_),
    .A2(_04466_),
    .A3(_04694_),
    .B1(_04697_),
    .C1(_04934_),
    .X(_04937_));
 sky130_fd_sc_hd__nand4_4 _15548_ (.A(_04937_),
    .B(_04257_),
    .C(_04255_),
    .D(_04476_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21oi_4 _15549_ (.A1(_04066_),
    .A2(_04259_),
    .B1(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand3_1 _15550_ (.A(_04473_),
    .B(_04697_),
    .C(_04699_),
    .Y(_04940_));
 sky130_fd_sc_hd__a2bb2oi_1 _15551_ (.A1_N(_04471_),
    .A2_N(_04694_),
    .B1(_04696_),
    .B2(_04931_),
    .Y(_04941_));
 sky130_fd_sc_hd__nand2_1 _15552_ (.A(_04940_),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__a21o_1 _15553_ (.A1(_04934_),
    .A2(_04942_),
    .B1(_04939_),
    .X(_04944_));
 sky130_fd_sc_hd__a21boi_1 _15554_ (.A1(_04920_),
    .A2(_04923_),
    .B1_N(_04921_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _15555_ (.A(_04921_),
    .B(_04926_),
    .Y(_04946_));
 sky130_fd_sc_hd__a21boi_2 _15556_ (.A1(_04864_),
    .A2(_04909_),
    .B1_N(_04910_),
    .Y(_04947_));
 sky130_fd_sc_hd__inv_2 _15557_ (.A(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__a21boi_2 _15558_ (.A1(_04862_),
    .A2(_04915_),
    .B1_N(_04863_),
    .Y(_04949_));
 sky130_fd_sc_hd__nand2_1 _15559_ (.A(_04863_),
    .B(_04917_),
    .Y(_04950_));
 sky130_fd_sc_hd__a21bo_1 _15560_ (.A1(_04893_),
    .A2(_04904_),
    .B1_N(_04894_),
    .X(_04951_));
 sky130_fd_sc_hd__a21oi_2 _15561_ (.A1(_04872_),
    .A2(_04880_),
    .B1(_04878_),
    .Y(_04952_));
 sky130_fd_sc_hd__a32o_1 _15562_ (.A1(net315),
    .A2(net267),
    .A3(net280),
    .B1(_04269_),
    .B2(net26),
    .X(_04953_));
 sky130_fd_sc_hd__nor2_1 _15563_ (.A(_03616_),
    .B(_04218_),
    .Y(_04955_));
 sky130_fd_sc_hd__a31oi_2 _15564_ (.A1(net266),
    .A2(net303),
    .A3(_04215_),
    .B1(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__a31o_1 _15565_ (.A1(net266),
    .A2(net303),
    .A3(_04215_),
    .B1(_04955_),
    .X(_04957_));
 sky130_fd_sc_hd__nor2_1 _15566_ (.A(_03725_),
    .B(_03737_),
    .Y(_04958_));
 sky130_fd_sc_hd__a31o_1 _15567_ (.A1(_05414_),
    .A2(_05446_),
    .A3(net285),
    .B1(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__nand2_1 _15568_ (.A(_04957_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__inv_2 _15569_ (.A(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__o221ai_4 _15570_ (.A1(_05457_),
    .A2(_03714_),
    .B1(_03737_),
    .B2(_03725_),
    .C1(_04956_),
    .Y(_04962_));
 sky130_fd_sc_hd__nand2_1 _15571_ (.A(_04959_),
    .B(_04956_),
    .Y(_04963_));
 sky130_fd_sc_hd__o221ai_2 _15572_ (.A1(_05457_),
    .A2(_03714_),
    .B1(_03737_),
    .B2(_03725_),
    .C1(_04957_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand3_2 _15573_ (.A(_04953_),
    .B(_04960_),
    .C(_04962_),
    .Y(_04966_));
 sky130_fd_sc_hd__inv_2 _15574_ (.A(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand3b_1 _15575_ (.A_N(_04953_),
    .B(_04963_),
    .C(_04964_),
    .Y(_04968_));
 sky130_fd_sc_hd__nand3b_2 _15576_ (.A_N(_04953_),
    .B(_04960_),
    .C(_04962_),
    .Y(_04969_));
 sky130_fd_sc_hd__nand3_1 _15577_ (.A(_04953_),
    .B(_04963_),
    .C(_04964_),
    .Y(_04970_));
 sky130_fd_sc_hd__o21ai_1 _15578_ (.A1(_04705_),
    .A2(_04712_),
    .B1(_04711_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand3_4 _15579_ (.A(_04971_),
    .B(_04968_),
    .C(_04966_),
    .Y(_04972_));
 sky130_fd_sc_hd__o2111a_1 _15580_ (.A1(_04705_),
    .A2(_04712_),
    .B1(_04969_),
    .C1(_04970_),
    .D1(_04711_),
    .X(_04973_));
 sky130_fd_sc_hd__o2111ai_4 _15581_ (.A1(_04705_),
    .A2(_04712_),
    .B1(_04969_),
    .C1(_04970_),
    .D1(_04711_),
    .Y(_04974_));
 sky130_fd_sc_hd__a21bo_1 _15582_ (.A1(_04972_),
    .A2(_04974_),
    .B1_N(_04952_),
    .X(_04975_));
 sky130_fd_sc_hd__o211ai_2 _15583_ (.A1(_04878_),
    .A2(_04883_),
    .B1(_04972_),
    .C1(_04974_),
    .Y(_04977_));
 sky130_fd_sc_hd__nand4_2 _15584_ (.A(_04879_),
    .B(_04884_),
    .C(_04972_),
    .D(_04974_),
    .Y(_04978_));
 sky130_fd_sc_hd__a22o_1 _15585_ (.A1(_04879_),
    .A2(_04884_),
    .B1(_04972_),
    .B2(_04974_),
    .X(_04979_));
 sky130_fd_sc_hd__o21ai_2 _15586_ (.A1(_04496_),
    .A2(_04499_),
    .B1(_04886_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2_1 _15587_ (.A(_04885_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand4_4 _15588_ (.A(_04885_),
    .B(_04978_),
    .C(_04979_),
    .D(_04980_),
    .Y(_04982_));
 sky130_fd_sc_hd__and3_2 _15589_ (.A(_04975_),
    .B(_04981_),
    .C(_04977_),
    .X(_04983_));
 sky130_fd_sc_hd__nand3_1 _15590_ (.A(_04975_),
    .B(_04981_),
    .C(_04977_),
    .Y(_04984_));
 sky130_fd_sc_hd__nor2_8 _15591_ (.A(net43),
    .B(_04124_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_8 _15592_ (.A(_04102_),
    .B(net45),
    .Y(_04986_));
 sky130_fd_sc_hd__nor2_8 _15593_ (.A(net45),
    .B(_04102_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand2_8 _15594_ (.A(_04124_),
    .B(net43),
    .Y(_04989_));
 sky130_fd_sc_hd__a21oi_1 _15595_ (.A1(_04986_),
    .A2(_04989_),
    .B1(_03176_),
    .Y(_04990_));
 sky130_fd_sc_hd__a22oi_2 _15596_ (.A1(net12),
    .A2(_04897_),
    .B1(_04539_),
    .B2(net243),
    .Y(_04991_));
 sky130_fd_sc_hd__a211o_1 _15597_ (.A1(_03176_),
    .A2(_04430_),
    .B1(_04481_),
    .C1(_04408_),
    .X(_04992_));
 sky130_fd_sc_hd__or3b_1 _15598_ (.A(_03396_),
    .B(net42),
    .C_N(net41),
    .X(_04993_));
 sky130_fd_sc_hd__o32a_1 _15599_ (.A1(_04481_),
    .A2(_04441_),
    .A3(_04408_),
    .B1(_03396_),
    .B2(_04483_),
    .X(_04994_));
 sky130_fd_sc_hd__a21oi_1 _15600_ (.A1(_04992_),
    .A2(_04993_),
    .B1(_04991_),
    .Y(_04995_));
 sky130_fd_sc_hd__a21o_1 _15601_ (.A1(_04992_),
    .A2(_04993_),
    .B1(_04991_),
    .X(_04996_));
 sky130_fd_sc_hd__nand2_1 _15602_ (.A(_04991_),
    .B(_04994_),
    .Y(_04997_));
 sky130_fd_sc_hd__a21oi_1 _15603_ (.A1(_04996_),
    .A2(_04997_),
    .B1(_04990_),
    .Y(_04999_));
 sky130_fd_sc_hd__and3_1 _15604_ (.A(_04996_),
    .B(_04997_),
    .C(_04990_),
    .X(_05000_));
 sky130_fd_sc_hd__o2bb2a_1 _15605_ (.A1_N(_04899_),
    .A2_N(_04901_),
    .B1(_04999_),
    .B2(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__or3b_2 _15606_ (.A(_04999_),
    .B(_05000_),
    .C_N(_04902_),
    .X(_05002_));
 sky130_fd_sc_hd__and2b_1 _15607_ (.A_N(_05001_),
    .B(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__a21o_1 _15608_ (.A1(_04982_),
    .A2(_04984_),
    .B1(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__and2_1 _15609_ (.A(_05003_),
    .B(_04982_),
    .X(_05005_));
 sky130_fd_sc_hd__nand2_1 _15610_ (.A(_05003_),
    .B(_04982_),
    .Y(_05006_));
 sky130_fd_sc_hd__o21ai_1 _15611_ (.A1(_04983_),
    .A2(_05006_),
    .B1(_05004_),
    .Y(_05007_));
 sky130_fd_sc_hd__o211ai_4 _15612_ (.A1(_04748_),
    .A2(_04742_),
    .B1(_04745_),
    .C1(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__o221ai_4 _15613_ (.A1(_04983_),
    .A2(_05006_),
    .B1(_04744_),
    .B2(_04751_),
    .C1(_05004_),
    .Y(_05010_));
 sky130_fd_sc_hd__a21oi_2 _15614_ (.A1(_05008_),
    .A2(_05010_),
    .B1(_04951_),
    .Y(_05011_));
 sky130_fd_sc_hd__a21o_1 _15615_ (.A1(_05008_),
    .A2(_05010_),
    .B1(_04951_),
    .X(_05012_));
 sky130_fd_sc_hd__and3_1 _15616_ (.A(_05010_),
    .B(_04951_),
    .C(_05008_),
    .X(_05013_));
 sky130_fd_sc_hd__nand3_2 _15617_ (.A(_05010_),
    .B(_04951_),
    .C(_05008_),
    .Y(_05014_));
 sky130_fd_sc_hd__nor2_1 _15618_ (.A(_05011_),
    .B(_05013_),
    .Y(_05015_));
 sky130_fd_sc_hd__nand2_2 _15619_ (.A(_05012_),
    .B(_05014_),
    .Y(_05016_));
 sky130_fd_sc_hd__a32o_1 _15620_ (.A1(_05841_),
    .A2(net265),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net29),
    .X(_05017_));
 sky130_fd_sc_hd__or3b_1 _15621_ (.A(_03916_),
    .B(net37),
    .C_N(net36),
    .X(_05018_));
 sky130_fd_sc_hd__o211ai_4 _15622_ (.A1(_04747_),
    .A2(net264),
    .B1(_01293_),
    .C1(_06486_),
    .Y(_05019_));
 sky130_fd_sc_hd__or3_2 _15623_ (.A(net36),
    .B(_03993_),
    .C(_03938_),
    .X(_05021_));
 sky130_fd_sc_hd__nand3_2 _15624_ (.A(_07242_),
    .B(_07253_),
    .C(_12330_),
    .Y(_05022_));
 sky130_fd_sc_hd__a22oi_4 _15625_ (.A1(_05018_),
    .A2(_05019_),
    .B1(_05021_),
    .B2(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__o2111a_1 _15626_ (.A1(_03916_),
    .A2(_01326_),
    .B1(_05019_),
    .C1(_05021_),
    .D1(_05022_),
    .X(_05024_));
 sky130_fd_sc_hd__o2111ai_1 _15627_ (.A1(_03916_),
    .A2(_01326_),
    .B1(_05019_),
    .C1(_05021_),
    .D1(_05022_),
    .Y(_05025_));
 sky130_fd_sc_hd__nor2_1 _15628_ (.A(_05023_),
    .B(_05024_),
    .Y(_05026_));
 sky130_fd_sc_hd__and2_1 _15629_ (.A(_05026_),
    .B(_05017_),
    .X(_05027_));
 sky130_fd_sc_hd__nor2_1 _15630_ (.A(_05017_),
    .B(_05026_),
    .Y(_05028_));
 sky130_fd_sc_hd__o21a_1 _15631_ (.A1(_05023_),
    .A2(_05024_),
    .B1(_05017_),
    .X(_05029_));
 sky130_fd_sc_hd__nor3_1 _15632_ (.A(_05017_),
    .B(_05023_),
    .C(_05024_),
    .Y(_05030_));
 sky130_fd_sc_hd__o32a_2 _15633_ (.A1(_11782_),
    .A2(_08689_),
    .A3(_08667_),
    .B1(_03949_),
    .B2(_11804_),
    .X(_05032_));
 sky130_fd_sc_hd__a32o_1 _15634_ (.A1(net256),
    .A2(_08700_),
    .A3(net252),
    .B1(_11793_),
    .B2(net32),
    .X(_05033_));
 sky130_fd_sc_hd__a31oi_4 _15635_ (.A1(net311),
    .A2(net295),
    .A3(net290),
    .B1(_10324_),
    .Y(_05034_));
 sky130_fd_sc_hd__a22oi_4 _15636_ (.A1(net2),
    .A2(_10335_),
    .B1(_09698_),
    .B2(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__o211ai_1 _15637_ (.A1(net261),
    .A2(_11387_),
    .B1(net291),
    .C1(_11354_),
    .Y(_05036_));
 sky130_fd_sc_hd__or3b_1 _15638_ (.A(net64),
    .B(_03982_),
    .C_N(net63),
    .X(_05037_));
 sky130_fd_sc_hd__a21oi_1 _15639_ (.A1(_05036_),
    .A2(_05037_),
    .B1(_05035_),
    .Y(_05038_));
 sky130_fd_sc_hd__a21o_1 _15640_ (.A1(_05036_),
    .A2(_05037_),
    .B1(_05035_),
    .X(_05039_));
 sky130_fd_sc_hd__o221a_2 _15641_ (.A1(_03982_),
    .A2(_08283_),
    .B1(net236),
    .B2(_08261_),
    .C1(_05035_),
    .X(_05040_));
 sky130_fd_sc_hd__o221ai_4 _15642_ (.A1(_03982_),
    .A2(_08283_),
    .B1(net236),
    .B2(_08261_),
    .C1(_05035_),
    .Y(_05041_));
 sky130_fd_sc_hd__o21ai_2 _15643_ (.A1(_05038_),
    .A2(_05040_),
    .B1(_05033_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand3_2 _15644_ (.A(_05039_),
    .B(_05041_),
    .C(_05032_),
    .Y(_05044_));
 sky130_fd_sc_hd__a21oi_1 _15645_ (.A1(_05033_),
    .A2(_05041_),
    .B1(_05038_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand3_1 _15646_ (.A(_05033_),
    .B(_05039_),
    .C(_05041_),
    .Y(_05046_));
 sky130_fd_sc_hd__o21ai_1 _15647_ (.A1(_05038_),
    .A2(_05040_),
    .B1(_05032_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_1 _15648_ (.A(_05043_),
    .B(_05044_),
    .Y(_05048_));
 sky130_fd_sc_hd__a22oi_4 _15649_ (.A1(_04729_),
    .A2(_04730_),
    .B1(_05043_),
    .B2(_05044_),
    .Y(_05049_));
 sky130_fd_sc_hd__a22o_1 _15650_ (.A1(_04729_),
    .A2(_04730_),
    .B1(_05043_),
    .B2(_05044_),
    .X(_05050_));
 sky130_fd_sc_hd__a21oi_1 _15651_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_04731_),
    .Y(_05051_));
 sky130_fd_sc_hd__a21o_1 _15652_ (.A1(_05046_),
    .A2(_05047_),
    .B1(_04731_),
    .X(_05052_));
 sky130_fd_sc_hd__o22ai_4 _15653_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_04731_),
    .B2(_05048_),
    .Y(_05054_));
 sky130_fd_sc_hd__o211ai_1 _15654_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_05050_),
    .C1(_05052_),
    .Y(_05055_));
 sky130_fd_sc_hd__o22ai_2 _15655_ (.A1(_05027_),
    .A2(_05028_),
    .B1(_05049_),
    .B2(_05051_),
    .Y(_05056_));
 sky130_fd_sc_hd__o21ai_2 _15656_ (.A1(_05049_),
    .A2(_05054_),
    .B1(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__o21a_1 _15657_ (.A1(_04820_),
    .A2(_04839_),
    .B1(_04838_),
    .X(_05058_));
 sky130_fd_sc_hd__o21ai_1 _15658_ (.A1(_04820_),
    .A2(_04839_),
    .B1(_04838_),
    .Y(_05059_));
 sky130_fd_sc_hd__a21oi_1 _15659_ (.A1(_05055_),
    .A2(_05056_),
    .B1(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__o211a_2 _15660_ (.A1(_05049_),
    .A2(_05054_),
    .B1(_05056_),
    .C1(_05059_),
    .X(_05061_));
 sky130_fd_sc_hd__o21ai_1 _15661_ (.A1(_04718_),
    .A2(_04737_),
    .B1(_04735_),
    .Y(_05062_));
 sky130_fd_sc_hd__o21bai_2 _15662_ (.A1(_05060_),
    .A2(_05061_),
    .B1_N(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__a22oi_4 _15663_ (.A1(_04735_),
    .A2(_04739_),
    .B1(_05057_),
    .B2(_05058_),
    .Y(_05065_));
 sky130_fd_sc_hd__o21ai_2 _15664_ (.A1(_05057_),
    .A2(_05058_),
    .B1(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__nand2_2 _15665_ (.A(_05063_),
    .B(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__o2bb2ai_1 _15666_ (.A1_N(_04845_),
    .A2_N(_04818_),
    .B1(_04815_),
    .B2(_04810_),
    .Y(_05068_));
 sky130_fd_sc_hd__a21boi_2 _15667_ (.A1(_04818_),
    .A2(_04845_),
    .B1_N(_04816_),
    .Y(_05069_));
 sky130_fd_sc_hd__a21oi_4 _15668_ (.A1(_04778_),
    .A2(_04807_),
    .B1(_04808_),
    .Y(_05070_));
 sky130_fd_sc_hd__o32ai_4 _15669_ (.A1(_04558_),
    .A2(_04353_),
    .A3(_04554_),
    .B1(_04375_),
    .B2(_04080_),
    .Y(_05071_));
 sky130_fd_sc_hd__o31ai_4 _15670_ (.A1(net262),
    .A2(net245),
    .A3(_04787_),
    .B1(net13),
    .Y(_05072_));
 sky130_fd_sc_hd__nand4b_4 _15671_ (.A_N(_11409_),
    .B(_04113_),
    .C(net309),
    .D(net282),
    .Y(_05073_));
 sky130_fd_sc_hd__nand4_4 _15672_ (.A(_06519_),
    .B(_03955_),
    .C(_04786_),
    .D(_04113_),
    .Y(_05074_));
 sky130_fd_sc_hd__o31a_4 _15673_ (.A1(net11),
    .A2(_04557_),
    .A3(_05073_),
    .B1(_05072_),
    .X(_05076_));
 sky130_fd_sc_hd__o21ai_4 _15674_ (.A1(_04787_),
    .A2(net208),
    .B1(net210),
    .Y(_05077_));
 sky130_fd_sc_hd__o211ai_2 _15675_ (.A1(_04787_),
    .A2(_05073_),
    .B1(net33),
    .C1(_05072_),
    .Y(_05078_));
 sky130_fd_sc_hd__nand3_1 _15676_ (.A(_04790_),
    .B(_04484_),
    .C(net185),
    .Y(_05079_));
 sky130_fd_sc_hd__nor2_2 _15677_ (.A(_04091_),
    .B(_04331_),
    .Y(_05080_));
 sky130_fd_sc_hd__or3_2 _15678_ (.A(net44),
    .B(_04091_),
    .C(_03286_),
    .X(_05081_));
 sky130_fd_sc_hd__nand4_2 _15679_ (.A(_05072_),
    .B(net183),
    .C(_05080_),
    .D(net33),
    .Y(_05082_));
 sky130_fd_sc_hd__nand3_4 _15680_ (.A(_05078_),
    .B(_05079_),
    .C(_05081_),
    .Y(_05083_));
 sky130_fd_sc_hd__a21oi_2 _15681_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_05071_),
    .Y(_05084_));
 sky130_fd_sc_hd__a21o_1 _15682_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_05071_),
    .X(_05085_));
 sky130_fd_sc_hd__o311a_2 _15683_ (.A1(_03286_),
    .A2(_05077_),
    .A3(_05081_),
    .B1(_05083_),
    .C1(_05071_),
    .X(_05087_));
 sky130_fd_sc_hd__nand3_1 _15684_ (.A(_05071_),
    .B(_05082_),
    .C(_05083_),
    .Y(_05088_));
 sky130_fd_sc_hd__a32oi_4 _15685_ (.A1(_04794_),
    .A2(_04795_),
    .A3(_04797_),
    .B1(_04799_),
    .B2(_04784_),
    .Y(_05089_));
 sky130_fd_sc_hd__a32o_2 _15686_ (.A1(_04794_),
    .A2(_04795_),
    .A3(_04797_),
    .B1(_04784_),
    .B2(_04799_),
    .X(_05090_));
 sky130_fd_sc_hd__a21oi_1 _15687_ (.A1(_05085_),
    .A2(_05088_),
    .B1(_05089_),
    .Y(_05091_));
 sky130_fd_sc_hd__o21ai_4 _15688_ (.A1(_05084_),
    .A2(_05087_),
    .B1(_05090_),
    .Y(_05092_));
 sky130_fd_sc_hd__and3_1 _15689_ (.A(_05085_),
    .B(_05088_),
    .C(_05089_),
    .X(_05093_));
 sky130_fd_sc_hd__nand3_2 _15690_ (.A(_05085_),
    .B(_05088_),
    .C(_05089_),
    .Y(_05094_));
 sky130_fd_sc_hd__o32a_2 _15691_ (.A1(_05238_),
    .A2(net247),
    .A3(_03957_),
    .B1(_05260_),
    .B2(_04048_),
    .X(_05095_));
 sky130_fd_sc_hd__a32o_2 _15692_ (.A1(_03952_),
    .A2(net232),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net7),
    .X(_05096_));
 sky130_fd_sc_hd__nand3_2 _15693_ (.A(net226),
    .B(net317),
    .C(_04409_),
    .Y(_05098_));
 sky130_fd_sc_hd__or3b_2 _15694_ (.A(net58),
    .B(_04069_),
    .C_N(net55),
    .X(_05099_));
 sky130_fd_sc_hd__and3b_1 _15695_ (.A_N(net59),
    .B(net8),
    .C(net58),
    .X(_05100_));
 sky130_fd_sc_hd__or3b_2 _15696_ (.A(net59),
    .B(_04059_),
    .C_N(net58),
    .X(_05101_));
 sky130_fd_sc_hd__nand3_1 _15697_ (.A(_04132_),
    .B(_04889_),
    .C(_04130_),
    .Y(_05102_));
 sky130_fd_sc_hd__a31oi_1 _15698_ (.A1(_04132_),
    .A2(_04889_),
    .A3(_04130_),
    .B1(_05100_),
    .Y(_05103_));
 sky130_fd_sc_hd__nand4_4 _15699_ (.A(_05098_),
    .B(_05099_),
    .C(_05101_),
    .D(_05102_),
    .Y(_05104_));
 sky130_fd_sc_hd__a221o_1 _15700_ (.A1(net7),
    .A2(_05249_),
    .B1(_03959_),
    .B2(_05227_),
    .C1(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__a21oi_2 _15701_ (.A1(_05098_),
    .A2(_05099_),
    .B1(_05103_),
    .Y(_05106_));
 sky130_fd_sc_hd__a22o_2 _15702_ (.A1(_05098_),
    .A2(_05099_),
    .B1(_05101_),
    .B2(_05102_),
    .X(_05107_));
 sky130_fd_sc_hd__a21o_2 _15703_ (.A1(_05096_),
    .A2(_05104_),
    .B1(_05106_),
    .X(_05109_));
 sky130_fd_sc_hd__a21oi_4 _15704_ (.A1(_05096_),
    .A2(_05104_),
    .B1(_05106_),
    .Y(_05110_));
 sky130_fd_sc_hd__o21ai_2 _15705_ (.A1(_05096_),
    .A2(_05104_),
    .B1(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__and3_1 _15706_ (.A(_05107_),
    .B(_05095_),
    .C(_05104_),
    .X(_05112_));
 sky130_fd_sc_hd__a21oi_2 _15707_ (.A1(_05104_),
    .A2(_05107_),
    .B1(_05095_),
    .Y(_05113_));
 sky130_fd_sc_hd__and3_1 _15708_ (.A(_05096_),
    .B(_05104_),
    .C(_05107_),
    .X(_05114_));
 sky130_fd_sc_hd__a21oi_1 _15709_ (.A1(_05104_),
    .A2(_05107_),
    .B1(_05096_),
    .Y(_05115_));
 sky130_fd_sc_hd__a22oi_2 _15710_ (.A1(_05106_),
    .A2(_05096_),
    .B1(_05105_),
    .B2(_05110_),
    .Y(_05116_));
 sky130_fd_sc_hd__o21ai_1 _15711_ (.A1(_05095_),
    .A2(_05107_),
    .B1(_05111_),
    .Y(_05117_));
 sky130_fd_sc_hd__o2bb2ai_4 _15712_ (.A1_N(_05092_),
    .A2_N(_05094_),
    .B1(_05112_),
    .B2(_05113_),
    .Y(_05118_));
 sky130_fd_sc_hd__o2111ai_4 _15713_ (.A1(_05095_),
    .A2(_05107_),
    .B1(_05111_),
    .C1(_05094_),
    .D1(_05092_),
    .Y(_05120_));
 sky130_fd_sc_hd__o2bb2ai_1 _15714_ (.A1_N(_05092_),
    .A2_N(_05094_),
    .B1(_05114_),
    .B2(_05115_),
    .Y(_05121_));
 sky130_fd_sc_hd__o21ai_1 _15715_ (.A1(_05112_),
    .A2(_05113_),
    .B1(_05092_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand3_4 _15716_ (.A(_05118_),
    .B(_05120_),
    .C(_05070_),
    .Y(_05123_));
 sky130_fd_sc_hd__a22oi_4 _15717_ (.A1(_04809_),
    .A2(_04811_),
    .B1(_05118_),
    .B2(_05120_),
    .Y(_05124_));
 sky130_fd_sc_hd__o221ai_4 _15718_ (.A1(_05093_),
    .A2(_05122_),
    .B1(_04808_),
    .B2(_04810_),
    .C1(_05121_),
    .Y(_05125_));
 sky130_fd_sc_hd__a21oi_2 _15719_ (.A1(_04825_),
    .A2(_04832_),
    .B1(_04829_),
    .Y(_05126_));
 sky130_fd_sc_hd__inv_2 _15720_ (.A(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__a32o_1 _15721_ (.A1(net235),
    .A2(_12999_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net4),
    .X(_05128_));
 sky130_fd_sc_hd__o211ai_4 _15722_ (.A1(net254),
    .A2(_00646_),
    .B1(net292),
    .C1(_00625_),
    .Y(_05129_));
 sky130_fd_sc_hd__or3b_2 _15723_ (.A(net62),
    .B(_04015_),
    .C_N(net61),
    .X(_05131_));
 sky130_fd_sc_hd__o211ai_4 _15724_ (.A1(net254),
    .A2(_02442_),
    .B1(net299),
    .C1(_02421_),
    .Y(_05132_));
 sky130_fd_sc_hd__or3b_1 _15725_ (.A(net61),
    .B(_04026_),
    .C_N(net60),
    .X(_05133_));
 sky130_fd_sc_hd__a22oi_2 _15726_ (.A1(_05129_),
    .A2(_05131_),
    .B1(_05132_),
    .B2(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__a22o_1 _15727_ (.A1(_05129_),
    .A2(_05131_),
    .B1(_05132_),
    .B2(_05133_),
    .X(_05135_));
 sky130_fd_sc_hd__o2111a_1 _15728_ (.A1(_04026_),
    .A2(net298),
    .B1(_05129_),
    .C1(_05131_),
    .D1(_05132_),
    .X(_05136_));
 sky130_fd_sc_hd__o2111ai_4 _15729_ (.A1(_04026_),
    .A2(net298),
    .B1(_05129_),
    .C1(_05131_),
    .D1(_05132_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand3_4 _15730_ (.A(_05128_),
    .B(_05135_),
    .C(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__o21bai_4 _15731_ (.A1(_05134_),
    .A2(_05136_),
    .B1_N(_05128_),
    .Y(_05139_));
 sky130_fd_sc_hd__a2bb2oi_2 _15732_ (.A1_N(_04765_),
    .A2_N(_04772_),
    .B1(_05138_),
    .B2(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__a21o_1 _15733_ (.A1(_05138_),
    .A2(_05139_),
    .B1(_04774_),
    .X(_05142_));
 sky130_fd_sc_hd__o211a_1 _15734_ (.A1(_04770_),
    .A2(_04773_),
    .B1(_05138_),
    .C1(_05139_),
    .X(_05143_));
 sky130_fd_sc_hd__o211ai_4 _15735_ (.A1(_04770_),
    .A2(_04773_),
    .B1(_05138_),
    .C1(_05139_),
    .Y(_05144_));
 sky130_fd_sc_hd__o221a_1 _15736_ (.A1(_04823_),
    .A2(_04831_),
    .B1(_05140_),
    .B2(_05143_),
    .C1(_04830_),
    .X(_05145_));
 sky130_fd_sc_hd__and3_1 _15737_ (.A(_05127_),
    .B(_05142_),
    .C(_05144_),
    .X(_05146_));
 sky130_fd_sc_hd__and3_1 _15738_ (.A(_05142_),
    .B(_05144_),
    .C(_05126_),
    .X(_05147_));
 sky130_fd_sc_hd__o2111ai_4 _15739_ (.A1(_04823_),
    .A2(_04831_),
    .B1(_05142_),
    .C1(_05144_),
    .D1(_04830_),
    .Y(_05148_));
 sky130_fd_sc_hd__o22a_1 _15740_ (.A1(_04829_),
    .A2(_04836_),
    .B1(_05140_),
    .B2(_05143_),
    .X(_05149_));
 sky130_fd_sc_hd__o21ai_2 _15741_ (.A1(_05140_),
    .A2(_05143_),
    .B1(_05127_),
    .Y(_05150_));
 sky130_fd_sc_hd__nand2_1 _15742_ (.A(_05148_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__a32oi_4 _15743_ (.A1(_05118_),
    .A2(_05120_),
    .A3(_05070_),
    .B1(_05148_),
    .B2(_05150_),
    .Y(_05153_));
 sky130_fd_sc_hd__o21ai_1 _15744_ (.A1(_05147_),
    .A2(_05149_),
    .B1(_05123_),
    .Y(_05154_));
 sky130_fd_sc_hd__o2bb2ai_1 _15745_ (.A1_N(_05123_),
    .A2_N(_05125_),
    .B1(_05145_),
    .B2(_05146_),
    .Y(_05155_));
 sky130_fd_sc_hd__o211ai_4 _15746_ (.A1(_05145_),
    .A2(_05146_),
    .B1(_05123_),
    .C1(_05125_),
    .Y(_05156_));
 sky130_fd_sc_hd__o2bb2ai_2 _15747_ (.A1_N(_05123_),
    .A2_N(_05125_),
    .B1(_05147_),
    .B2(_05149_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand3_2 _15748_ (.A(_05069_),
    .B(_05156_),
    .C(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__o211ai_4 _15749_ (.A1(_05124_),
    .A2(_05154_),
    .B1(_05068_),
    .C1(_05155_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand4_2 _15750_ (.A(_05063_),
    .B(_05066_),
    .C(_05158_),
    .D(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__a22o_1 _15751_ (.A1(_05063_),
    .A2(_05066_),
    .B1(_05158_),
    .B2(_05159_),
    .X(_05161_));
 sky130_fd_sc_hd__nand3_2 _15752_ (.A(_05067_),
    .B(_05158_),
    .C(_05159_),
    .Y(_05162_));
 sky130_fd_sc_hd__a21o_1 _15753_ (.A1(_05158_),
    .A2(_05159_),
    .B1(_05067_),
    .X(_05164_));
 sky130_fd_sc_hd__a32o_1 _15754_ (.A1(_04757_),
    .A2(_04847_),
    .A3(_04848_),
    .B1(_04855_),
    .B2(_04755_),
    .X(_05165_));
 sky130_fd_sc_hd__o211a_1 _15755_ (.A1(_04854_),
    .A2(_04860_),
    .B1(_05160_),
    .C1(_05161_),
    .X(_05166_));
 sky130_fd_sc_hd__o211ai_4 _15756_ (.A1(_04854_),
    .A2(_04860_),
    .B1(_05160_),
    .C1(_05161_),
    .Y(_05167_));
 sky130_fd_sc_hd__o2111ai_4 _15757_ (.A1(_04755_),
    .A2(_04852_),
    .B1(_04855_),
    .C1(_05162_),
    .D1(_05164_),
    .Y(_05168_));
 sky130_fd_sc_hd__a21o_1 _15758_ (.A1(_05167_),
    .A2(_05168_),
    .B1(_05016_),
    .X(_05169_));
 sky130_fd_sc_hd__o211ai_4 _15759_ (.A1(_05011_),
    .A2(_05013_),
    .B1(_05167_),
    .C1(_05168_),
    .Y(_05170_));
 sky130_fd_sc_hd__a22o_1 _15760_ (.A1(_05012_),
    .A2(_05014_),
    .B1(_05167_),
    .B2(_05168_),
    .X(_05171_));
 sky130_fd_sc_hd__nand4_1 _15761_ (.A(_05012_),
    .B(_05014_),
    .C(_05167_),
    .D(_05168_),
    .Y(_05172_));
 sky130_fd_sc_hd__a21oi_2 _15762_ (.A1(_05169_),
    .A2(_05170_),
    .B1(_04949_),
    .Y(_05173_));
 sky130_fd_sc_hd__a22o_1 _15763_ (.A1(_04863_),
    .A2(_04917_),
    .B1(_05169_),
    .B2(_05170_),
    .X(_05175_));
 sky130_fd_sc_hd__and3_1 _15764_ (.A(_05169_),
    .B(_05170_),
    .C(_04949_),
    .X(_05176_));
 sky130_fd_sc_hd__o21ai_1 _15765_ (.A1(_05173_),
    .A2(_05176_),
    .B1(_04947_),
    .Y(_05177_));
 sky130_fd_sc_hd__nand3b_1 _15766_ (.A_N(_05176_),
    .B(_04948_),
    .C(_05175_),
    .Y(_05178_));
 sky130_fd_sc_hd__a211o_1 _15767_ (.A1(_05171_),
    .A2(_05172_),
    .B1(_04948_),
    .C1(_04950_),
    .X(_05179_));
 sky130_fd_sc_hd__a31oi_2 _15768_ (.A1(_04950_),
    .A2(_05171_),
    .A3(_05172_),
    .B1(_04948_),
    .Y(_05180_));
 sky130_fd_sc_hd__a31oi_2 _15769_ (.A1(_05169_),
    .A2(_05170_),
    .A3(_04949_),
    .B1(_04947_),
    .Y(_05181_));
 sky130_fd_sc_hd__o21ai_1 _15770_ (.A1(_05176_),
    .A2(_05180_),
    .B1(_05179_),
    .Y(_05182_));
 sky130_fd_sc_hd__nand3_2 _15771_ (.A(_04946_),
    .B(_05177_),
    .C(_05178_),
    .Y(_05183_));
 sky130_fd_sc_hd__o211ai_2 _15772_ (.A1(_04947_),
    .A2(_05175_),
    .B1(_04945_),
    .C1(_05182_),
    .Y(_05184_));
 sky130_fd_sc_hd__nand2_1 _15773_ (.A(_05183_),
    .B(_05184_),
    .Y(_05186_));
 sky130_fd_sc_hd__a221oi_2 _15774_ (.A1(_04691_),
    .A2(_04928_),
    .B1(_05183_),
    .B2(_05184_),
    .C1(_04929_),
    .Y(_05187_));
 sky130_fd_sc_hd__a21oi_1 _15775_ (.A1(_04930_),
    .A2(_04932_),
    .B1(_05186_),
    .Y(_05188_));
 sky130_fd_sc_hd__or2_1 _15776_ (.A(_04930_),
    .B(_05186_),
    .X(_05189_));
 sky130_fd_sc_hd__nor2_1 _15777_ (.A(_05187_),
    .B(_05188_),
    .Y(_05190_));
 sky130_fd_sc_hd__xor2_1 _15778_ (.A(_04944_),
    .B(_05190_),
    .X(net77));
 sky130_fd_sc_hd__a2bb2o_1 _15779_ (.A1_N(_04932_),
    .A2_N(_05186_),
    .B1(_05190_),
    .B2(_04944_),
    .X(_05191_));
 sky130_fd_sc_hd__a31o_1 _15780_ (.A1(_04975_),
    .A2(_04977_),
    .A3(_04981_),
    .B1(_05003_),
    .X(_05192_));
 sky130_fd_sc_hd__a21o_1 _15781_ (.A1(_04953_),
    .A2(_04962_),
    .B1(_04961_),
    .X(_05193_));
 sky130_fd_sc_hd__a21oi_1 _15782_ (.A1(_05017_),
    .A2(_05025_),
    .B1(_05023_),
    .Y(_05194_));
 sky130_fd_sc_hd__a21o_1 _15783_ (.A1(_05017_),
    .A2(_05025_),
    .B1(_05023_),
    .X(_05196_));
 sky130_fd_sc_hd__a32oi_4 _15784_ (.A1(net266),
    .A2(net303),
    .A3(net280),
    .B1(_04269_),
    .B2(net27),
    .Y(_05197_));
 sky130_fd_sc_hd__o211ai_1 _15785_ (.A1(_04747_),
    .A2(_05436_),
    .B1(_04215_),
    .C1(_05414_),
    .Y(_05198_));
 sky130_fd_sc_hd__a32oi_4 _15786_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_04215_),
    .B1(_04217_),
    .B2(net28),
    .Y(_05199_));
 sky130_fd_sc_hd__or3_2 _15787_ (.A(net39),
    .B(_04037_),
    .C(_03835_),
    .X(_05200_));
 sky130_fd_sc_hd__nand4_2 _15788_ (.A(_04037_),
    .B(_05841_),
    .C(net265),
    .D(net39),
    .Y(_05201_));
 sky130_fd_sc_hd__o31a_1 _15789_ (.A1(_03835_),
    .A2(_04037_),
    .A3(net39),
    .B1(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__o2111a_1 _15790_ (.A1(_03725_),
    .A2(_04218_),
    .B1(_05198_),
    .C1(_05200_),
    .D1(_05201_),
    .X(_05203_));
 sky130_fd_sc_hd__a21oi_1 _15791_ (.A1(_05200_),
    .A2(_05201_),
    .B1(_05199_),
    .Y(_05204_));
 sky130_fd_sc_hd__o21bai_1 _15792_ (.A1(_05199_),
    .A2(_05202_),
    .B1_N(_05197_),
    .Y(_05205_));
 sky130_fd_sc_hd__o21ai_1 _15793_ (.A1(_05203_),
    .A2(_05204_),
    .B1(_05197_),
    .Y(_05206_));
 sky130_fd_sc_hd__a211o_1 _15794_ (.A1(_05200_),
    .A2(_05201_),
    .B1(_05197_),
    .C1(_05199_),
    .X(_05207_));
 sky130_fd_sc_hd__nand4_1 _15795_ (.A(_05197_),
    .B(_05199_),
    .C(_05200_),
    .D(_05201_),
    .Y(_05208_));
 sky130_fd_sc_hd__a31o_1 _15796_ (.A1(_05199_),
    .A2(_05200_),
    .A3(_05201_),
    .B1(_05197_),
    .X(_05209_));
 sky130_fd_sc_hd__o21ai_1 _15797_ (.A1(_05199_),
    .A2(_05202_),
    .B1(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__o21a_1 _15798_ (.A1(_05199_),
    .A2(_05202_),
    .B1(_05209_),
    .X(_05211_));
 sky130_fd_sc_hd__o211ai_1 _15799_ (.A1(_05199_),
    .A2(_05202_),
    .B1(_05208_),
    .C1(_05209_),
    .Y(_05212_));
 sky130_fd_sc_hd__o211a_1 _15800_ (.A1(_05203_),
    .A2(_05205_),
    .B1(_05206_),
    .C1(_05196_),
    .X(_05213_));
 sky130_fd_sc_hd__o211ai_2 _15801_ (.A1(_05203_),
    .A2(_05205_),
    .B1(_05206_),
    .C1(_05196_),
    .Y(_05214_));
 sky130_fd_sc_hd__nand3_2 _15802_ (.A(_05212_),
    .B(_05194_),
    .C(_05207_),
    .Y(_05215_));
 sky130_fd_sc_hd__a21oi_1 _15803_ (.A1(_05214_),
    .A2(_05215_),
    .B1(_05193_),
    .Y(_05217_));
 sky130_fd_sc_hd__a221o_1 _15804_ (.A1(_04957_),
    .A2(_04959_),
    .B1(_05214_),
    .B2(_05215_),
    .C1(_04967_),
    .X(_05218_));
 sky130_fd_sc_hd__and3_1 _15805_ (.A(_05193_),
    .B(_05214_),
    .C(_05215_),
    .X(_05219_));
 sky130_fd_sc_hd__o211ai_1 _15806_ (.A1(_04961_),
    .A2(_04967_),
    .B1(_05214_),
    .C1(_05215_),
    .Y(_05220_));
 sky130_fd_sc_hd__o21ai_1 _15807_ (.A1(_04952_),
    .A2(_04973_),
    .B1(_04972_),
    .Y(_05221_));
 sky130_fd_sc_hd__o221ai_4 _15808_ (.A1(_04952_),
    .A2(_04973_),
    .B1(_05217_),
    .B2(_05219_),
    .C1(_04972_),
    .Y(_05222_));
 sky130_fd_sc_hd__and3_2 _15809_ (.A(_05218_),
    .B(_05220_),
    .C(_05221_),
    .X(_05223_));
 sky130_fd_sc_hd__nand3_2 _15810_ (.A(_05218_),
    .B(_05220_),
    .C(_05221_),
    .Y(_05224_));
 sky130_fd_sc_hd__and2b_4 _15811_ (.A_N(net45),
    .B(net46),
    .X(_05225_));
 sky130_fd_sc_hd__nand2_8 _15812_ (.A(_04124_),
    .B(net46),
    .Y(_05226_));
 sky130_fd_sc_hd__nor2_8 _15813_ (.A(net46),
    .B(_04124_),
    .Y(_05228_));
 sky130_fd_sc_hd__or2_4 _15814_ (.A(net46),
    .B(_04124_),
    .X(_05229_));
 sky130_fd_sc_hd__o21ai_1 _15815_ (.A1(net276),
    .A2(_05228_),
    .B1(net1),
    .Y(_05230_));
 sky130_fd_sc_hd__a21o_1 _15816_ (.A1(_04997_),
    .A2(_04990_),
    .B1(_04995_),
    .X(_05231_));
 sky130_fd_sc_hd__a22o_1 _15817_ (.A1(net12),
    .A2(_04988_),
    .B1(_04539_),
    .B2(_04985_),
    .X(_05232_));
 sky130_fd_sc_hd__o32a_1 _15818_ (.A1(_04896_),
    .A2(_04441_),
    .A3(_04408_),
    .B1(_03396_),
    .B2(_04898_),
    .X(_05233_));
 sky130_fd_sc_hd__a32o_1 _15819_ (.A1(net243),
    .A2(_04452_),
    .A3(net318),
    .B1(net23),
    .B2(_04897_),
    .X(_05234_));
 sky130_fd_sc_hd__a32o_1 _15820_ (.A1(net315),
    .A2(net267),
    .A3(net279),
    .B1(_04482_),
    .B2(net26),
    .X(_05235_));
 sky130_fd_sc_hd__nand2_1 _15821_ (.A(_05234_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__o221ai_4 _15822_ (.A1(_04758_),
    .A2(_04481_),
    .B1(_04483_),
    .B2(_03506_),
    .C1(_05233_),
    .Y(_05237_));
 sky130_fd_sc_hd__nand3_1 _15823_ (.A(_05232_),
    .B(_05236_),
    .C(_05237_),
    .Y(_05239_));
 sky130_fd_sc_hd__a21o_1 _15824_ (.A1(_05236_),
    .A2(_05237_),
    .B1(_05232_),
    .X(_05240_));
 sky130_fd_sc_hd__o211ai_2 _15825_ (.A1(_04995_),
    .A2(_05000_),
    .B1(_05239_),
    .C1(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__a21o_1 _15826_ (.A1(_05239_),
    .A2(_05240_),
    .B1(_05231_),
    .X(_05242_));
 sky130_fd_sc_hd__nand2_1 _15827_ (.A(_05241_),
    .B(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__o2111a_1 _15828_ (.A1(net276),
    .A2(_05228_),
    .B1(net1),
    .C1(_05241_),
    .D1(_05242_),
    .X(_05244_));
 sky130_fd_sc_hd__and2_1 _15829_ (.A(_05230_),
    .B(_05243_),
    .X(_05245_));
 sky130_fd_sc_hd__and3_1 _15830_ (.A(_05230_),
    .B(_05241_),
    .C(_05242_),
    .X(_05246_));
 sky130_fd_sc_hd__o211a_1 _15831_ (.A1(net276),
    .A2(_05228_),
    .B1(net1),
    .C1(_05243_),
    .X(_05247_));
 sky130_fd_sc_hd__o2bb2ai_2 _15832_ (.A1_N(_05222_),
    .A2_N(_05224_),
    .B1(_05244_),
    .B2(_05245_),
    .Y(_05248_));
 sky130_fd_sc_hd__o21ai_4 _15833_ (.A1(_05246_),
    .A2(_05247_),
    .B1(_05222_),
    .Y(_05250_));
 sky130_fd_sc_hd__o21ai_2 _15834_ (.A1(_05223_),
    .A2(_05250_),
    .B1(_05248_),
    .Y(_05251_));
 sky130_fd_sc_hd__nor2_1 _15835_ (.A(_05061_),
    .B(_05065_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_2 _15836_ (.A(_05251_),
    .B(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__o221ai_4 _15837_ (.A1(_05223_),
    .A2(_05250_),
    .B1(_05061_),
    .B2(_05065_),
    .C1(_05248_),
    .Y(_05254_));
 sky130_fd_sc_hd__a22oi_4 _15838_ (.A1(_04982_),
    .A2(_05192_),
    .B1(_05253_),
    .B2(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__o22a_1 _15839_ (.A1(_04983_),
    .A2(_05005_),
    .B1(_05252_),
    .B2(_05251_),
    .X(_05256_));
 sky130_fd_sc_hd__o211a_1 _15840_ (.A1(_04983_),
    .A2(_05005_),
    .B1(_05253_),
    .C1(_05254_),
    .X(_05257_));
 sky130_fd_sc_hd__nand2_1 _15841_ (.A(_05256_),
    .B(_05253_),
    .Y(_05258_));
 sky130_fd_sc_hd__a21oi_1 _15842_ (.A1(_05253_),
    .A2(_05256_),
    .B1(_05255_),
    .Y(_05259_));
 sky130_fd_sc_hd__a21o_1 _15843_ (.A1(_05253_),
    .A2(_05256_),
    .B1(_05255_),
    .X(_05261_));
 sky130_fd_sc_hd__a32oi_4 _15844_ (.A1(_05069_),
    .A2(_05156_),
    .A3(_05157_),
    .B1(_05159_),
    .B2(_05067_),
    .Y(_05262_));
 sky130_fd_sc_hd__a21oi_1 _15845_ (.A1(_05123_),
    .A2(_05151_),
    .B1(_05124_),
    .Y(_05263_));
 sky130_fd_sc_hd__a21oi_1 _15846_ (.A1(_05092_),
    .A2(_05117_),
    .B1(_05093_),
    .Y(_05264_));
 sky130_fd_sc_hd__o32ai_4 _15847_ (.A1(_05084_),
    .A2(_05090_),
    .A3(_05087_),
    .B1(_05116_),
    .B2(_05091_),
    .Y(_05265_));
 sky130_fd_sc_hd__o22a_1 _15848_ (.A1(_04059_),
    .A2(_05260_),
    .B1(_04133_),
    .B2(_05238_),
    .X(_05266_));
 sky130_fd_sc_hd__a32o_1 _15849_ (.A1(_04132_),
    .A2(_05227_),
    .A3(net230),
    .B1(_05249_),
    .B2(net8),
    .X(_05267_));
 sky130_fd_sc_hd__and3b_1 _15850_ (.A_N(net59),
    .B(net9),
    .C(net58),
    .X(_05268_));
 sky130_fd_sc_hd__a31oi_4 _15851_ (.A1(net224),
    .A2(net305),
    .A3(net188),
    .B1(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__o211ai_2 _15852_ (.A1(net232),
    .A2(_04557_),
    .B1(net317),
    .C1(_04555_),
    .Y(_05270_));
 sky130_fd_sc_hd__or3b_1 _15853_ (.A(net58),
    .B(_04080_),
    .C_N(net55),
    .X(_05272_));
 sky130_fd_sc_hd__a32oi_2 _15854_ (.A1(_04555_),
    .A2(_04559_),
    .A3(net317),
    .B1(_04649_),
    .B2(net10),
    .Y(_05273_));
 sky130_fd_sc_hd__a21oi_2 _15855_ (.A1(_05270_),
    .A2(_05272_),
    .B1(_05269_),
    .Y(_05274_));
 sky130_fd_sc_hd__a21o_1 _15856_ (.A1(_05270_),
    .A2(_05272_),
    .B1(_05269_),
    .X(_05275_));
 sky130_fd_sc_hd__o211a_1 _15857_ (.A1(_04080_),
    .A2(net316),
    .B1(_05270_),
    .C1(_05269_),
    .X(_05276_));
 sky130_fd_sc_hd__o221ai_4 _15858_ (.A1(_04080_),
    .A2(net316),
    .B1(_04562_),
    .B2(_04638_),
    .C1(_05269_),
    .Y(_05277_));
 sky130_fd_sc_hd__a21oi_1 _15859_ (.A1(_05275_),
    .A2(_05277_),
    .B1(_05266_),
    .Y(_05278_));
 sky130_fd_sc_hd__o21ai_4 _15860_ (.A1(_05274_),
    .A2(_05276_),
    .B1(_05267_),
    .Y(_05279_));
 sky130_fd_sc_hd__nor3_1 _15861_ (.A(_05267_),
    .B(_05274_),
    .C(_05276_),
    .Y(_05280_));
 sky130_fd_sc_hd__nand3_2 _15862_ (.A(_05275_),
    .B(_05277_),
    .C(_05266_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(_05279_),
    .B(_05281_),
    .Y(_05283_));
 sky130_fd_sc_hd__a32oi_4 _15864_ (.A1(net33),
    .A2(_05076_),
    .A3(_05080_),
    .B1(_05083_),
    .B2(_05071_),
    .Y(_05284_));
 sky130_fd_sc_hd__a32o_1 _15865_ (.A1(net33),
    .A2(_05076_),
    .A3(_05080_),
    .B1(_05083_),
    .B2(_05071_),
    .X(_05285_));
 sky130_fd_sc_hd__nor2_1 _15866_ (.A(_04091_),
    .B(_04375_),
    .Y(_05286_));
 sky130_fd_sc_hd__o311a_1 _15867_ (.A1(net7),
    .A2(net249),
    .A3(_04787_),
    .B1(_04342_),
    .C1(_04790_),
    .X(_05287_));
 sky130_fd_sc_hd__a21oi_1 _15868_ (.A1(_04342_),
    .A2(_04792_),
    .B1(_05286_),
    .Y(_05288_));
 sky130_fd_sc_hd__a31o_1 _15869_ (.A1(_04790_),
    .A2(_04342_),
    .A3(net185),
    .B1(_05286_),
    .X(_05289_));
 sky130_fd_sc_hd__o21bai_4 _15870_ (.A1(_04787_),
    .A2(net208),
    .B1_N(_04135_),
    .Y(_05290_));
 sky130_fd_sc_hd__nor2_4 _15871_ (.A(net13),
    .B(net14),
    .Y(_05291_));
 sky130_fd_sc_hd__nand4_4 _15872_ (.A(_06519_),
    .B(_03955_),
    .C(net277),
    .D(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nand2_8 _15873_ (.A(net181),
    .B(net180),
    .Y(_05294_));
 sky130_fd_sc_hd__nand3_2 _15874_ (.A(net181),
    .B(net180),
    .C(net33),
    .Y(_05295_));
 sky130_fd_sc_hd__o211ai_1 _15875_ (.A1(_04787_),
    .A2(_05073_),
    .B1(_04484_),
    .C1(_05072_),
    .Y(_05296_));
 sky130_fd_sc_hd__nor2_1 _15876_ (.A(_04113_),
    .B(_04331_),
    .Y(_05297_));
 sky130_fd_sc_hd__or3_1 _15877_ (.A(net44),
    .B(_04113_),
    .C(_03286_),
    .X(_05298_));
 sky130_fd_sc_hd__a31oi_2 _15878_ (.A1(_05072_),
    .A2(net183),
    .A3(_04484_),
    .B1(_05297_),
    .Y(_05299_));
 sky130_fd_sc_hd__nand3_2 _15879_ (.A(_05295_),
    .B(_05296_),
    .C(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__and3_2 _15880_ (.A(net13),
    .B(_04320_),
    .C(_04135_),
    .X(_05301_));
 sky130_fd_sc_hd__or4_1 _15881_ (.A(net44),
    .B(net14),
    .C(_04113_),
    .D(_03286_),
    .X(_05302_));
 sky130_fd_sc_hd__a211o_1 _15882_ (.A1(_05299_),
    .A2(_05295_),
    .B1(_05301_),
    .C1(_05289_),
    .X(_05303_));
 sky130_fd_sc_hd__a21o_1 _15883_ (.A1(_05300_),
    .A2(_05302_),
    .B1(_05288_),
    .X(_05305_));
 sky130_fd_sc_hd__a21o_1 _15884_ (.A1(_05300_),
    .A2(_05302_),
    .B1(_05289_),
    .X(_05306_));
 sky130_fd_sc_hd__o2bb2ai_2 _15885_ (.A1_N(_05295_),
    .A2_N(_05299_),
    .B1(_05286_),
    .B2(_05287_),
    .Y(_05307_));
 sky130_fd_sc_hd__nand3_2 _15886_ (.A(_05305_),
    .B(_05284_),
    .C(_05303_),
    .Y(_05308_));
 sky130_fd_sc_hd__o211a_2 _15887_ (.A1(_05307_),
    .A2(_05301_),
    .B1(_05285_),
    .C1(_05306_),
    .X(_05309_));
 sky130_fd_sc_hd__o211ai_4 _15888_ (.A1(_05307_),
    .A2(_05301_),
    .B1(_05285_),
    .C1(_05306_),
    .Y(_05310_));
 sky130_fd_sc_hd__nand4_2 _15889_ (.A(_05279_),
    .B(_05281_),
    .C(_05308_),
    .D(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__a22o_1 _15890_ (.A1(_05279_),
    .A2(_05281_),
    .B1(_05308_),
    .B2(_05310_),
    .X(_05312_));
 sky130_fd_sc_hd__a32oi_4 _15891_ (.A1(_05305_),
    .A2(_05284_),
    .A3(_05303_),
    .B1(_05281_),
    .B2(_05279_),
    .Y(_05313_));
 sky130_fd_sc_hd__o21ai_2 _15892_ (.A1(_05278_),
    .A2(_05280_),
    .B1(_05308_),
    .Y(_05314_));
 sky130_fd_sc_hd__and3_1 _15893_ (.A(_05283_),
    .B(_05308_),
    .C(_05310_),
    .X(_05316_));
 sky130_fd_sc_hd__a21o_1 _15894_ (.A1(_05308_),
    .A2(_05310_),
    .B1(_05283_),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_1 _15895_ (.A(_05265_),
    .B(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__o211ai_4 _15896_ (.A1(_05314_),
    .A2(_05309_),
    .B1(_05265_),
    .C1(_05317_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand3_4 _15897_ (.A(_05312_),
    .B(_05264_),
    .C(_05311_),
    .Y(_05320_));
 sky130_fd_sc_hd__and2_1 _15898_ (.A(_05135_),
    .B(_05138_),
    .X(_05321_));
 sky130_fd_sc_hd__nand2_1 _15899_ (.A(_05135_),
    .B(_05138_),
    .Y(_05322_));
 sky130_fd_sc_hd__and3_1 _15900_ (.A(_03927_),
    .B(net6),
    .C(net61),
    .X(_05323_));
 sky130_fd_sc_hd__a31oi_2 _15901_ (.A1(_02421_),
    .A2(net249),
    .A3(net292),
    .B1(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__a31o_1 _15902_ (.A1(_02421_),
    .A2(net249),
    .A3(net292),
    .B1(_05323_),
    .X(_05325_));
 sky130_fd_sc_hd__o21ai_1 _15903_ (.A1(net263),
    .A2(net246),
    .B1(net299),
    .Y(_05327_));
 sky130_fd_sc_hd__o22ai_2 _15904_ (.A1(_04048_),
    .A2(net298),
    .B1(net247),
    .B2(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__nand2_2 _15905_ (.A(_05325_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__o221ai_4 _15906_ (.A1(_04048_),
    .A2(net298),
    .B1(_03961_),
    .B2(_05699_),
    .C1(_05324_),
    .Y(_05330_));
 sky130_fd_sc_hd__a32o_1 _15907_ (.A1(_00625_),
    .A2(net250),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net5),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_1 _15908_ (.A1(_05329_),
    .A2(_05330_),
    .B1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__a21o_1 _15909_ (.A1(_05329_),
    .A2(_05330_),
    .B1(_05331_),
    .X(_05333_));
 sky130_fd_sc_hd__and3_1 _15910_ (.A(_05329_),
    .B(_05330_),
    .C(_05331_),
    .X(_05334_));
 sky130_fd_sc_hd__nand3_4 _15911_ (.A(_05329_),
    .B(_05330_),
    .C(_05331_),
    .Y(_05335_));
 sky130_fd_sc_hd__nor2_1 _15912_ (.A(_05332_),
    .B(_05334_),
    .Y(_05336_));
 sky130_fd_sc_hd__a21oi_2 _15913_ (.A1(_05333_),
    .A2(_05335_),
    .B1(_05109_),
    .Y(_05338_));
 sky130_fd_sc_hd__o21ai_2 _15914_ (.A1(_05332_),
    .A2(_05334_),
    .B1(_05110_),
    .Y(_05339_));
 sky130_fd_sc_hd__nand3_2 _15915_ (.A(_05333_),
    .B(_05335_),
    .C(_05109_),
    .Y(_05340_));
 sky130_fd_sc_hd__a21oi_2 _15916_ (.A1(_05339_),
    .A2(_05340_),
    .B1(_05322_),
    .Y(_05341_));
 sky130_fd_sc_hd__a21oi_1 _15917_ (.A1(_05135_),
    .A2(_05138_),
    .B1(_05338_),
    .Y(_05342_));
 sky130_fd_sc_hd__and3_1 _15918_ (.A(_05322_),
    .B(_05339_),
    .C(_05340_),
    .X(_05343_));
 sky130_fd_sc_hd__and3_1 _15919_ (.A(_05339_),
    .B(_05340_),
    .C(_05321_),
    .X(_05344_));
 sky130_fd_sc_hd__a21oi_1 _15920_ (.A1(_05339_),
    .A2(_05340_),
    .B1(_05321_),
    .Y(_05345_));
 sky130_fd_sc_hd__a21oi_2 _15921_ (.A1(_05342_),
    .A2(_05340_),
    .B1(_05341_),
    .Y(_05346_));
 sky130_fd_sc_hd__o211ai_4 _15922_ (.A1(_05341_),
    .A2(_05343_),
    .B1(_05319_),
    .C1(_05320_),
    .Y(_05347_));
 sky130_fd_sc_hd__o2bb2ai_2 _15923_ (.A1_N(_05319_),
    .A2_N(_05320_),
    .B1(_05344_),
    .B2(_05345_),
    .Y(_05349_));
 sky130_fd_sc_hd__a21oi_2 _15924_ (.A1(_05319_),
    .A2(_05320_),
    .B1(_05346_),
    .Y(_05350_));
 sky130_fd_sc_hd__o2bb2ai_1 _15925_ (.A1_N(_05319_),
    .A2_N(_05320_),
    .B1(_05341_),
    .B2(_05343_),
    .Y(_05351_));
 sky130_fd_sc_hd__o211ai_2 _15926_ (.A1(_05344_),
    .A2(_05345_),
    .B1(_05319_),
    .C1(_05320_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand3_4 _15927_ (.A(_05349_),
    .B(_05263_),
    .C(_05347_),
    .Y(_05353_));
 sky130_fd_sc_hd__o21ai_2 _15928_ (.A1(_05124_),
    .A2(_05153_),
    .B1(_05352_),
    .Y(_05354_));
 sky130_fd_sc_hd__a2bb2oi_2 _15929_ (.A1_N(_05124_),
    .A2_N(_05153_),
    .B1(_05347_),
    .B2(_05349_),
    .Y(_05355_));
 sky130_fd_sc_hd__o211ai_2 _15930_ (.A1(_05124_),
    .A2(_05153_),
    .B1(_05351_),
    .C1(_05352_),
    .Y(_05356_));
 sky130_fd_sc_hd__o22a_1 _15931_ (.A1(_06552_),
    .A2(_02869_),
    .B1(_02891_),
    .B2(_03916_),
    .X(_05357_));
 sky130_fd_sc_hd__a32o_1 _15932_ (.A1(_06486_),
    .A2(net261),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net30),
    .X(_05358_));
 sky130_fd_sc_hd__nor2_1 _15933_ (.A(_03938_),
    .B(_01326_),
    .Y(_05360_));
 sky130_fd_sc_hd__a31oi_4 _15934_ (.A1(_07242_),
    .A2(net257),
    .A3(_01293_),
    .B1(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__or3_1 _15935_ (.A(net36),
    .B(_03993_),
    .C(_03949_),
    .X(_05362_));
 sky130_fd_sc_hd__o211ai_4 _15936_ (.A1(net261),
    .A2(_08656_),
    .B1(_12330_),
    .C1(_08700_),
    .Y(_05363_));
 sky130_fd_sc_hd__a21oi_2 _15937_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05361_),
    .Y(_05364_));
 sky130_fd_sc_hd__a21o_1 _15938_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05361_),
    .X(_05365_));
 sky130_fd_sc_hd__o211ai_2 _15939_ (.A1(_03949_),
    .A2(_12363_),
    .B1(_05363_),
    .C1(_05361_),
    .Y(_05366_));
 sky130_fd_sc_hd__a21oi_2 _15940_ (.A1(_05365_),
    .A2(_05366_),
    .B1(_05358_),
    .Y(_05367_));
 sky130_fd_sc_hd__and3_1 _15941_ (.A(_05358_),
    .B(_05365_),
    .C(_05366_),
    .X(_05368_));
 sky130_fd_sc_hd__or3b_1 _15942_ (.A(_05357_),
    .B(_05364_),
    .C_N(_05366_),
    .X(_05369_));
 sky130_fd_sc_hd__a22oi_2 _15943_ (.A1(_09709_),
    .A2(net252),
    .B1(_11793_),
    .B2(net2),
    .Y(_05371_));
 sky130_fd_sc_hd__nand3_2 _15944_ (.A(net235),
    .B(net251),
    .C(net291),
    .Y(_05372_));
 sky130_fd_sc_hd__or3b_2 _15945_ (.A(net64),
    .B(_04004_),
    .C_N(net63),
    .X(_05373_));
 sky130_fd_sc_hd__o211ai_4 _15946_ (.A1(net261),
    .A2(_11387_),
    .B1(net289),
    .C1(_11354_),
    .Y(_05374_));
 sky130_fd_sc_hd__or3b_2 _15947_ (.A(net34),
    .B(_03982_),
    .C_N(net64),
    .X(_05375_));
 sky130_fd_sc_hd__a22oi_4 _15948_ (.A1(_05372_),
    .A2(_05373_),
    .B1(_05374_),
    .B2(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__a22o_1 _15949_ (.A1(_05372_),
    .A2(_05373_),
    .B1(_05374_),
    .B2(_05375_),
    .X(_05377_));
 sky130_fd_sc_hd__o2111a_2 _15950_ (.A1(_03982_),
    .A2(_10346_),
    .B1(_05372_),
    .C1(_05373_),
    .D1(_05374_),
    .X(_05378_));
 sky130_fd_sc_hd__o2111ai_1 _15951_ (.A1(_03982_),
    .A2(_10346_),
    .B1(_05372_),
    .C1(_05373_),
    .D1(_05374_),
    .Y(_05379_));
 sky130_fd_sc_hd__o21bai_4 _15952_ (.A1(_05376_),
    .A2(_05378_),
    .B1_N(_05371_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand3_2 _15953_ (.A(_05377_),
    .B(_05379_),
    .C(_05371_),
    .Y(_05382_));
 sky130_fd_sc_hd__a21oi_2 _15954_ (.A1(_05380_),
    .A2(_05382_),
    .B1(_05045_),
    .Y(_05383_));
 sky130_fd_sc_hd__a21o_2 _15955_ (.A1(_05380_),
    .A2(_05382_),
    .B1(_05045_),
    .X(_05384_));
 sky130_fd_sc_hd__and3_1 _15956_ (.A(_05045_),
    .B(_05380_),
    .C(_05382_),
    .X(_05385_));
 sky130_fd_sc_hd__o2111ai_4 _15957_ (.A1(_05032_),
    .A2(_05040_),
    .B1(_05380_),
    .C1(_05382_),
    .D1(_05039_),
    .Y(_05386_));
 sky130_fd_sc_hd__nand4b_4 _15958_ (.A_N(_05367_),
    .B(_05369_),
    .C(_05384_),
    .D(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__o22a_1 _15959_ (.A1(_05367_),
    .A2(_05368_),
    .B1(_05383_),
    .B2(_05385_),
    .X(_05388_));
 sky130_fd_sc_hd__o22ai_4 _15960_ (.A1(_05367_),
    .A2(_05368_),
    .B1(_05383_),
    .B2(_05385_),
    .Y(_05389_));
 sky130_fd_sc_hd__o21ai_4 _15961_ (.A1(_05126_),
    .A2(_05140_),
    .B1(_05144_),
    .Y(_05390_));
 sky130_fd_sc_hd__a21oi_4 _15962_ (.A1(_05387_),
    .A2(_05389_),
    .B1(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _15963_ (.A(_05390_),
    .B(_05387_),
    .Y(_05393_));
 sky130_fd_sc_hd__and3_1 _15964_ (.A(_05390_),
    .B(_05389_),
    .C(_05387_),
    .X(_05394_));
 sky130_fd_sc_hd__nand3_1 _15965_ (.A(_05390_),
    .B(_05389_),
    .C(_05387_),
    .Y(_05395_));
 sky130_fd_sc_hd__o31a_1 _15966_ (.A1(_05027_),
    .A2(_05028_),
    .A3(_05051_),
    .B1(_05050_),
    .X(_05396_));
 sky130_fd_sc_hd__o21bai_1 _15967_ (.A1(_05391_),
    .A2(_05394_),
    .B1_N(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__nand3b_1 _15968_ (.A_N(_05391_),
    .B(_05395_),
    .C(_05396_),
    .Y(_05398_));
 sky130_fd_sc_hd__o211a_1 _15969_ (.A1(_05391_),
    .A2(_05394_),
    .B1(_05050_),
    .C1(_05054_),
    .X(_05399_));
 sky130_fd_sc_hd__a211oi_2 _15970_ (.A1(_05050_),
    .A2(_05054_),
    .B1(_05391_),
    .C1(_05394_),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_1 _15971_ (.A(_05397_),
    .B(_05398_),
    .Y(_05401_));
 sky130_fd_sc_hd__o2bb2ai_4 _15972_ (.A1_N(_05353_),
    .A2_N(_05356_),
    .B1(_05399_),
    .B2(_05400_),
    .Y(_05402_));
 sky130_fd_sc_hd__nand2_1 _15973_ (.A(_05353_),
    .B(_05401_),
    .Y(_05404_));
 sky130_fd_sc_hd__o211ai_2 _15974_ (.A1(_05350_),
    .A2(_05354_),
    .B1(_05401_),
    .C1(_05353_),
    .Y(_05405_));
 sky130_fd_sc_hd__o211a_1 _15975_ (.A1(_05355_),
    .A2(_05404_),
    .B1(_05262_),
    .C1(_05402_),
    .X(_05406_));
 sky130_fd_sc_hd__o211ai_4 _15976_ (.A1(_05355_),
    .A2(_05404_),
    .B1(_05262_),
    .C1(_05402_),
    .Y(_05407_));
 sky130_fd_sc_hd__a21oi_4 _15977_ (.A1(_05402_),
    .A2(_05405_),
    .B1(_05262_),
    .Y(_05408_));
 sky130_fd_sc_hd__a21o_1 _15978_ (.A1(_05402_),
    .A2(_05405_),
    .B1(_05262_),
    .X(_05409_));
 sky130_fd_sc_hd__o21ai_2 _15979_ (.A1(_05406_),
    .A2(_05408_),
    .B1(_05259_),
    .Y(_05410_));
 sky130_fd_sc_hd__o211ai_4 _15980_ (.A1(_05255_),
    .A2(_05257_),
    .B1(_05407_),
    .C1(_05409_),
    .Y(_05411_));
 sky130_fd_sc_hd__o22ai_2 _15981_ (.A1(_05255_),
    .A2(_05257_),
    .B1(_05406_),
    .B2(_05408_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand3_1 _15982_ (.A(_05409_),
    .B(_05259_),
    .C(_05407_),
    .Y(_05413_));
 sky130_fd_sc_hd__a32oi_4 _15983_ (.A1(_05162_),
    .A2(_05164_),
    .A3(_05165_),
    .B1(_05167_),
    .B2(_05016_),
    .Y(_05415_));
 sky130_fd_sc_hd__a21oi_2 _15984_ (.A1(_05015_),
    .A2(_05168_),
    .B1(_05166_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21oi_2 _15985_ (.A1(_05412_),
    .A2(_05413_),
    .B1(_05415_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand3_1 _15986_ (.A(_05410_),
    .B(_05411_),
    .C(_05416_),
    .Y(_05418_));
 sky130_fd_sc_hd__a21oi_2 _15987_ (.A1(_05410_),
    .A2(_05411_),
    .B1(_05416_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand3_2 _15988_ (.A(_05412_),
    .B(_05415_),
    .C(_05413_),
    .Y(_05420_));
 sky130_fd_sc_hd__and2_1 _15989_ (.A(_05010_),
    .B(_05014_),
    .X(_05421_));
 sky130_fd_sc_hd__a21oi_2 _15990_ (.A1(_05010_),
    .A2(_05014_),
    .B1(_05002_),
    .Y(_05422_));
 sky130_fd_sc_hd__a21o_1 _15991_ (.A1(_05010_),
    .A2(_05014_),
    .B1(_05002_),
    .X(_05423_));
 sky130_fd_sc_hd__and3_1 _15992_ (.A(_05002_),
    .B(_05010_),
    .C(_05014_),
    .X(_05424_));
 sky130_fd_sc_hd__or2_2 _15993_ (.A(_05422_),
    .B(_05424_),
    .X(_05426_));
 sky130_fd_sc_hd__o21ai_1 _15994_ (.A1(_05417_),
    .A2(_05419_),
    .B1(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__a31o_1 _15995_ (.A1(_05410_),
    .A2(_05411_),
    .A3(_05416_),
    .B1(_05426_),
    .X(_05428_));
 sky130_fd_sc_hd__o211ai_2 _15996_ (.A1(_05422_),
    .A2(_05424_),
    .B1(_05418_),
    .C1(_05420_),
    .Y(_05429_));
 sky130_fd_sc_hd__a21o_1 _15997_ (.A1(_05418_),
    .A2(_05420_),
    .B1(_05426_),
    .X(_05430_));
 sky130_fd_sc_hd__o221ai_4 _15998_ (.A1(_05173_),
    .A2(_05181_),
    .B1(_05419_),
    .B2(_05428_),
    .C1(_05427_),
    .Y(_05431_));
 sky130_fd_sc_hd__inv_2 _15999_ (.A(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__o211a_1 _16000_ (.A1(_05176_),
    .A2(_05180_),
    .B1(_05429_),
    .C1(_05430_),
    .X(_05433_));
 sky130_fd_sc_hd__o211ai_1 _16001_ (.A1(_05176_),
    .A2(_05180_),
    .B1(_05429_),
    .C1(_05430_),
    .Y(_05434_));
 sky130_fd_sc_hd__nand2_1 _16002_ (.A(_05431_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__a32o_1 _16003_ (.A1(_04946_),
    .A2(_05177_),
    .A3(_05178_),
    .B1(_05431_),
    .B2(_05434_),
    .X(_05437_));
 sky130_fd_sc_hd__nand4_1 _16004_ (.A(_04946_),
    .B(_05177_),
    .C(_05178_),
    .D(_05431_),
    .Y(_05438_));
 sky130_fd_sc_hd__nor2_1 _16005_ (.A(_05183_),
    .B(_05435_),
    .Y(_05439_));
 sky130_fd_sc_hd__or2_1 _16006_ (.A(_05183_),
    .B(_05435_),
    .X(_05440_));
 sky130_fd_sc_hd__o21ai_1 _16007_ (.A1(_05438_),
    .A2(_05433_),
    .B1(_05437_),
    .Y(_05441_));
 sky130_fd_sc_hd__o221a_1 _16008_ (.A1(_05438_),
    .A2(_05433_),
    .B1(_05186_),
    .B2(_04930_),
    .C1(_05437_),
    .X(_05442_));
 sky130_fd_sc_hd__a41o_1 _16009_ (.A1(_04929_),
    .A2(_05183_),
    .A3(_05184_),
    .A4(_05435_),
    .B1(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__xor2_1 _16010_ (.A(_05191_),
    .B(_05443_),
    .X(net78));
 sky130_fd_sc_hd__o32ai_2 _16011_ (.A1(_04932_),
    .A2(_05186_),
    .A3(_05441_),
    .B1(_05435_),
    .B2(_05189_),
    .Y(_05444_));
 sky130_fd_sc_hd__nor3_2 _16012_ (.A(_05187_),
    .B(_05441_),
    .C(_05188_),
    .Y(_05445_));
 sky130_fd_sc_hd__a21oi_1 _16013_ (.A1(_04944_),
    .A2(_05445_),
    .B1(_05444_),
    .Y(_05447_));
 sky130_fd_sc_hd__o21ai_1 _16014_ (.A1(_05261_),
    .A2(_05408_),
    .B1(_05407_),
    .Y(_05448_));
 sky130_fd_sc_hd__o22ai_4 _16015_ (.A1(_05388_),
    .A2(_05393_),
    .B1(_05396_),
    .B2(_05391_),
    .Y(_05449_));
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(_05236_),
    .B(_05239_),
    .Y(_05450_));
 sky130_fd_sc_hd__a32o_1 _16017_ (.A1(_04985_),
    .A2(_04452_),
    .A3(net318),
    .B1(net23),
    .B2(_04988_),
    .X(_05451_));
 sky130_fd_sc_hd__a32o_1 _16018_ (.A1(net266),
    .A2(net303),
    .A3(net279),
    .B1(_04482_),
    .B2(net27),
    .X(_05452_));
 sky130_fd_sc_hd__o32a_1 _16019_ (.A1(_04896_),
    .A2(net306),
    .A3(_04703_),
    .B1(_03506_),
    .B2(_04898_),
    .X(_05453_));
 sky130_fd_sc_hd__a32o_1 _16020_ (.A1(net243),
    .A2(_04747_),
    .A3(net315),
    .B1(net26),
    .B2(_04897_),
    .X(_05454_));
 sky130_fd_sc_hd__nand2_1 _16021_ (.A(_05452_),
    .B(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__o221ai_4 _16022_ (.A1(_05020_),
    .A2(_04481_),
    .B1(_04483_),
    .B2(_03616_),
    .C1(_05453_),
    .Y(_05456_));
 sky130_fd_sc_hd__nand3_1 _16023_ (.A(_05451_),
    .B(_05455_),
    .C(_05456_),
    .Y(_05458_));
 sky130_fd_sc_hd__a21o_1 _16024_ (.A1(_05455_),
    .A2(_05456_),
    .B1(_05451_),
    .X(_05459_));
 sky130_fd_sc_hd__a21o_1 _16025_ (.A1(_05458_),
    .A2(_05459_),
    .B1(_05450_),
    .X(_05460_));
 sky130_fd_sc_hd__nand3_2 _16026_ (.A(_05450_),
    .B(_05458_),
    .C(_05459_),
    .Y(_05461_));
 sky130_fd_sc_hd__and2b_4 _16027_ (.A_N(net46),
    .B(net47),
    .X(_05462_));
 sky130_fd_sc_hd__nand2b_4 _16028_ (.A_N(net46),
    .B(net47),
    .Y(_05463_));
 sky130_fd_sc_hd__and2b_4 _16029_ (.A_N(net47),
    .B(net46),
    .X(_05464_));
 sky130_fd_sc_hd__nand2b_4 _16030_ (.A_N(net47),
    .B(net46),
    .Y(_05465_));
 sky130_fd_sc_hd__a21oi_2 _16031_ (.A1(_05463_),
    .A2(_05465_),
    .B1(_03176_),
    .Y(_05466_));
 sky130_fd_sc_hd__a22o_1 _16032_ (.A1(net12),
    .A2(_05228_),
    .B1(_04539_),
    .B2(net276),
    .X(_05467_));
 sky130_fd_sc_hd__nand2_2 _16033_ (.A(_05467_),
    .B(_05466_),
    .Y(_05469_));
 sky130_fd_sc_hd__a221o_1 _16034_ (.A1(_04539_),
    .A2(net276),
    .B1(_05228_),
    .B2(net12),
    .C1(_05466_),
    .X(_05470_));
 sky130_fd_sc_hd__and4_2 _16035_ (.A(_05460_),
    .B(_05461_),
    .C(_05469_),
    .D(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__a22oi_2 _16036_ (.A1(_05460_),
    .A2(_05461_),
    .B1(_05469_),
    .B2(_05470_),
    .Y(_05472_));
 sky130_fd_sc_hd__nor2_1 _16037_ (.A(_05471_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__a21oi_1 _16038_ (.A1(_05193_),
    .A2(_05215_),
    .B1(_05213_),
    .Y(_05474_));
 sky130_fd_sc_hd__nor2_1 _16039_ (.A(_03916_),
    .B(_03737_),
    .Y(_05475_));
 sky130_fd_sc_hd__a31o_1 _16040_ (.A1(_06486_),
    .A2(net261),
    .A3(net285),
    .B1(_05475_),
    .X(_05476_));
 sky130_fd_sc_hd__nor2_1 _16041_ (.A(_03835_),
    .B(_04218_),
    .Y(_05477_));
 sky130_fd_sc_hd__a31oi_1 _16042_ (.A1(_05841_),
    .A2(net265),
    .A3(_04215_),
    .B1(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__a31o_1 _16043_ (.A1(_05841_),
    .A2(net265),
    .A3(_04215_),
    .B1(_05477_),
    .X(_05480_));
 sky130_fd_sc_hd__o221ai_2 _16044_ (.A1(_06552_),
    .A2(_03714_),
    .B1(_03737_),
    .B2(_03916_),
    .C1(_05478_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(_05476_),
    .B(_05480_),
    .Y(_05482_));
 sky130_fd_sc_hd__a32o_1 _16046_ (.A1(_05414_),
    .A2(_05446_),
    .A3(net280),
    .B1(_04269_),
    .B2(net28),
    .X(_05483_));
 sky130_fd_sc_hd__a21o_1 _16047_ (.A1(_05481_),
    .A2(_05482_),
    .B1(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__nand3_2 _16048_ (.A(_05481_),
    .B(_05482_),
    .C(_05483_),
    .Y(_05485_));
 sky130_fd_sc_hd__a31oi_2 _16049_ (.A1(_05361_),
    .A2(_05362_),
    .A3(_05363_),
    .B1(_05357_),
    .Y(_05486_));
 sky130_fd_sc_hd__a21o_1 _16050_ (.A1(_05358_),
    .A2(_05366_),
    .B1(_05364_),
    .X(_05487_));
 sky130_fd_sc_hd__a21oi_2 _16051_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__o211a_1 _16052_ (.A1(_05364_),
    .A2(_05486_),
    .B1(_05485_),
    .C1(_05484_),
    .X(_05489_));
 sky130_fd_sc_hd__o211ai_4 _16053_ (.A1(_05364_),
    .A2(_05486_),
    .B1(_05485_),
    .C1(_05484_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_2 _16054_ (.A1(_05488_),
    .A2(_05489_),
    .B1(_05211_),
    .Y(_05492_));
 sky130_fd_sc_hd__nor2_1 _16055_ (.A(_05211_),
    .B(_05488_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand3b_2 _16056_ (.A_N(_05488_),
    .B(_05491_),
    .C(_05210_),
    .Y(_05494_));
 sky130_fd_sc_hd__a21boi_1 _16057_ (.A1(_05492_),
    .A2(_05494_),
    .B1_N(_05474_),
    .Y(_05495_));
 sky130_fd_sc_hd__a21bo_1 _16058_ (.A1(_05492_),
    .A2(_05494_),
    .B1_N(_05474_),
    .X(_05496_));
 sky130_fd_sc_hd__o211a_1 _16059_ (.A1(_05213_),
    .A2(_05219_),
    .B1(_05492_),
    .C1(_05494_),
    .X(_05497_));
 sky130_fd_sc_hd__o211ai_1 _16060_ (.A1(_05213_),
    .A2(_05219_),
    .B1(_05492_),
    .C1(_05494_),
    .Y(_05498_));
 sky130_fd_sc_hd__o22ai_2 _16061_ (.A1(_05471_),
    .A2(_05472_),
    .B1(_05495_),
    .B2(_05497_),
    .Y(_05499_));
 sky130_fd_sc_hd__nand3_2 _16062_ (.A(_05496_),
    .B(_05498_),
    .C(_05473_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand3_4 _16063_ (.A(_05499_),
    .B(_05500_),
    .C(_05449_),
    .Y(_05502_));
 sky130_fd_sc_hd__a21o_1 _16064_ (.A1(_05499_),
    .A2(_05500_),
    .B1(_05449_),
    .X(_05503_));
 sky130_fd_sc_hd__o31a_1 _16065_ (.A1(_05223_),
    .A2(_05246_),
    .A3(_05247_),
    .B1(_05222_),
    .X(_05504_));
 sky130_fd_sc_hd__a22o_1 _16066_ (.A1(_05224_),
    .A2(_05250_),
    .B1(_05502_),
    .B2(_05503_),
    .X(_05505_));
 sky130_fd_sc_hd__nand4_2 _16067_ (.A(_05224_),
    .B(_05250_),
    .C(_05502_),
    .D(_05503_),
    .Y(_05506_));
 sky130_fd_sc_hd__a21o_1 _16068_ (.A1(_05502_),
    .A2(_05503_),
    .B1(_05504_),
    .X(_05507_));
 sky130_fd_sc_hd__nand3_4 _16069_ (.A(_05502_),
    .B(_05503_),
    .C(_05504_),
    .Y(_05508_));
 sky130_fd_sc_hd__nand2_1 _16070_ (.A(_05507_),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(_05505_),
    .B(_05506_),
    .Y(_05510_));
 sky130_fd_sc_hd__a21boi_1 _16072_ (.A1(_05320_),
    .A2(_05346_),
    .B1_N(_05319_),
    .Y(_05511_));
 sky130_fd_sc_hd__o2bb2ai_2 _16073_ (.A1_N(_05346_),
    .A2_N(_05320_),
    .B1(_05316_),
    .B2(_05318_),
    .Y(_05513_));
 sky130_fd_sc_hd__a21oi_1 _16074_ (.A1(_05325_),
    .A2(_05328_),
    .B1(_05334_),
    .Y(_05514_));
 sky130_fd_sc_hd__o21ai_2 _16075_ (.A1(_05269_),
    .A2(_05273_),
    .B1(_05266_),
    .Y(_05515_));
 sky130_fd_sc_hd__a21oi_1 _16076_ (.A1(_05269_),
    .A2(_05273_),
    .B1(_05266_),
    .Y(_05516_));
 sky130_fd_sc_hd__a32o_2 _16077_ (.A1(_02421_),
    .A2(net249),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net6),
    .X(_05517_));
 sky130_fd_sc_hd__nand3_2 _16078_ (.A(_04132_),
    .B(net299),
    .C(net230),
    .Y(_05518_));
 sky130_fd_sc_hd__or3b_1 _16079_ (.A(net61),
    .B(_04059_),
    .C_N(net60),
    .X(_05519_));
 sky130_fd_sc_hd__and3_1 _16080_ (.A(_03927_),
    .B(net7),
    .C(net61),
    .X(_05520_));
 sky130_fd_sc_hd__o21ai_1 _16081_ (.A1(net263),
    .A2(net246),
    .B1(net292),
    .Y(_05521_));
 sky130_fd_sc_hd__a21oi_1 _16082_ (.A1(net7),
    .A2(net249),
    .B1(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__o22a_1 _16083_ (.A1(_04048_),
    .A2(_06859_),
    .B1(net247),
    .B2(_05521_),
    .X(_05524_));
 sky130_fd_sc_hd__o211ai_4 _16084_ (.A1(_04059_),
    .A2(net298),
    .B1(_05518_),
    .C1(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__o2bb2ai_2 _16085_ (.A1_N(_05518_),
    .A2_N(_05519_),
    .B1(_05520_),
    .B2(_05522_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand3b_1 _16086_ (.A_N(_05517_),
    .B(_05525_),
    .C(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21bo_1 _16087_ (.A1(_05525_),
    .A2(_05526_),
    .B1_N(_05517_),
    .X(_05528_));
 sky130_fd_sc_hd__a21boi_4 _16088_ (.A1(_05517_),
    .A2(_05525_),
    .B1_N(_05526_),
    .Y(_05529_));
 sky130_fd_sc_hd__a21o_1 _16089_ (.A1(_05525_),
    .A2(_05526_),
    .B1(_05517_),
    .X(_05530_));
 sky130_fd_sc_hd__nand3_2 _16090_ (.A(_05517_),
    .B(_05525_),
    .C(_05526_),
    .Y(_05531_));
 sky130_fd_sc_hd__a22oi_4 _16091_ (.A1(_05277_),
    .A2(_05515_),
    .B1(_05530_),
    .B2(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__a22o_1 _16092_ (.A1(_05277_),
    .A2(_05515_),
    .B1(_05530_),
    .B2(_05531_),
    .X(_05533_));
 sky130_fd_sc_hd__a2bb2oi_1 _16093_ (.A1_N(_05274_),
    .A2_N(_05516_),
    .B1(_05527_),
    .B2(_05528_),
    .Y(_05535_));
 sky130_fd_sc_hd__nand4_2 _16094_ (.A(_05277_),
    .B(_05515_),
    .C(_05530_),
    .D(_05531_),
    .Y(_05536_));
 sky130_fd_sc_hd__o2bb2a_1 _16095_ (.A1_N(_05329_),
    .A2_N(_05335_),
    .B1(_05532_),
    .B2(_05535_),
    .X(_05537_));
 sky130_fd_sc_hd__a22o_1 _16096_ (.A1(_05329_),
    .A2(_05335_),
    .B1(_05533_),
    .B2(_05536_),
    .X(_05538_));
 sky130_fd_sc_hd__and3_1 _16097_ (.A(_05533_),
    .B(_05536_),
    .C(_05514_),
    .X(_05539_));
 sky130_fd_sc_hd__nand4_2 _16098_ (.A(_05329_),
    .B(_05335_),
    .C(_05533_),
    .D(_05536_),
    .Y(_05540_));
 sky130_fd_sc_hd__o21ai_1 _16099_ (.A1(_05532_),
    .A2(_05535_),
    .B1(_05514_),
    .Y(_05541_));
 sky130_fd_sc_hd__a211o_1 _16100_ (.A1(_05329_),
    .A2(_05335_),
    .B1(_05532_),
    .C1(_05535_),
    .X(_05542_));
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(_05538_),
    .B(_05540_),
    .Y(_05543_));
 sky130_fd_sc_hd__a21oi_1 _16102_ (.A1(_05283_),
    .A2(_05308_),
    .B1(_05309_),
    .Y(_05544_));
 sky130_fd_sc_hd__a22o_1 _16103_ (.A1(_04135_),
    .A2(_05297_),
    .B1(_05300_),
    .B2(_05289_),
    .X(_05546_));
 sky130_fd_sc_hd__a21oi_2 _16104_ (.A1(_05289_),
    .A2(_05300_),
    .B1(_05301_),
    .Y(_05547_));
 sky130_fd_sc_hd__a41oi_4 _16105_ (.A1(_06519_),
    .A2(_03955_),
    .A3(net277),
    .A4(_05291_),
    .B1(_04146_),
    .Y(_05548_));
 sky130_fd_sc_hd__a41o_4 _16106_ (.A1(_06519_),
    .A2(_03955_),
    .A3(_04786_),
    .A4(_05291_),
    .B1(_04146_),
    .X(_05549_));
 sky130_fd_sc_hd__and3_4 _16107_ (.A(_04113_),
    .B(_04135_),
    .C(_04146_),
    .X(_05550_));
 sky130_fd_sc_hd__nand2_8 _16108_ (.A(_05291_),
    .B(_04146_),
    .Y(_05551_));
 sky130_fd_sc_hd__nor4_2 _16109_ (.A(net262),
    .B(net245),
    .C(_04787_),
    .D(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand4_4 _16110_ (.A(_06519_),
    .B(_03955_),
    .C(net277),
    .D(_05550_),
    .Y(_05553_));
 sky130_fd_sc_hd__o21ai_4 _16111_ (.A1(_04789_),
    .A2(_05551_),
    .B1(_05549_),
    .Y(_05554_));
 sky130_fd_sc_hd__o211ai_2 _16112_ (.A1(net185),
    .A2(_05551_),
    .B1(net33),
    .C1(_05549_),
    .Y(_05555_));
 sky130_fd_sc_hd__nand3_1 _16113_ (.A(net181),
    .B(net180),
    .C(_04484_),
    .Y(_05557_));
 sky130_fd_sc_hd__or3_1 _16114_ (.A(net44),
    .B(_04135_),
    .C(_03286_),
    .X(_05558_));
 sky130_fd_sc_hd__and4b_1 _16115_ (.A_N(net44),
    .B(_04146_),
    .C(net14),
    .D(net33),
    .X(_05559_));
 sky130_fd_sc_hd__or4_2 _16116_ (.A(net44),
    .B(net15),
    .C(_04135_),
    .D(_03286_),
    .X(_05560_));
 sky130_fd_sc_hd__nand3_4 _16117_ (.A(_05555_),
    .B(_05557_),
    .C(_05558_),
    .Y(_05561_));
 sky130_fd_sc_hd__o41ai_1 _16118_ (.A1(_03286_),
    .A2(net44),
    .A3(_04135_),
    .A4(net15),
    .B1(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__nor2_1 _16119_ (.A(_04113_),
    .B(_04375_),
    .Y(_05563_));
 sky130_fd_sc_hd__o311a_1 _16120_ (.A1(net11),
    .A2(_04557_),
    .A3(_05073_),
    .B1(_04342_),
    .C1(net212),
    .X(_05564_));
 sky130_fd_sc_hd__a31oi_2 _16121_ (.A1(net212),
    .A2(net183),
    .A3(_04342_),
    .B1(_05563_),
    .Y(_05565_));
 sky130_fd_sc_hd__a31o_1 _16122_ (.A1(net212),
    .A2(net183),
    .A3(_04342_),
    .B1(_05563_),
    .X(_05566_));
 sky130_fd_sc_hd__o2bb2ai_2 _16123_ (.A1_N(_05560_),
    .A2_N(_05561_),
    .B1(_05563_),
    .B2(_05564_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand3_2 _16124_ (.A(_05560_),
    .B(_05561_),
    .C(_05565_),
    .Y(_05569_));
 sky130_fd_sc_hd__o221a_1 _16125_ (.A1(_04113_),
    .A2(_04375_),
    .B1(_05077_),
    .B2(_04353_),
    .C1(_05562_),
    .X(_05570_));
 sky130_fd_sc_hd__nand2_1 _16126_ (.A(_05562_),
    .B(_05565_),
    .Y(_05571_));
 sky130_fd_sc_hd__a311o_1 _16127_ (.A1(_05555_),
    .A2(_05557_),
    .A3(_05558_),
    .B1(_05559_),
    .C1(_05565_),
    .X(_05572_));
 sky130_fd_sc_hd__a32o_1 _16128_ (.A1(_05560_),
    .A2(_05561_),
    .A3(_05566_),
    .B1(_05307_),
    .B2(_05302_),
    .X(_05573_));
 sky130_fd_sc_hd__a21oi_2 _16129_ (.A1(_05568_),
    .A2(_05569_),
    .B1(_05547_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand3_4 _16130_ (.A(_05571_),
    .B(_05572_),
    .C(_05546_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand3_4 _16131_ (.A(_05547_),
    .B(_05568_),
    .C(_05569_),
    .Y(_05576_));
 sky130_fd_sc_hd__inv_2 _16132_ (.A(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__o21ai_1 _16133_ (.A1(_05570_),
    .A2(_05573_),
    .B1(_05576_),
    .Y(_05579_));
 sky130_fd_sc_hd__a32oi_4 _16134_ (.A1(net224),
    .A2(_05227_),
    .A3(net188),
    .B1(_05249_),
    .B2(net9),
    .Y(_05580_));
 sky130_fd_sc_hd__or3b_2 _16135_ (.A(net58),
    .B(_04091_),
    .C_N(net55),
    .X(_05581_));
 sky130_fd_sc_hd__o221ai_4 _16136_ (.A1(net232),
    .A2(_04787_),
    .B1(_04091_),
    .B2(_04558_),
    .C1(net317),
    .Y(_05582_));
 sky130_fd_sc_hd__a31oi_2 _16137_ (.A1(_11420_),
    .A2(net282),
    .A3(_04556_),
    .B1(_04900_),
    .Y(_05583_));
 sky130_fd_sc_hd__a22oi_4 _16138_ (.A1(net10),
    .A2(_04911_),
    .B1(_05583_),
    .B2(_04555_),
    .Y(_05584_));
 sky130_fd_sc_hd__a21oi_4 _16139_ (.A1(_05581_),
    .A2(_05582_),
    .B1(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__a21o_1 _16140_ (.A1(_05581_),
    .A2(_05582_),
    .B1(_05584_),
    .X(_05586_));
 sky130_fd_sc_hd__o211a_2 _16141_ (.A1(_04091_),
    .A2(net316),
    .B1(_05582_),
    .C1(_05584_),
    .X(_05587_));
 sky130_fd_sc_hd__o211ai_1 _16142_ (.A1(_04091_),
    .A2(net316),
    .B1(_05582_),
    .C1(_05584_),
    .Y(_05588_));
 sky130_fd_sc_hd__a31o_1 _16143_ (.A1(_05584_),
    .A2(_05582_),
    .A3(_05581_),
    .B1(_05580_),
    .X(_05590_));
 sky130_fd_sc_hd__o21ai_2 _16144_ (.A1(_05580_),
    .A2(_05587_),
    .B1(_05586_),
    .Y(_05591_));
 sky130_fd_sc_hd__nor2_1 _16145_ (.A(_05585_),
    .B(_05590_),
    .Y(_05592_));
 sky130_fd_sc_hd__a21oi_1 _16146_ (.A1(_05586_),
    .A2(_05588_),
    .B1(_05580_),
    .Y(_05593_));
 sky130_fd_sc_hd__and3_1 _16147_ (.A(_05586_),
    .B(_05588_),
    .C(_05580_),
    .X(_05594_));
 sky130_fd_sc_hd__o21a_1 _16148_ (.A1(_05585_),
    .A2(_05587_),
    .B1(_05580_),
    .X(_05595_));
 sky130_fd_sc_hd__o21ai_2 _16149_ (.A1(_05585_),
    .A2(_05587_),
    .B1(_05580_),
    .Y(_05596_));
 sky130_fd_sc_hd__o21ai_1 _16150_ (.A1(_05585_),
    .A2(_05590_),
    .B1(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__o2bb2ai_1 _16151_ (.A1_N(_05575_),
    .A2_N(_05576_),
    .B1(_05593_),
    .B2(_05594_),
    .Y(_05598_));
 sky130_fd_sc_hd__o211ai_2 _16152_ (.A1(_05592_),
    .A2(_05595_),
    .B1(_05575_),
    .C1(_05576_),
    .Y(_05599_));
 sky130_fd_sc_hd__o21a_1 _16153_ (.A1(_05592_),
    .A2(_05595_),
    .B1(_05575_),
    .X(_05601_));
 sky130_fd_sc_hd__o211ai_4 _16154_ (.A1(_05585_),
    .A2(_05590_),
    .B1(_05596_),
    .C1(_05576_),
    .Y(_05602_));
 sky130_fd_sc_hd__o21ai_2 _16155_ (.A1(_05570_),
    .A2(_05573_),
    .B1(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__o21a_1 _16156_ (.A1(_05570_),
    .A2(_05573_),
    .B1(_05602_),
    .X(_05604_));
 sky130_fd_sc_hd__o2bb2ai_2 _16157_ (.A1_N(_05575_),
    .A2_N(_05576_),
    .B1(_05592_),
    .B2(_05595_),
    .Y(_05605_));
 sky130_fd_sc_hd__o211ai_2 _16158_ (.A1(_05593_),
    .A2(_05594_),
    .B1(_05575_),
    .C1(_05576_),
    .Y(_05606_));
 sky130_fd_sc_hd__nand3_4 _16159_ (.A(_05544_),
    .B(_05598_),
    .C(_05599_),
    .Y(_05607_));
 sky130_fd_sc_hd__inv_2 _16160_ (.A(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__a22oi_2 _16161_ (.A1(_05310_),
    .A2(_05314_),
    .B1(_05579_),
    .B2(_05597_),
    .Y(_05609_));
 sky130_fd_sc_hd__o221a_2 _16162_ (.A1(_05309_),
    .A2(_05313_),
    .B1(_05574_),
    .B2(_05602_),
    .C1(_05605_),
    .X(_05610_));
 sky130_fd_sc_hd__o221ai_4 _16163_ (.A1(_05309_),
    .A2(_05313_),
    .B1(_05574_),
    .B2(_05602_),
    .C1(_05605_),
    .Y(_05612_));
 sky130_fd_sc_hd__a22o_1 _16164_ (.A1(_05538_),
    .A2(_05540_),
    .B1(_05607_),
    .B2(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__a21oi_2 _16165_ (.A1(_05609_),
    .A2(_05606_),
    .B1(_05543_),
    .Y(_05614_));
 sky130_fd_sc_hd__nand4_2 _16166_ (.A(_05538_),
    .B(_05540_),
    .C(_05607_),
    .D(_05612_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_2 _16167_ (.A1(_05537_),
    .A2(_05539_),
    .B1(_05607_),
    .Y(_05616_));
 sky130_fd_sc_hd__a22o_1 _16168_ (.A1(_05541_),
    .A2(_05542_),
    .B1(_05607_),
    .B2(_05612_),
    .X(_05617_));
 sky130_fd_sc_hd__o211a_1 _16169_ (.A1(_05616_),
    .A2(_05610_),
    .B1(_05513_),
    .C1(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__o211ai_4 _16170_ (.A1(_05616_),
    .A2(_05610_),
    .B1(_05513_),
    .C1(_05617_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand3_4 _16171_ (.A(_05511_),
    .B(_05613_),
    .C(_05615_),
    .Y(_05620_));
 sky130_fd_sc_hd__o31a_2 _16172_ (.A1(_05367_),
    .A2(_05368_),
    .A3(_05385_),
    .B1(_05384_),
    .X(_05621_));
 sky130_fd_sc_hd__a31oi_2 _16173_ (.A1(_05109_),
    .A2(_05333_),
    .A3(_05335_),
    .B1(_05322_),
    .Y(_05623_));
 sky130_fd_sc_hd__a31o_1 _16174_ (.A1(_05109_),
    .A2(_05333_),
    .A3(_05335_),
    .B1(_05322_),
    .X(_05624_));
 sky130_fd_sc_hd__a32o_1 _16175_ (.A1(_07242_),
    .A2(net257),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net31),
    .X(_05625_));
 sky130_fd_sc_hd__a31oi_2 _16176_ (.A1(net310),
    .A2(net294),
    .A3(net290),
    .B1(_12341_),
    .Y(_05626_));
 sky130_fd_sc_hd__a22oi_2 _16177_ (.A1(net2),
    .A2(_12352_),
    .B1(_09698_),
    .B2(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__o211ai_2 _16178_ (.A1(net261),
    .A2(_08656_),
    .B1(_01293_),
    .C1(_08700_),
    .Y(_05628_));
 sky130_fd_sc_hd__or3b_1 _16179_ (.A(_03949_),
    .B(net37),
    .C_N(net36),
    .X(_05629_));
 sky130_fd_sc_hd__a21oi_1 _16180_ (.A1(_05628_),
    .A2(_05629_),
    .B1(_05627_),
    .Y(_05630_));
 sky130_fd_sc_hd__a21o_1 _16181_ (.A1(_05628_),
    .A2(_05629_),
    .B1(_05627_),
    .X(_05631_));
 sky130_fd_sc_hd__o211ai_2 _16182_ (.A1(_03949_),
    .A2(_01326_),
    .B1(_05628_),
    .C1(_05627_),
    .Y(_05632_));
 sky130_fd_sc_hd__a21oi_2 _16183_ (.A1(_05631_),
    .A2(_05632_),
    .B1(_05625_),
    .Y(_05634_));
 sky130_fd_sc_hd__and3_1 _16184_ (.A(_05625_),
    .B(_05631_),
    .C(_05632_),
    .X(_05635_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_05634_),
    .B(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__o221a_1 _16186_ (.A1(_09720_),
    .A2(_11782_),
    .B1(_11804_),
    .B2(_03960_),
    .C1(_05377_),
    .X(_05637_));
 sky130_fd_sc_hd__nor2_1 _16187_ (.A(_05371_),
    .B(_05378_),
    .Y(_05638_));
 sky130_fd_sc_hd__a32o_2 _16188_ (.A1(_11354_),
    .A2(net254),
    .A3(net252),
    .B1(_11793_),
    .B2(net3),
    .X(_05639_));
 sky130_fd_sc_hd__or3b_1 _16189_ (.A(net64),
    .B(_04015_),
    .C_N(net63),
    .X(_05640_));
 sky130_fd_sc_hd__o211ai_2 _16190_ (.A1(net254),
    .A2(_00646_),
    .B1(net291),
    .C1(_00625_),
    .Y(_05641_));
 sky130_fd_sc_hd__a32oi_4 _16191_ (.A1(net235),
    .A2(net251),
    .A3(net289),
    .B1(_10335_),
    .B2(net4),
    .Y(_05642_));
 sky130_fd_sc_hd__o211a_1 _16192_ (.A1(_04015_),
    .A2(_08283_),
    .B1(_05641_),
    .C1(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__o221ai_4 _16193_ (.A1(_04015_),
    .A2(_08283_),
    .B1(_00668_),
    .B2(_08261_),
    .C1(_05642_),
    .Y(_05645_));
 sky130_fd_sc_hd__a21oi_2 _16194_ (.A1(_05640_),
    .A2(_05641_),
    .B1(_05642_),
    .Y(_05646_));
 sky130_fd_sc_hd__a21o_1 _16195_ (.A1(_05640_),
    .A2(_05641_),
    .B1(_05642_),
    .X(_05647_));
 sky130_fd_sc_hd__nand3b_2 _16196_ (.A_N(_05639_),
    .B(_05645_),
    .C(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_2 _16197_ (.A1(_05643_),
    .A2(_05646_),
    .B1(_05639_),
    .Y(_05649_));
 sky130_fd_sc_hd__o221a_1 _16198_ (.A1(net236),
    .A2(_11782_),
    .B1(_11804_),
    .B2(_03982_),
    .C1(_05647_),
    .X(_05650_));
 sky130_fd_sc_hd__a21o_1 _16199_ (.A1(_05645_),
    .A2(_05647_),
    .B1(_05639_),
    .X(_05651_));
 sky130_fd_sc_hd__nand3_1 _16200_ (.A(_05639_),
    .B(_05645_),
    .C(_05647_),
    .Y(_05652_));
 sky130_fd_sc_hd__a2bb2oi_2 _16201_ (.A1_N(_05376_),
    .A2_N(_05638_),
    .B1(_05648_),
    .B2(_05649_),
    .Y(_05653_));
 sky130_fd_sc_hd__o211ai_2 _16202_ (.A1(_05376_),
    .A2(_05638_),
    .B1(_05651_),
    .C1(_05652_),
    .Y(_05654_));
 sky130_fd_sc_hd__o211a_1 _16203_ (.A1(_05378_),
    .A2(_05637_),
    .B1(_05648_),
    .C1(_05649_),
    .X(_05656_));
 sky130_fd_sc_hd__o211ai_2 _16204_ (.A1(_05378_),
    .A2(_05637_),
    .B1(_05648_),
    .C1(_05649_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand3_4 _16205_ (.A(_05654_),
    .B(_05657_),
    .C(_05636_),
    .Y(_05658_));
 sky130_fd_sc_hd__o22ai_4 _16206_ (.A1(_05634_),
    .A2(_05635_),
    .B1(_05653_),
    .B2(_05656_),
    .Y(_05659_));
 sky130_fd_sc_hd__a2bb2oi_4 _16207_ (.A1_N(_05338_),
    .A2_N(_05623_),
    .B1(_05658_),
    .B2(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__o2111a_1 _16208_ (.A1(_05109_),
    .A2(_05336_),
    .B1(_05624_),
    .C1(_05658_),
    .D1(_05659_),
    .X(_05661_));
 sky130_fd_sc_hd__o2111ai_4 _16209_ (.A1(_05109_),
    .A2(_05336_),
    .B1(_05624_),
    .C1(_05658_),
    .D1(_05659_),
    .Y(_05662_));
 sky130_fd_sc_hd__o211a_1 _16210_ (.A1(_05660_),
    .A2(_05661_),
    .B1(_05384_),
    .C1(_05387_),
    .X(_05663_));
 sky130_fd_sc_hd__a211oi_1 _16211_ (.A1(_05384_),
    .A2(_05387_),
    .B1(_05660_),
    .C1(_05661_),
    .Y(_05664_));
 sky130_fd_sc_hd__o2bb2a_1 _16212_ (.A1_N(_05384_),
    .A2_N(_05387_),
    .B1(_05660_),
    .B2(_05661_),
    .X(_05665_));
 sky130_fd_sc_hd__and3b_1 _16213_ (.A_N(_05660_),
    .B(_05662_),
    .C(_05621_),
    .X(_05667_));
 sky130_fd_sc_hd__o2bb2ai_1 _16214_ (.A1_N(_05619_),
    .A2_N(_05620_),
    .B1(_05663_),
    .B2(_05664_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21a_1 _16215_ (.A1(_05665_),
    .A2(_05667_),
    .B1(_05620_),
    .X(_05669_));
 sky130_fd_sc_hd__o211ai_2 _16216_ (.A1(_05665_),
    .A2(_05667_),
    .B1(_05619_),
    .C1(_05620_),
    .Y(_05670_));
 sky130_fd_sc_hd__o211ai_1 _16217_ (.A1(_05663_),
    .A2(_05664_),
    .B1(_05619_),
    .C1(_05620_),
    .Y(_05671_));
 sky130_fd_sc_hd__o2bb2ai_1 _16218_ (.A1_N(_05619_),
    .A2_N(_05620_),
    .B1(_05665_),
    .B2(_05667_),
    .Y(_05672_));
 sky130_fd_sc_hd__o2bb2ai_1 _16219_ (.A1_N(_05353_),
    .A2_N(_05401_),
    .B1(_05354_),
    .B2(_05350_),
    .Y(_05673_));
 sky130_fd_sc_hd__a21oi_1 _16220_ (.A1(_05353_),
    .A2(_05401_),
    .B1(_05355_),
    .Y(_05674_));
 sky130_fd_sc_hd__and3_1 _16221_ (.A(_05671_),
    .B(_05672_),
    .C(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__nand3_2 _16222_ (.A(_05671_),
    .B(_05672_),
    .C(_05674_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand3_4 _16223_ (.A(_05668_),
    .B(_05673_),
    .C(_05670_),
    .Y(_05678_));
 sky130_fd_sc_hd__nand4_2 _16224_ (.A(_05505_),
    .B(_05506_),
    .C(_05676_),
    .D(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__a22o_1 _16225_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_05676_),
    .B2(_05678_),
    .X(_05680_));
 sky130_fd_sc_hd__nand4_1 _16226_ (.A(_05507_),
    .B(_05508_),
    .C(_05676_),
    .D(_05678_),
    .Y(_05681_));
 sky130_fd_sc_hd__a22o_1 _16227_ (.A1(_05507_),
    .A2(_05508_),
    .B1(_05676_),
    .B2(_05678_),
    .X(_05682_));
 sky130_fd_sc_hd__nand3_2 _16228_ (.A(_05682_),
    .B(_05448_),
    .C(_05681_),
    .Y(_05683_));
 sky130_fd_sc_hd__o2111ai_4 _16229_ (.A1(_05408_),
    .A2(_05261_),
    .B1(_05407_),
    .C1(_05679_),
    .D1(_05680_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21a_2 _16230_ (.A1(_05230_),
    .A2(_05243_),
    .B1(_05241_),
    .X(_05685_));
 sky130_fd_sc_hd__o21a_1 _16231_ (.A1(_05251_),
    .A2(_05252_),
    .B1(_05258_),
    .X(_05686_));
 sky130_fd_sc_hd__a21oi_2 _16232_ (.A1(_05254_),
    .A2(_05258_),
    .B1(_05685_),
    .Y(_05687_));
 sky130_fd_sc_hd__a21o_1 _16233_ (.A1(_05254_),
    .A2(_05258_),
    .B1(_05685_),
    .X(_05689_));
 sky130_fd_sc_hd__and3_1 _16234_ (.A(_05254_),
    .B(_05258_),
    .C(_05685_),
    .X(_05690_));
 sky130_fd_sc_hd__and2b_1 _16235_ (.A_N(_05685_),
    .B(_05686_),
    .X(_05691_));
 sky130_fd_sc_hd__a21boi_1 _16236_ (.A1(_05254_),
    .A2(_05258_),
    .B1_N(_05685_),
    .Y(_05692_));
 sky130_fd_sc_hd__o211ai_2 _16237_ (.A1(_05687_),
    .A2(_05690_),
    .B1(_05683_),
    .C1(_05684_),
    .Y(_05693_));
 sky130_fd_sc_hd__o2bb2ai_1 _16238_ (.A1_N(_05683_),
    .A2_N(_05684_),
    .B1(_05691_),
    .B2(_05692_),
    .Y(_05694_));
 sky130_fd_sc_hd__o2bb2ai_1 _16239_ (.A1_N(_05683_),
    .A2_N(_05684_),
    .B1(_05687_),
    .B2(_05690_),
    .Y(_05695_));
 sky130_fd_sc_hd__o211ai_1 _16240_ (.A1(_05691_),
    .A2(_05692_),
    .B1(_05683_),
    .C1(_05684_),
    .Y(_05696_));
 sky130_fd_sc_hd__a32oi_2 _16241_ (.A1(_05410_),
    .A2(_05411_),
    .A3(_05416_),
    .B1(_05420_),
    .B2(_05426_),
    .Y(_05697_));
 sky130_fd_sc_hd__o2111ai_4 _16242_ (.A1(_05426_),
    .A2(_05417_),
    .B1(_05420_),
    .C1(_05693_),
    .D1(_05694_),
    .Y(_05698_));
 sky130_fd_sc_hd__nand3_2 _16243_ (.A(_05695_),
    .B(_05697_),
    .C(_05696_),
    .Y(_05700_));
 sky130_fd_sc_hd__a2bb2o_1 _16244_ (.A1_N(_05421_),
    .A2_N(_05002_),
    .B1(_05700_),
    .B2(_05698_),
    .X(_05701_));
 sky130_fd_sc_hd__o211ai_1 _16245_ (.A1(_05421_),
    .A2(_05002_),
    .B1(_05700_),
    .C1(_05698_),
    .Y(_05702_));
 sky130_fd_sc_hd__a21o_1 _16246_ (.A1(_05698_),
    .A2(_05700_),
    .B1(_05423_),
    .X(_05703_));
 sky130_fd_sc_hd__nand3_1 _16247_ (.A(_05698_),
    .B(_05700_),
    .C(_05422_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand3_1 _16248_ (.A(_05431_),
    .B(_05702_),
    .C(_05703_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand3_1 _16249_ (.A(_05701_),
    .B(_05704_),
    .C(_05432_),
    .Y(_05706_));
 sky130_fd_sc_hd__inv_2 _16250_ (.A(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand2_1 _16251_ (.A(_05705_),
    .B(_05706_),
    .Y(_05708_));
 sky130_fd_sc_hd__and3_1 _16252_ (.A(_05439_),
    .B(_05701_),
    .C(_05704_),
    .X(_05709_));
 sky130_fd_sc_hd__or4b_1 _16253_ (.A(_05183_),
    .B(_05432_),
    .C(_05433_),
    .D_N(_05705_),
    .X(_05711_));
 sky130_fd_sc_hd__a21oi_2 _16254_ (.A1(_05440_),
    .A2(_05708_),
    .B1(_05709_),
    .Y(_05712_));
 sky130_fd_sc_hd__xnor2_1 _16255_ (.A(_05447_),
    .B(_05712_),
    .Y(net79));
 sky130_fd_sc_hd__o21ai_1 _16256_ (.A1(_05687_),
    .A2(_05690_),
    .B1(_05683_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _16257_ (.A(_05684_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__a32o_1 _16258_ (.A1(_05450_),
    .A2(_05458_),
    .A3(_05459_),
    .B1(_05466_),
    .B2(_05467_),
    .X(_05715_));
 sky130_fd_sc_hd__or2_4 _16259_ (.A(_05461_),
    .B(_05469_),
    .X(_05716_));
 sky130_fd_sc_hd__a21oi_4 _16260_ (.A1(_05715_),
    .A2(_05716_),
    .B1(_05471_),
    .Y(_05717_));
 sky130_fd_sc_hd__and2_1 _16261_ (.A(_05502_),
    .B(_05508_),
    .X(_05718_));
 sky130_fd_sc_hd__a21oi_4 _16262_ (.A1(_05502_),
    .A2(_05508_),
    .B1(_05717_),
    .Y(_05719_));
 sky130_fd_sc_hd__inv_2 _16263_ (.A(_05719_),
    .Y(_05721_));
 sky130_fd_sc_hd__and3_1 _16264_ (.A(_05502_),
    .B(_05508_),
    .C(_05717_),
    .X(_05722_));
 sky130_fd_sc_hd__and2b_1 _16265_ (.A_N(_05717_),
    .B(_05718_),
    .X(_05723_));
 sky130_fd_sc_hd__a221oi_2 _16266_ (.A1(_05502_),
    .A2(_05508_),
    .B1(_05715_),
    .B2(_05716_),
    .C1(_05471_),
    .Y(_05724_));
 sky130_fd_sc_hd__nor2_1 _16267_ (.A(_05719_),
    .B(_05722_),
    .Y(_05725_));
 sky130_fd_sc_hd__and3_1 _16268_ (.A(_05505_),
    .B(_05506_),
    .C(_05678_),
    .X(_05726_));
 sky130_fd_sc_hd__o21ai_1 _16269_ (.A1(_05509_),
    .A2(_05675_),
    .B1(_05678_),
    .Y(_05727_));
 sky130_fd_sc_hd__a21boi_1 _16270_ (.A1(_05510_),
    .A2(_05676_),
    .B1_N(_05678_),
    .Y(_05728_));
 sky130_fd_sc_hd__o21ai_1 _16271_ (.A1(_05621_),
    .A2(_05660_),
    .B1(_05662_),
    .Y(_05729_));
 sky130_fd_sc_hd__a21o_1 _16272_ (.A1(_05625_),
    .A2(_05632_),
    .B1(_05630_),
    .X(_05730_));
 sky130_fd_sc_hd__a21oi_1 _16273_ (.A1(_05625_),
    .A2(_05632_),
    .B1(_05630_),
    .Y(_05732_));
 sky130_fd_sc_hd__and3_1 _16274_ (.A(_05841_),
    .B(net265),
    .C(net280),
    .X(_05733_));
 sky130_fd_sc_hd__nor2_1 _16275_ (.A(_03835_),
    .B(_04270_),
    .Y(_05734_));
 sky130_fd_sc_hd__a31o_1 _16276_ (.A1(_05841_),
    .A2(net265),
    .A3(net280),
    .B1(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__nand4_2 _16277_ (.A(_04037_),
    .B(_07242_),
    .C(net257),
    .D(net39),
    .Y(_05736_));
 sky130_fd_sc_hd__or3_1 _16278_ (.A(net39),
    .B(_04037_),
    .C(_03938_),
    .X(_05737_));
 sky130_fd_sc_hd__nor2_1 _16279_ (.A(_03916_),
    .B(_04218_),
    .Y(_05738_));
 sky130_fd_sc_hd__a31oi_4 _16280_ (.A1(_06486_),
    .A2(net261),
    .A3(_04215_),
    .B1(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__o311a_1 _16281_ (.A1(_03938_),
    .A2(_04037_),
    .A3(net39),
    .B1(_05739_),
    .C1(_05736_),
    .X(_05740_));
 sky130_fd_sc_hd__o221ai_4 _16282_ (.A1(_07263_),
    .A2(_03714_),
    .B1(_03737_),
    .B2(_03938_),
    .C1(_05739_),
    .Y(_05741_));
 sky130_fd_sc_hd__a21oi_1 _16283_ (.A1(_05736_),
    .A2(_05737_),
    .B1(_05739_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21o_1 _16284_ (.A1(_05736_),
    .A2(_05737_),
    .B1(_05739_),
    .X(_05744_));
 sky130_fd_sc_hd__nand3b_1 _16285_ (.A_N(_05735_),
    .B(_05741_),
    .C(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__o22ai_1 _16286_ (.A1(_05733_),
    .A2(_05734_),
    .B1(_05740_),
    .B2(_05743_),
    .Y(_05746_));
 sky130_fd_sc_hd__nor2_1 _16287_ (.A(_05735_),
    .B(_05743_),
    .Y(_05747_));
 sky130_fd_sc_hd__a21o_1 _16288_ (.A1(_05735_),
    .A2(_05741_),
    .B1(_05743_),
    .X(_05748_));
 sky130_fd_sc_hd__a31o_2 _16289_ (.A1(_05736_),
    .A2(_05737_),
    .A3(_05739_),
    .B1(_05747_),
    .X(_05749_));
 sky130_fd_sc_hd__o211ai_1 _16290_ (.A1(_05733_),
    .A2(_05734_),
    .B1(_05741_),
    .C1(_05744_),
    .Y(_05750_));
 sky130_fd_sc_hd__o21bai_1 _16291_ (.A1(_05740_),
    .A2(_05743_),
    .B1_N(_05735_),
    .Y(_05751_));
 sky130_fd_sc_hd__nand3_2 _16292_ (.A(_05730_),
    .B(_05750_),
    .C(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand3_2 _16293_ (.A(_05732_),
    .B(_05745_),
    .C(_05746_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2_1 _16294_ (.A(_05482_),
    .B(_05485_),
    .Y(_05755_));
 sky130_fd_sc_hd__a21oi_1 _16295_ (.A1(_05752_),
    .A2(_05754_),
    .B1(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__a21o_1 _16296_ (.A1(_05752_),
    .A2(_05754_),
    .B1(_05755_),
    .X(_05757_));
 sky130_fd_sc_hd__and3_1 _16297_ (.A(_05752_),
    .B(_05754_),
    .C(_05755_),
    .X(_05758_));
 sky130_fd_sc_hd__nand3_2 _16298_ (.A(_05752_),
    .B(_05754_),
    .C(_05755_),
    .Y(_05759_));
 sky130_fd_sc_hd__o221ai_4 _16299_ (.A1(_05211_),
    .A2(_05488_),
    .B1(_05756_),
    .B2(_05758_),
    .C1(_05491_),
    .Y(_05760_));
 sky130_fd_sc_hd__o211ai_4 _16300_ (.A1(_05489_),
    .A2(_05493_),
    .B1(_05757_),
    .C1(_05759_),
    .Y(_05761_));
 sky130_fd_sc_hd__and2b_4 _16301_ (.A_N(net47),
    .B(net48),
    .X(_05762_));
 sky130_fd_sc_hd__nand2b_4 _16302_ (.A_N(net47),
    .B(net48),
    .Y(_05763_));
 sky130_fd_sc_hd__and2b_4 _16303_ (.A_N(net48),
    .B(net47),
    .X(_05765_));
 sky130_fd_sc_hd__nand2b_4 _16304_ (.A_N(net48),
    .B(net47),
    .Y(_05766_));
 sky130_fd_sc_hd__a21oi_1 _16305_ (.A1(_05763_),
    .A2(_05766_),
    .B1(_03176_),
    .Y(_05767_));
 sky130_fd_sc_hd__o2bb2a_1 _16306_ (.A1_N(net12),
    .A2_N(_05464_),
    .B1(_05463_),
    .B2(_04528_),
    .X(_05768_));
 sky130_fd_sc_hd__a32o_1 _16307_ (.A1(net318),
    .A2(_04452_),
    .A3(net276),
    .B1(_05228_),
    .B2(net23),
    .X(_05769_));
 sky130_fd_sc_hd__nand2b_1 _16308_ (.A_N(_05768_),
    .B(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__a221o_1 _16309_ (.A1(_04539_),
    .A2(_05462_),
    .B1(_05464_),
    .B2(net12),
    .C1(_05769_),
    .X(_05771_));
 sky130_fd_sc_hd__o2111ai_1 _16310_ (.A1(net275),
    .A2(_05765_),
    .B1(_05771_),
    .C1(net1),
    .D1(_05770_),
    .Y(_05772_));
 sky130_fd_sc_hd__a21o_1 _16311_ (.A1(_05770_),
    .A2(_05771_),
    .B1(_05767_),
    .X(_05773_));
 sky130_fd_sc_hd__nand2_1 _16312_ (.A(_05772_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__a32o_1 _16313_ (.A1(_04985_),
    .A2(_04747_),
    .A3(net315),
    .B1(net26),
    .B2(_04988_),
    .X(_05776_));
 sky130_fd_sc_hd__or3b_1 _16314_ (.A(_03616_),
    .B(net43),
    .C_N(net42),
    .X(_05777_));
 sky130_fd_sc_hd__nand3_2 _16315_ (.A(net266),
    .B(net303),
    .C(net243),
    .Y(_05778_));
 sky130_fd_sc_hd__or3b_2 _16316_ (.A(_03725_),
    .B(net42),
    .C_N(net41),
    .X(_05779_));
 sky130_fd_sc_hd__o211ai_4 _16317_ (.A1(_04747_),
    .A2(_05436_),
    .B1(net279),
    .C1(_05414_),
    .Y(_05780_));
 sky130_fd_sc_hd__a22oi_4 _16318_ (.A1(_05777_),
    .A2(_05778_),
    .B1(_05779_),
    .B2(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__o2111a_1 _16319_ (.A1(_03616_),
    .A2(_04898_),
    .B1(_05778_),
    .C1(_05779_),
    .D1(_05780_),
    .X(_05782_));
 sky130_fd_sc_hd__o2111ai_4 _16320_ (.A1(_03616_),
    .A2(_04898_),
    .B1(_05778_),
    .C1(_05779_),
    .D1(_05780_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21ai_1 _16321_ (.A1(_05781_),
    .A2(_05782_),
    .B1(_05776_),
    .Y(_05784_));
 sky130_fd_sc_hd__or3_1 _16322_ (.A(_05776_),
    .B(_05781_),
    .C(_05782_),
    .X(_05785_));
 sky130_fd_sc_hd__a21boi_1 _16323_ (.A1(_05451_),
    .A2(_05456_),
    .B1_N(_05455_),
    .Y(_05787_));
 sky130_fd_sc_hd__a21oi_2 _16324_ (.A1(_05784_),
    .A2(_05785_),
    .B1(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__and3_1 _16325_ (.A(_05784_),
    .B(_05785_),
    .C(_05787_),
    .X(_05789_));
 sky130_fd_sc_hd__a31o_1 _16326_ (.A1(_05784_),
    .A2(_05785_),
    .A3(_05787_),
    .B1(_05774_),
    .X(_05790_));
 sky130_fd_sc_hd__o21ai_1 _16327_ (.A1(_05788_),
    .A2(_05789_),
    .B1(_05774_),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_1 _16328_ (.A1(_05788_),
    .A2(_05790_),
    .B1(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__o21a_1 _16329_ (.A1(_05788_),
    .A2(_05790_),
    .B1(_05791_),
    .X(_05793_));
 sky130_fd_sc_hd__a21o_1 _16330_ (.A1(_05760_),
    .A2(_05761_),
    .B1(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__o2111a_1 _16331_ (.A1(_05788_),
    .A2(_05790_),
    .B1(_05791_),
    .C1(_05761_),
    .D1(_05760_),
    .X(_05795_));
 sky130_fd_sc_hd__nand3_1 _16332_ (.A(_05760_),
    .B(_05792_),
    .C(_05761_),
    .Y(_05796_));
 sky130_fd_sc_hd__a21o_1 _16333_ (.A1(_05760_),
    .A2(_05761_),
    .B1(_05792_),
    .X(_05798_));
 sky130_fd_sc_hd__nand3b_4 _16334_ (.A_N(_05795_),
    .B(_05729_),
    .C(_05794_),
    .Y(_05799_));
 sky130_fd_sc_hd__o2111ai_4 _16335_ (.A1(_05621_),
    .A2(_05660_),
    .B1(_05662_),
    .C1(_05796_),
    .D1(_05798_),
    .Y(_05800_));
 sky130_fd_sc_hd__a21o_1 _16336_ (.A1(_05496_),
    .A2(_05473_),
    .B1(_05497_),
    .X(_05801_));
 sky130_fd_sc_hd__a21oi_2 _16337_ (.A1(_05799_),
    .A2(_05800_),
    .B1(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__a21o_1 _16338_ (.A1(_05799_),
    .A2(_05800_),
    .B1(_05801_),
    .X(_05803_));
 sky130_fd_sc_hd__and3_1 _16339_ (.A(_05799_),
    .B(_05800_),
    .C(_05801_),
    .X(_05804_));
 sky130_fd_sc_hd__nand3_4 _16340_ (.A(_05799_),
    .B(_05800_),
    .C(_05801_),
    .Y(_05805_));
 sky130_fd_sc_hd__nand2_1 _16341_ (.A(_05803_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21ai_1 _16342_ (.A1(_05663_),
    .A2(_05664_),
    .B1(_05619_),
    .Y(_05807_));
 sky130_fd_sc_hd__nand2_2 _16343_ (.A(_05620_),
    .B(_05807_),
    .Y(_05809_));
 sky130_fd_sc_hd__a32o_1 _16344_ (.A1(net235),
    .A2(net251),
    .A3(net252),
    .B1(_11793_),
    .B2(net4),
    .X(_05810_));
 sky130_fd_sc_hd__o211ai_4 _16345_ (.A1(net254),
    .A2(_00646_),
    .B1(net289),
    .C1(_00625_),
    .Y(_05811_));
 sky130_fd_sc_hd__or3b_2 _16346_ (.A(net34),
    .B(_04015_),
    .C_N(net64),
    .X(_05812_));
 sky130_fd_sc_hd__nor2_1 _16347_ (.A(_04026_),
    .B(_08283_),
    .Y(_05813_));
 sky130_fd_sc_hd__or3b_1 _16348_ (.A(net64),
    .B(_04026_),
    .C_N(net63),
    .X(_05814_));
 sky130_fd_sc_hd__o311a_1 _16349_ (.A1(net261),
    .A2(_11387_),
    .A3(_02442_),
    .B1(net291),
    .C1(_02421_),
    .X(_05815_));
 sky130_fd_sc_hd__o211ai_4 _16350_ (.A1(net254),
    .A2(_02442_),
    .B1(net291),
    .C1(_02421_),
    .Y(_05816_));
 sky130_fd_sc_hd__o211ai_2 _16351_ (.A1(_04015_),
    .A2(_10346_),
    .B1(_05811_),
    .C1(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__o2111ai_4 _16352_ (.A1(_04026_),
    .A2(_08283_),
    .B1(_05811_),
    .C1(_05812_),
    .D1(_05816_),
    .Y(_05818_));
 sky130_fd_sc_hd__a22oi_1 _16353_ (.A1(_05811_),
    .A2(_05812_),
    .B1(_05814_),
    .B2(_05816_),
    .Y(_05820_));
 sky130_fd_sc_hd__o2bb2ai_2 _16354_ (.A1_N(_05811_),
    .A2_N(_05812_),
    .B1(_05813_),
    .B2(_05815_),
    .Y(_05821_));
 sky130_fd_sc_hd__o211a_1 _16355_ (.A1(_05813_),
    .A2(_05817_),
    .B1(_05821_),
    .C1(_05810_),
    .X(_05822_));
 sky130_fd_sc_hd__o211ai_2 _16356_ (.A1(_05813_),
    .A2(_05817_),
    .B1(_05821_),
    .C1(_05810_),
    .Y(_05823_));
 sky130_fd_sc_hd__a21oi_1 _16357_ (.A1(_05818_),
    .A2(_05821_),
    .B1(_05810_),
    .Y(_05824_));
 sky130_fd_sc_hd__a21o_1 _16358_ (.A1(_05818_),
    .A2(_05821_),
    .B1(_05810_),
    .X(_05825_));
 sky130_fd_sc_hd__o22ai_4 _16359_ (.A1(_05643_),
    .A2(_05650_),
    .B1(_05822_),
    .B2(_05824_),
    .Y(_05826_));
 sky130_fd_sc_hd__o2111ai_4 _16360_ (.A1(_05646_),
    .A2(_05639_),
    .B1(_05645_),
    .C1(_05823_),
    .D1(_05825_),
    .Y(_05827_));
 sky130_fd_sc_hd__inv_2 _16361_ (.A(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__o32a_1 _16362_ (.A1(_02869_),
    .A2(_08689_),
    .A3(_08667_),
    .B1(_03949_),
    .B2(_02891_),
    .X(_05829_));
 sky130_fd_sc_hd__a32o_1 _16363_ (.A1(net256),
    .A2(_08700_),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net32),
    .X(_05831_));
 sky130_fd_sc_hd__o211ai_2 _16364_ (.A1(net261),
    .A2(_09665_),
    .B1(_01293_),
    .C1(_09698_),
    .Y(_05832_));
 sky130_fd_sc_hd__or3b_2 _16365_ (.A(_03960_),
    .B(net37),
    .C_N(net36),
    .X(_05833_));
 sky130_fd_sc_hd__o2111ai_4 _16366_ (.A1(net261),
    .A2(_11387_),
    .B1(net36),
    .C1(_11354_),
    .D1(_03993_),
    .Y(_05834_));
 sky130_fd_sc_hd__or3_2 _16367_ (.A(net36),
    .B(_03993_),
    .C(_03982_),
    .X(_05835_));
 sky130_fd_sc_hd__a22oi_4 _16368_ (.A1(_05832_),
    .A2(_05833_),
    .B1(_05834_),
    .B2(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__and4_1 _16369_ (.A(_05832_),
    .B(_05833_),
    .C(_05834_),
    .D(_05835_),
    .X(_05837_));
 sky130_fd_sc_hd__nand4_1 _16370_ (.A(_05832_),
    .B(_05833_),
    .C(_05834_),
    .D(_05835_),
    .Y(_05838_));
 sky130_fd_sc_hd__o21a_1 _16371_ (.A1(_05836_),
    .A2(_05837_),
    .B1(_05829_),
    .X(_05839_));
 sky130_fd_sc_hd__nor3_1 _16372_ (.A(_05829_),
    .B(_05836_),
    .C(_05837_),
    .Y(_05840_));
 sky130_fd_sc_hd__o21a_1 _16373_ (.A1(_05836_),
    .A2(_05837_),
    .B1(_05831_),
    .X(_05842_));
 sky130_fd_sc_hd__nor3_1 _16374_ (.A(_05831_),
    .B(_05836_),
    .C(_05837_),
    .Y(_05843_));
 sky130_fd_sc_hd__o2bb2ai_1 _16375_ (.A1_N(_05826_),
    .A2_N(_05827_),
    .B1(_05839_),
    .B2(_05840_),
    .Y(_05844_));
 sky130_fd_sc_hd__o211a_2 _16376_ (.A1(_05842_),
    .A2(_05843_),
    .B1(_05826_),
    .C1(_05827_),
    .X(_05845_));
 sky130_fd_sc_hd__o211ai_4 _16377_ (.A1(_05842_),
    .A2(_05843_),
    .B1(_05826_),
    .C1(_05827_),
    .Y(_05846_));
 sky130_fd_sc_hd__o21ai_2 _16378_ (.A1(_05514_),
    .A2(_05532_),
    .B1(_05536_),
    .Y(_05847_));
 sky130_fd_sc_hd__a21o_2 _16379_ (.A1(_05844_),
    .A2(_05846_),
    .B1(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__nand2_1 _16380_ (.A(_05847_),
    .B(_05844_),
    .Y(_05849_));
 sky130_fd_sc_hd__nand3_2 _16381_ (.A(_05847_),
    .B(_05846_),
    .C(_05844_),
    .Y(_05850_));
 sky130_fd_sc_hd__a21o_2 _16382_ (.A1(_05636_),
    .A2(_05657_),
    .B1(_05653_),
    .X(_05851_));
 sky130_fd_sc_hd__a21oi_2 _16383_ (.A1(_05848_),
    .A2(_05850_),
    .B1(_05851_),
    .Y(_05853_));
 sky130_fd_sc_hd__a21o_1 _16384_ (.A1(_05848_),
    .A2(_05850_),
    .B1(_05851_),
    .X(_05854_));
 sky130_fd_sc_hd__o211ai_4 _16385_ (.A1(_05845_),
    .A2(_05849_),
    .B1(_05851_),
    .C1(_05848_),
    .Y(_05855_));
 sky130_fd_sc_hd__inv_2 _16386_ (.A(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _16387_ (.A(_05854_),
    .B(_05855_),
    .Y(_05857_));
 sky130_fd_sc_hd__a31o_1 _16388_ (.A1(_05541_),
    .A2(_05542_),
    .A3(_05607_),
    .B1(_05610_),
    .X(_05858_));
 sky130_fd_sc_hd__a22oi_2 _16389_ (.A1(_05609_),
    .A2(_05606_),
    .B1(_05543_),
    .B2(_05607_),
    .Y(_05859_));
 sky130_fd_sc_hd__and3_1 _16390_ (.A(_03952_),
    .B(net232),
    .C(_07658_),
    .X(_05860_));
 sky130_fd_sc_hd__nor2_1 _16391_ (.A(_04048_),
    .B(_07691_),
    .Y(_05861_));
 sky130_fd_sc_hd__a31o_1 _16392_ (.A1(_03952_),
    .A2(net232),
    .A3(_07658_),
    .B1(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__nand3_2 _16393_ (.A(net224),
    .B(net299),
    .C(net188),
    .Y(_05864_));
 sky130_fd_sc_hd__or3b_1 _16394_ (.A(net61),
    .B(_04069_),
    .C_N(net60),
    .X(_05865_));
 sky130_fd_sc_hd__and3_1 _16395_ (.A(_03927_),
    .B(net8),
    .C(net61),
    .X(_05866_));
 sky130_fd_sc_hd__and3_1 _16396_ (.A(_04132_),
    .B(net292),
    .C(net230),
    .X(_05867_));
 sky130_fd_sc_hd__a31oi_2 _16397_ (.A1(_04132_),
    .A2(net292),
    .A3(net230),
    .B1(_05866_),
    .Y(_05868_));
 sky130_fd_sc_hd__o211ai_4 _16398_ (.A1(_04069_),
    .A2(net298),
    .B1(_05864_),
    .C1(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__o2bb2ai_4 _16399_ (.A1_N(_05864_),
    .A2_N(_05865_),
    .B1(_05866_),
    .B2(_05867_),
    .Y(_05870_));
 sky130_fd_sc_hd__o211a_1 _16400_ (.A1(_05860_),
    .A2(_05861_),
    .B1(_05869_),
    .C1(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__o211ai_4 _16401_ (.A1(_05860_),
    .A2(_05861_),
    .B1(_05869_),
    .C1(_05870_),
    .Y(_05872_));
 sky130_fd_sc_hd__a21oi_1 _16402_ (.A1(_05869_),
    .A2(_05870_),
    .B1(_05862_),
    .Y(_05873_));
 sky130_fd_sc_hd__a21o_1 _16403_ (.A1(_05869_),
    .A2(_05870_),
    .B1(_05862_),
    .X(_05875_));
 sky130_fd_sc_hd__a21oi_1 _16404_ (.A1(_05872_),
    .A2(_05875_),
    .B1(_05591_),
    .Y(_05876_));
 sky130_fd_sc_hd__o221ai_4 _16405_ (.A1(_05580_),
    .A2(_05587_),
    .B1(_05871_),
    .B2(_05873_),
    .C1(_05586_),
    .Y(_05877_));
 sky130_fd_sc_hd__nand3_4 _16406_ (.A(_05591_),
    .B(_05872_),
    .C(_05875_),
    .Y(_05878_));
 sky130_fd_sc_hd__a21bo_1 _16407_ (.A1(_05877_),
    .A2(_05878_),
    .B1_N(_05529_),
    .X(_05879_));
 sky130_fd_sc_hd__nand3b_2 _16408_ (.A_N(_05529_),
    .B(_05877_),
    .C(_05878_),
    .Y(_05880_));
 sky130_fd_sc_hd__a21oi_1 _16409_ (.A1(_05877_),
    .A2(_05878_),
    .B1(_05529_),
    .Y(_05881_));
 sky130_fd_sc_hd__a21o_1 _16410_ (.A1(_05877_),
    .A2(_05878_),
    .B1(_05529_),
    .X(_05882_));
 sky130_fd_sc_hd__and3_1 _16411_ (.A(_05529_),
    .B(_05877_),
    .C(_05878_),
    .X(_05883_));
 sky130_fd_sc_hd__nand3_1 _16412_ (.A(_05529_),
    .B(_05877_),
    .C(_05878_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand2_1 _16413_ (.A(_05879_),
    .B(_05880_),
    .Y(_05886_));
 sky130_fd_sc_hd__nor2_1 _16414_ (.A(_04080_),
    .B(_05260_),
    .Y(_05887_));
 sky130_fd_sc_hd__o311a_1 _16415_ (.A1(net7),
    .A2(net249),
    .A3(_04557_),
    .B1(_05227_),
    .C1(net219),
    .X(_05888_));
 sky130_fd_sc_hd__o32a_1 _16416_ (.A1(_04558_),
    .A2(_05238_),
    .A3(_04554_),
    .B1(_05260_),
    .B2(_04080_),
    .X(_05889_));
 sky130_fd_sc_hd__a31o_1 _16417_ (.A1(net219),
    .A2(_04559_),
    .A3(_05227_),
    .B1(_05887_),
    .X(_05890_));
 sky130_fd_sc_hd__nand3_2 _16418_ (.A(net212),
    .B(net183),
    .C(net317),
    .Y(_05891_));
 sky130_fd_sc_hd__nor2_1 _16419_ (.A(_04113_),
    .B(net316),
    .Y(_05892_));
 sky130_fd_sc_hd__or3b_2 _16420_ (.A(net58),
    .B(_04113_),
    .C_N(net55),
    .X(_05893_));
 sky130_fd_sc_hd__a31oi_1 _16421_ (.A1(net212),
    .A2(net183),
    .A3(net317),
    .B1(_05892_),
    .Y(_05894_));
 sky130_fd_sc_hd__a31o_1 _16422_ (.A1(net212),
    .A2(net183),
    .A3(net317),
    .B1(_05892_),
    .X(_05895_));
 sky130_fd_sc_hd__or3b_2 _16423_ (.A(net59),
    .B(_04091_),
    .C_N(net58),
    .X(_05897_));
 sky130_fd_sc_hd__nand3_2 _16424_ (.A(net215),
    .B(net305),
    .C(net185),
    .Y(_05898_));
 sky130_fd_sc_hd__a32oi_1 _16425_ (.A1(_04790_),
    .A2(net305),
    .A3(net185),
    .B1(_04911_),
    .B2(net11),
    .Y(_05899_));
 sky130_fd_sc_hd__nand2_1 _16426_ (.A(_05897_),
    .B(_05898_),
    .Y(_05900_));
 sky130_fd_sc_hd__nand4_4 _16427_ (.A(_05891_),
    .B(_05893_),
    .C(_05897_),
    .D(_05898_),
    .Y(_05901_));
 sky130_fd_sc_hd__nor2_1 _16428_ (.A(_05890_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__a22oi_2 _16429_ (.A1(_05891_),
    .A2(_05893_),
    .B1(_05897_),
    .B2(_05898_),
    .Y(_05903_));
 sky130_fd_sc_hd__a22o_1 _16430_ (.A1(_05891_),
    .A2(_05893_),
    .B1(_05897_),
    .B2(_05898_),
    .X(_05904_));
 sky130_fd_sc_hd__o21ai_1 _16431_ (.A1(_05894_),
    .A2(_05899_),
    .B1(_05889_),
    .Y(_05905_));
 sky130_fd_sc_hd__a21o_1 _16432_ (.A1(_05890_),
    .A2(_05901_),
    .B1(_05903_),
    .X(_05906_));
 sky130_fd_sc_hd__a21oi_4 _16433_ (.A1(_05890_),
    .A2(_05901_),
    .B1(_05903_),
    .Y(_05908_));
 sky130_fd_sc_hd__o211ai_1 _16434_ (.A1(_05887_),
    .A2(_05888_),
    .B1(_05895_),
    .C1(_05900_),
    .Y(_05909_));
 sky130_fd_sc_hd__a21oi_2 _16435_ (.A1(_05901_),
    .A2(_05904_),
    .B1(_05889_),
    .Y(_05910_));
 sky130_fd_sc_hd__and3_1 _16436_ (.A(_05904_),
    .B(_05889_),
    .C(_05901_),
    .X(_05911_));
 sky130_fd_sc_hd__a211o_1 _16437_ (.A1(_05901_),
    .A2(_05904_),
    .B1(_05887_),
    .C1(_05888_),
    .X(_05912_));
 sky130_fd_sc_hd__o211ai_2 _16438_ (.A1(_05887_),
    .A2(_05888_),
    .B1(_05901_),
    .C1(_05904_),
    .Y(_05913_));
 sky130_fd_sc_hd__a31oi_1 _16439_ (.A1(_05901_),
    .A2(_05905_),
    .A3(_05909_),
    .B1(_05902_),
    .Y(_05914_));
 sky130_fd_sc_hd__a31o_1 _16440_ (.A1(_05901_),
    .A2(_05905_),
    .A3(_05909_),
    .B1(_05902_),
    .X(_05915_));
 sky130_fd_sc_hd__nor2_2 _16441_ (.A(_04135_),
    .B(_04375_),
    .Y(_05916_));
 sky130_fd_sc_hd__and3_2 _16442_ (.A(net181),
    .B(net180),
    .C(_04342_),
    .X(_05917_));
 sky130_fd_sc_hd__a31oi_4 _16443_ (.A1(net181),
    .A2(net180),
    .A3(_04342_),
    .B1(_05916_),
    .Y(_05919_));
 sky130_fd_sc_hd__a31o_1 _16444_ (.A1(net181),
    .A2(net180),
    .A3(_04342_),
    .B1(_05916_),
    .X(_05920_));
 sky130_fd_sc_hd__o211ai_4 _16445_ (.A1(net185),
    .A2(_05551_),
    .B1(_04484_),
    .C1(_05549_),
    .Y(_05921_));
 sky130_fd_sc_hd__nor2_1 _16446_ (.A(_04146_),
    .B(_04331_),
    .Y(_05922_));
 sky130_fd_sc_hd__or3_1 _16447_ (.A(net44),
    .B(_04146_),
    .C(_03286_),
    .X(_05923_));
 sky130_fd_sc_hd__nor4_4 _16448_ (.A(net13),
    .B(net14),
    .C(net15),
    .D(net16),
    .Y(_05924_));
 sky130_fd_sc_hd__nand3_4 _16449_ (.A(_04406_),
    .B(_04785_),
    .C(_04157_),
    .Y(_05925_));
 sky130_fd_sc_hd__nor2_8 _16450_ (.A(_05551_),
    .B(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__nand2_8 _16451_ (.A(net278),
    .B(_05924_),
    .Y(_05927_));
 sky130_fd_sc_hd__nand4_4 _16452_ (.A(net311),
    .B(net293),
    .C(net278),
    .D(_05924_),
    .Y(_05928_));
 sky130_fd_sc_hd__nor3_4 _16453_ (.A(net262),
    .B(net244),
    .C(_05927_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand3_4 _16454_ (.A(_06519_),
    .B(_03955_),
    .C(_05926_),
    .Y(_05931_));
 sky130_fd_sc_hd__a41oi_4 _16455_ (.A1(_06519_),
    .A2(_03955_),
    .A3(net277),
    .A4(_05550_),
    .B1(_04157_),
    .Y(_05932_));
 sky130_fd_sc_hd__a41o_4 _16456_ (.A1(_06519_),
    .A2(_03955_),
    .A3(net277),
    .A4(_05550_),
    .B1(_04157_),
    .X(_05933_));
 sky130_fd_sc_hd__o32a_1 _16457_ (.A1(net7),
    .A2(net248),
    .A3(_05927_),
    .B1(_04157_),
    .B2(net207),
    .X(_05934_));
 sky130_fd_sc_hd__o2bb2ai_4 _16458_ (.A1_N(net16),
    .A2_N(_05553_),
    .B1(_05927_),
    .B2(net233),
    .Y(_05935_));
 sky130_fd_sc_hd__o211ai_4 _16459_ (.A1(net232),
    .A2(_05927_),
    .B1(net33),
    .C1(_05933_),
    .Y(_05936_));
 sky130_fd_sc_hd__and4_1 _16460_ (.A(_05933_),
    .B(_05922_),
    .C(net33),
    .D(net175),
    .X(_05937_));
 sky130_fd_sc_hd__nand4_4 _16461_ (.A(_05933_),
    .B(_05922_),
    .C(net33),
    .D(net175),
    .Y(_05938_));
 sky130_fd_sc_hd__o311a_1 _16462_ (.A1(_03286_),
    .A2(net44),
    .A3(_04146_),
    .B1(_05921_),
    .C1(_05936_),
    .X(_05939_));
 sky130_fd_sc_hd__o221ai_4 _16463_ (.A1(_04146_),
    .A2(_04331_),
    .B1(net155),
    .B2(_03286_),
    .C1(_05921_),
    .Y(_05941_));
 sky130_fd_sc_hd__o21bai_2 _16464_ (.A1(_05937_),
    .A2(_05939_),
    .B1_N(_05920_),
    .Y(_05942_));
 sky130_fd_sc_hd__o211ai_4 _16465_ (.A1(_05916_),
    .A2(_05917_),
    .B1(_05938_),
    .C1(_05941_),
    .Y(_05943_));
 sky130_fd_sc_hd__nand3_2 _16466_ (.A(_05941_),
    .B(_05919_),
    .C(_05938_),
    .Y(_05944_));
 sky130_fd_sc_hd__o22ai_4 _16467_ (.A1(_05916_),
    .A2(_05917_),
    .B1(_05937_),
    .B2(_05939_),
    .Y(_05945_));
 sky130_fd_sc_hd__o31a_1 _16468_ (.A1(_05559_),
    .A2(_05563_),
    .A3(_05564_),
    .B1(_05561_),
    .X(_05946_));
 sky130_fd_sc_hd__a21oi_4 _16469_ (.A1(_05561_),
    .A2(_05566_),
    .B1(_05559_),
    .Y(_05947_));
 sky130_fd_sc_hd__and3_1 _16470_ (.A(_05944_),
    .B(_05945_),
    .C(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__nand3_4 _16471_ (.A(_05944_),
    .B(_05945_),
    .C(_05947_),
    .Y(_05949_));
 sky130_fd_sc_hd__nand3_4 _16472_ (.A(_05942_),
    .B(_05943_),
    .C(_05946_),
    .Y(_05950_));
 sky130_fd_sc_hd__a31oi_2 _16473_ (.A1(_05942_),
    .A2(_05943_),
    .A3(_05946_),
    .B1(_05914_),
    .Y(_05952_));
 sky130_fd_sc_hd__a32oi_4 _16474_ (.A1(_05944_),
    .A2(_05945_),
    .A3(_05947_),
    .B1(_05950_),
    .B2(_05915_),
    .Y(_05953_));
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(_05949_),
    .B(_05950_),
    .Y(_05954_));
 sky130_fd_sc_hd__a22oi_2 _16476_ (.A1(_05912_),
    .A2(_05913_),
    .B1(_05949_),
    .B2(_05950_),
    .Y(_05955_));
 sky130_fd_sc_hd__a22o_1 _16477_ (.A1(_05912_),
    .A2(_05913_),
    .B1(_05949_),
    .B2(_05950_),
    .X(_05956_));
 sky130_fd_sc_hd__o21ai_1 _16478_ (.A1(_05910_),
    .A2(_05911_),
    .B1(_05950_),
    .Y(_05957_));
 sky130_fd_sc_hd__o211a_1 _16479_ (.A1(_05910_),
    .A2(_05911_),
    .B1(_05949_),
    .C1(_05950_),
    .X(_05958_));
 sky130_fd_sc_hd__o211ai_4 _16480_ (.A1(_05910_),
    .A2(_05911_),
    .B1(_05949_),
    .C1(_05950_),
    .Y(_05959_));
 sky130_fd_sc_hd__o2bb2ai_2 _16481_ (.A1_N(_05915_),
    .A2_N(_05954_),
    .B1(_05957_),
    .B2(_05948_),
    .Y(_05960_));
 sky130_fd_sc_hd__a21oi_1 _16482_ (.A1(_05956_),
    .A2(_05959_),
    .B1(_05603_),
    .Y(_05961_));
 sky130_fd_sc_hd__o22ai_4 _16483_ (.A1(_05577_),
    .A2(_05601_),
    .B1(_05955_),
    .B2(_05958_),
    .Y(_05963_));
 sky130_fd_sc_hd__and3_1 _16484_ (.A(_05956_),
    .B(_05959_),
    .C(_05603_),
    .X(_05964_));
 sky130_fd_sc_hd__nand3_4 _16485_ (.A(_05956_),
    .B(_05959_),
    .C(_05603_),
    .Y(_05965_));
 sky130_fd_sc_hd__a22oi_4 _16486_ (.A1(_05882_),
    .A2(_05884_),
    .B1(_05960_),
    .B2(_05604_),
    .Y(_05966_));
 sky130_fd_sc_hd__o32a_2 _16487_ (.A1(_05577_),
    .A2(_05601_),
    .A3(_05960_),
    .B1(_05886_),
    .B2(_05961_),
    .X(_05967_));
 sky130_fd_sc_hd__o21ai_1 _16488_ (.A1(_05886_),
    .A2(_05961_),
    .B1(_05965_),
    .Y(_05968_));
 sky130_fd_sc_hd__o211a_2 _16489_ (.A1(_05881_),
    .A2(_05883_),
    .B1(_05963_),
    .C1(_05965_),
    .X(_05969_));
 sky130_fd_sc_hd__o211ai_2 _16490_ (.A1(_05881_),
    .A2(_05883_),
    .B1(_05963_),
    .C1(_05965_),
    .Y(_05970_));
 sky130_fd_sc_hd__a22oi_4 _16491_ (.A1(_05879_),
    .A2(_05880_),
    .B1(_05963_),
    .B2(_05965_),
    .Y(_05971_));
 sky130_fd_sc_hd__a22o_1 _16492_ (.A1(_05879_),
    .A2(_05880_),
    .B1(_05963_),
    .B2(_05965_),
    .X(_05972_));
 sky130_fd_sc_hd__nand2_2 _16493_ (.A(_05972_),
    .B(_05858_),
    .Y(_05974_));
 sky130_fd_sc_hd__a211oi_4 _16494_ (.A1(_05966_),
    .A2(_05965_),
    .B1(_05859_),
    .C1(_05971_),
    .Y(_05975_));
 sky130_fd_sc_hd__nand3_1 _16495_ (.A(_05972_),
    .B(_05858_),
    .C(_05970_),
    .Y(_05976_));
 sky130_fd_sc_hd__a2bb2oi_4 _16496_ (.A1_N(_05608_),
    .A2_N(_05614_),
    .B1(_05970_),
    .B2(_05972_),
    .Y(_05977_));
 sky130_fd_sc_hd__o22ai_4 _16497_ (.A1(_05608_),
    .A2(_05614_),
    .B1(_05969_),
    .B2(_05971_),
    .Y(_05978_));
 sky130_fd_sc_hd__o221ai_4 _16498_ (.A1(_05853_),
    .A2(_05856_),
    .B1(_05969_),
    .B2(_05974_),
    .C1(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21bai_4 _16499_ (.A1(_05975_),
    .A2(_05977_),
    .B1_N(_05857_),
    .Y(_05980_));
 sky130_fd_sc_hd__nand3b_2 _16500_ (.A_N(_05857_),
    .B(_05976_),
    .C(_05978_),
    .Y(_05981_));
 sky130_fd_sc_hd__o22ai_4 _16501_ (.A1(_05853_),
    .A2(_05856_),
    .B1(_05975_),
    .B2(_05977_),
    .Y(_05982_));
 sky130_fd_sc_hd__o211a_1 _16502_ (.A1(_05618_),
    .A2(_05669_),
    .B1(_05981_),
    .C1(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__o211ai_4 _16503_ (.A1(_05618_),
    .A2(_05669_),
    .B1(_05981_),
    .C1(_05982_),
    .Y(_05985_));
 sky130_fd_sc_hd__nand3_4 _16504_ (.A(_05980_),
    .B(_05809_),
    .C(_05979_),
    .Y(_05986_));
 sky130_fd_sc_hd__a31oi_4 _16505_ (.A1(_05980_),
    .A2(_05809_),
    .A3(_05979_),
    .B1(_05806_),
    .Y(_05987_));
 sky130_fd_sc_hd__nand2_1 _16506_ (.A(_05987_),
    .B(_05985_),
    .Y(_05988_));
 sky130_fd_sc_hd__inv_2 _16507_ (.A(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__a2bb2oi_1 _16508_ (.A1_N(_05802_),
    .A2_N(_05804_),
    .B1(_05985_),
    .B2(_05986_),
    .Y(_05990_));
 sky130_fd_sc_hd__a22o_1 _16509_ (.A1(_05803_),
    .A2(_05805_),
    .B1(_05985_),
    .B2(_05986_),
    .X(_05991_));
 sky130_fd_sc_hd__o211ai_2 _16510_ (.A1(_05802_),
    .A2(_05804_),
    .B1(_05985_),
    .C1(_05986_),
    .Y(_05992_));
 sky130_fd_sc_hd__a21o_1 _16511_ (.A1(_05985_),
    .A2(_05986_),
    .B1(_05806_),
    .X(_05993_));
 sky130_fd_sc_hd__nand2_1 _16512_ (.A(_05991_),
    .B(_05727_),
    .Y(_05994_));
 sky130_fd_sc_hd__a211oi_2 _16513_ (.A1(_05985_),
    .A2(_05987_),
    .B1(_05728_),
    .C1(_05990_),
    .Y(_05996_));
 sky130_fd_sc_hd__nand3_1 _16514_ (.A(_05991_),
    .B(_05727_),
    .C(_05988_),
    .Y(_05997_));
 sky130_fd_sc_hd__a2bb2oi_1 _16515_ (.A1_N(_05675_),
    .A2_N(_05726_),
    .B1(_05988_),
    .B2(_05991_),
    .Y(_05998_));
 sky130_fd_sc_hd__o2111ai_4 _16516_ (.A1(_05509_),
    .A2(_05675_),
    .B1(_05678_),
    .C1(_05992_),
    .D1(_05993_),
    .Y(_05999_));
 sky130_fd_sc_hd__o211ai_1 _16517_ (.A1(_05723_),
    .A2(_05724_),
    .B1(_05997_),
    .C1(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__o22ai_1 _16518_ (.A1(_05719_),
    .A2(_05722_),
    .B1(_05996_),
    .B2(_05998_),
    .Y(_06001_));
 sky130_fd_sc_hd__o22ai_2 _16519_ (.A1(_05723_),
    .A2(_05724_),
    .B1(_05996_),
    .B2(_05998_),
    .Y(_06002_));
 sky130_fd_sc_hd__o211ai_2 _16520_ (.A1(_05719_),
    .A2(_05722_),
    .B1(_05997_),
    .C1(_05999_),
    .Y(_06003_));
 sky130_fd_sc_hd__a21oi_1 _16521_ (.A1(_06002_),
    .A2(_06003_),
    .B1(_05714_),
    .Y(_06004_));
 sky130_fd_sc_hd__nand3b_1 _16522_ (.A_N(_05714_),
    .B(_06000_),
    .C(_06001_),
    .Y(_06005_));
 sky130_fd_sc_hd__a22oi_1 _16523_ (.A1(_05684_),
    .A2(_05713_),
    .B1(_06000_),
    .B2(_06001_),
    .Y(_06007_));
 sky130_fd_sc_hd__nand3_2 _16524_ (.A(_05714_),
    .B(_06002_),
    .C(_06003_),
    .Y(_06008_));
 sky130_fd_sc_hd__a21o_1 _16525_ (.A1(_06005_),
    .A2(_06008_),
    .B1(_05689_),
    .X(_06009_));
 sky130_fd_sc_hd__o211ai_2 _16526_ (.A1(_05685_),
    .A2(_05686_),
    .B1(_06005_),
    .C1(_06008_),
    .Y(_06010_));
 sky130_fd_sc_hd__o22ai_1 _16527_ (.A1(_05685_),
    .A2(_05686_),
    .B1(_06004_),
    .B2(_06007_),
    .Y(_06011_));
 sky130_fd_sc_hd__nand3_1 _16528_ (.A(_06005_),
    .B(_06008_),
    .C(_05687_),
    .Y(_06012_));
 sky130_fd_sc_hd__a21bo_1 _16529_ (.A1(_05422_),
    .A2(_05698_),
    .B1_N(_05700_),
    .X(_06013_));
 sky130_fd_sc_hd__a21boi_1 _16530_ (.A1(_05698_),
    .A2(_05422_),
    .B1_N(_05700_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand3_1 _16531_ (.A(_06009_),
    .B(_06010_),
    .C(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__a21oi_2 _16532_ (.A1(_06009_),
    .A2(_06010_),
    .B1(_06014_),
    .Y(_06016_));
 sky130_fd_sc_hd__nand3_1 _16533_ (.A(_06011_),
    .B(_06012_),
    .C(_06013_),
    .Y(_06018_));
 sky130_fd_sc_hd__a32o_2 _16534_ (.A1(_05432_),
    .A2(_05701_),
    .A3(_05704_),
    .B1(_06015_),
    .B2(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__nand2_1 _16535_ (.A(_05707_),
    .B(_06015_),
    .Y(_06020_));
 sky130_fd_sc_hd__a22oi_1 _16536_ (.A1(_05440_),
    .A2(_05708_),
    .B1(_05447_),
    .B2(_05711_),
    .Y(_06021_));
 sky130_fd_sc_hd__a21oi_1 _16537_ (.A1(_06019_),
    .A2(_06020_),
    .B1(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__and3_1 _16538_ (.A(_06019_),
    .B(_06020_),
    .C(_06021_),
    .X(_06023_));
 sky130_fd_sc_hd__nor2_1 _16539_ (.A(_06022_),
    .B(_06023_),
    .Y(net80));
 sky130_fd_sc_hd__o2bb2ai_2 _16540_ (.A1_N(_05725_),
    .A2_N(_05999_),
    .B1(_05994_),
    .B2(_05989_),
    .Y(_06024_));
 sky130_fd_sc_hd__a21oi_2 _16541_ (.A1(_05999_),
    .A2(_05725_),
    .B1(_05996_),
    .Y(_06025_));
 sky130_fd_sc_hd__and2b_4 _16542_ (.A_N(net48),
    .B(net49),
    .X(_06026_));
 sky130_fd_sc_hd__nand2b_4 _16543_ (.A_N(net48),
    .B(net49),
    .Y(_06028_));
 sky130_fd_sc_hd__and2b_4 _16544_ (.A_N(net49),
    .B(net48),
    .X(_06029_));
 sky130_fd_sc_hd__nand2b_4 _16545_ (.A_N(net49),
    .B(net48),
    .Y(_06030_));
 sky130_fd_sc_hd__a21oi_1 _16546_ (.A1(_06028_),
    .A2(_06030_),
    .B1(_03176_),
    .Y(_06031_));
 sky130_fd_sc_hd__a21bo_1 _16547_ (.A1(_05767_),
    .A2(_05771_),
    .B1_N(_05770_),
    .X(_06032_));
 sky130_fd_sc_hd__o211a_1 _16548_ (.A1(_06026_),
    .A2(_06029_),
    .B1(net1),
    .C1(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__nor2_1 _16549_ (.A(_06031_),
    .B(_06032_),
    .Y(_06034_));
 sky130_fd_sc_hd__or2_2 _16550_ (.A(_06033_),
    .B(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__o21ba_1 _16551_ (.A1(_05774_),
    .A2(_05789_),
    .B1_N(_05788_),
    .X(_06036_));
 sky130_fd_sc_hd__nor2_2 _16552_ (.A(_06035_),
    .B(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__and3b_2 _16553_ (.A_N(_05788_),
    .B(_05790_),
    .C(_06035_),
    .X(_06039_));
 sky130_fd_sc_hd__or2_1 _16554_ (.A(_06037_),
    .B(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__o21ai_1 _16555_ (.A1(_06037_),
    .A2(_06039_),
    .B1(_05716_),
    .Y(_06041_));
 sky130_fd_sc_hd__o41ai_4 _16556_ (.A1(_05461_),
    .A2(_05469_),
    .A3(_06037_),
    .A4(_06039_),
    .B1(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__a21oi_4 _16557_ (.A1(_05799_),
    .A2(_05805_),
    .B1(_06042_),
    .Y(_06043_));
 sky130_fd_sc_hd__and3_1 _16558_ (.A(_05799_),
    .B(_05805_),
    .C(_06042_),
    .X(_06044_));
 sky130_fd_sc_hd__and3b_1 _16559_ (.A_N(_06042_),
    .B(_05805_),
    .C(_05799_),
    .X(_06045_));
 sky130_fd_sc_hd__a21boi_2 _16560_ (.A1(_05799_),
    .A2(_05805_),
    .B1_N(_06042_),
    .Y(_06046_));
 sky130_fd_sc_hd__nor2_1 _16561_ (.A(_06043_),
    .B(_06044_),
    .Y(_06047_));
 sky130_fd_sc_hd__nor2_1 _16562_ (.A(_06045_),
    .B(_06046_),
    .Y(_06048_));
 sky130_fd_sc_hd__o21ai_4 _16563_ (.A1(_05802_),
    .A2(_05804_),
    .B1(_05985_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_1 _16564_ (.A(_05986_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__a22o_1 _16565_ (.A1(net12),
    .A2(_05765_),
    .B1(_04539_),
    .B2(net275),
    .X(_06052_));
 sky130_fd_sc_hd__a32oi_2 _16566_ (.A1(net318),
    .A2(_04452_),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net23),
    .Y(_06053_));
 sky130_fd_sc_hd__and3_1 _16567_ (.A(net313),
    .B(_04747_),
    .C(net276),
    .X(_06054_));
 sky130_fd_sc_hd__and3b_1 _16568_ (.A_N(net46),
    .B(net45),
    .C(net26),
    .X(_06055_));
 sky130_fd_sc_hd__a31oi_1 _16569_ (.A1(net313),
    .A2(_04747_),
    .A3(net276),
    .B1(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__nor2_1 _16570_ (.A(_06053_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__o21bai_1 _16571_ (.A1(_06054_),
    .A2(_06055_),
    .B1_N(_06053_),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_1 _16572_ (.A(_06053_),
    .B(_06056_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand3_1 _16573_ (.A(_06052_),
    .B(_06058_),
    .C(_06059_),
    .Y(_06061_));
 sky130_fd_sc_hd__a21o_1 _16574_ (.A1(_06058_),
    .A2(_06059_),
    .B1(_06052_),
    .X(_06062_));
 sky130_fd_sc_hd__nand2_1 _16575_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__a21oi_4 _16576_ (.A1(_05776_),
    .A2(_05783_),
    .B1(_05781_),
    .Y(_06064_));
 sky130_fd_sc_hd__o22a_2 _16577_ (.A1(_05020_),
    .A2(_04986_),
    .B1(_04989_),
    .B2(_03616_),
    .X(_06065_));
 sky130_fd_sc_hd__or3b_1 _16578_ (.A(_03835_),
    .B(net42),
    .C_N(net41),
    .X(_06066_));
 sky130_fd_sc_hd__nand3_2 _16579_ (.A(_05841_),
    .B(net265),
    .C(net279),
    .Y(_06067_));
 sky130_fd_sc_hd__o21a_1 _16580_ (.A1(_03835_),
    .A2(_04483_),
    .B1(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__and3_1 _16581_ (.A(_04102_),
    .B(net42),
    .C(net28),
    .X(_06069_));
 sky130_fd_sc_hd__a31oi_4 _16582_ (.A1(_05414_),
    .A2(_05446_),
    .A3(net243),
    .B1(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__a21oi_2 _16583_ (.A1(_06066_),
    .A2(_06067_),
    .B1(_06070_),
    .Y(_06072_));
 sky130_fd_sc_hd__a21o_1 _16584_ (.A1(_06066_),
    .A2(_06067_),
    .B1(_06070_),
    .X(_06073_));
 sky130_fd_sc_hd__o211a_1 _16585_ (.A1(_03835_),
    .A2(_04483_),
    .B1(_06067_),
    .C1(_06070_),
    .X(_06074_));
 sky130_fd_sc_hd__nand3b_4 _16586_ (.A_N(_06074_),
    .B(_06065_),
    .C(_06073_),
    .Y(_06075_));
 sky130_fd_sc_hd__o21bai_4 _16587_ (.A1(_06072_),
    .A2(_06074_),
    .B1_N(_06065_),
    .Y(_06076_));
 sky130_fd_sc_hd__a21oi_4 _16588_ (.A1(_06075_),
    .A2(_06076_),
    .B1(_06064_),
    .Y(_06077_));
 sky130_fd_sc_hd__a21o_1 _16589_ (.A1(_06075_),
    .A2(_06076_),
    .B1(_06064_),
    .X(_06078_));
 sky130_fd_sc_hd__and3_1 _16590_ (.A(_06075_),
    .B(_06076_),
    .C(_06064_),
    .X(_06079_));
 sky130_fd_sc_hd__a31oi_2 _16591_ (.A1(_06064_),
    .A2(_06075_),
    .A3(_06076_),
    .B1(_06063_),
    .Y(_06080_));
 sky130_fd_sc_hd__a31o_1 _16592_ (.A1(_06064_),
    .A2(_06075_),
    .A3(_06076_),
    .B1(_06063_),
    .X(_06081_));
 sky130_fd_sc_hd__o21ai_1 _16593_ (.A1(_06077_),
    .A2(_06079_),
    .B1(_06063_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_4 _16594_ (.A1(_06077_),
    .A2(_06081_),
    .B1(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__a21boi_1 _16595_ (.A1(_05754_),
    .A2(_05755_),
    .B1_N(_05752_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand2_1 _16596_ (.A(_05752_),
    .B(_05759_),
    .Y(_06086_));
 sky130_fd_sc_hd__a21o_2 _16597_ (.A1(_05831_),
    .A2(_05838_),
    .B1(_05836_),
    .X(_06087_));
 sky130_fd_sc_hd__a32o_1 _16598_ (.A1(_06486_),
    .A2(net261),
    .A3(net280),
    .B1(_04269_),
    .B2(net30),
    .X(_06088_));
 sky130_fd_sc_hd__nor2_1 _16599_ (.A(_03938_),
    .B(_04218_),
    .Y(_06089_));
 sky130_fd_sc_hd__a31oi_4 _16600_ (.A1(_07242_),
    .A2(net257),
    .A3(_04215_),
    .B1(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__or3_1 _16601_ (.A(net39),
    .B(_04037_),
    .C(_03949_),
    .X(_06091_));
 sky130_fd_sc_hd__o211ai_4 _16602_ (.A1(net261),
    .A2(_08656_),
    .B1(net285),
    .C1(_08700_),
    .Y(_06092_));
 sky130_fd_sc_hd__o311a_4 _16603_ (.A1(_03949_),
    .A2(_04037_),
    .A3(net39),
    .B1(_06092_),
    .C1(_06090_),
    .X(_06094_));
 sky130_fd_sc_hd__o221ai_4 _16604_ (.A1(_08711_),
    .A2(_03714_),
    .B1(_03737_),
    .B2(_03949_),
    .C1(_06090_),
    .Y(_06095_));
 sky130_fd_sc_hd__a21oi_4 _16605_ (.A1(_06091_),
    .A2(_06092_),
    .B1(_06090_),
    .Y(_06096_));
 sky130_fd_sc_hd__a21o_2 _16606_ (.A1(_06091_),
    .A2(_06092_),
    .B1(_06090_),
    .X(_06097_));
 sky130_fd_sc_hd__o21bai_4 _16607_ (.A1(_06094_),
    .A2(_06096_),
    .B1_N(_06088_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_2 _16608_ (.A(_06088_),
    .B(_06097_),
    .Y(_06099_));
 sky130_fd_sc_hd__and3_1 _16609_ (.A(_06088_),
    .B(_06095_),
    .C(_06097_),
    .X(_06100_));
 sky130_fd_sc_hd__nand3_2 _16610_ (.A(_06088_),
    .B(_06095_),
    .C(_06097_),
    .Y(_06101_));
 sky130_fd_sc_hd__o211a_1 _16611_ (.A1(_06094_),
    .A2(_06099_),
    .B1(_06098_),
    .C1(_06087_),
    .X(_06102_));
 sky130_fd_sc_hd__o211ai_4 _16612_ (.A1(_06094_),
    .A2(_06099_),
    .B1(_06098_),
    .C1(_06087_),
    .Y(_06103_));
 sky130_fd_sc_hd__a21oi_4 _16613_ (.A1(_06098_),
    .A2(_06101_),
    .B1(_06087_),
    .Y(_06105_));
 sky130_fd_sc_hd__nand3b_1 _16614_ (.A_N(_06105_),
    .B(_05748_),
    .C(_06103_),
    .Y(_06106_));
 sky130_fd_sc_hd__o22ai_2 _16615_ (.A1(_05740_),
    .A2(_05747_),
    .B1(_06102_),
    .B2(_06105_),
    .Y(_06107_));
 sky130_fd_sc_hd__a211o_1 _16616_ (.A1(_06098_),
    .A2(_06101_),
    .B1(_05748_),
    .C1(_06087_),
    .X(_06108_));
 sky130_fd_sc_hd__a31oi_1 _16617_ (.A1(_06087_),
    .A2(_06098_),
    .A3(_06101_),
    .B1(_05748_),
    .Y(_06109_));
 sky130_fd_sc_hd__o21ai_1 _16618_ (.A1(_05749_),
    .A2(_06105_),
    .B1(_06103_),
    .Y(_06110_));
 sky130_fd_sc_hd__o21ai_1 _16619_ (.A1(_06105_),
    .A2(_06109_),
    .B1(_06108_),
    .Y(_06111_));
 sky130_fd_sc_hd__o211a_1 _16620_ (.A1(_05749_),
    .A2(_06103_),
    .B1(_06085_),
    .C1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__o211ai_2 _16621_ (.A1(_05749_),
    .A2(_06103_),
    .B1(_06085_),
    .C1(_06111_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand3_2 _16622_ (.A(_06086_),
    .B(_06106_),
    .C(_06107_),
    .Y(_06114_));
 sky130_fd_sc_hd__a31o_1 _16623_ (.A1(_06086_),
    .A2(_06106_),
    .A3(_06107_),
    .B1(_06084_),
    .X(_06116_));
 sky130_fd_sc_hd__a21bo_1 _16624_ (.A1(_06113_),
    .A2(_06114_),
    .B1_N(_06084_),
    .X(_06117_));
 sky130_fd_sc_hd__nand3_1 _16625_ (.A(_06084_),
    .B(_06113_),
    .C(_06114_),
    .Y(_06118_));
 sky130_fd_sc_hd__a21o_1 _16626_ (.A1(_06113_),
    .A2(_06114_),
    .B1(_06084_),
    .X(_06119_));
 sky130_fd_sc_hd__o2bb2ai_2 _16627_ (.A1_N(_05848_),
    .A2_N(_05851_),
    .B1(_05849_),
    .B2(_05845_),
    .Y(_06120_));
 sky130_fd_sc_hd__nand4_2 _16628_ (.A(_05850_),
    .B(_05855_),
    .C(_06118_),
    .D(_06119_),
    .Y(_06121_));
 sky130_fd_sc_hd__o211ai_4 _16629_ (.A1(_06112_),
    .A2(_06116_),
    .B1(_06117_),
    .C1(_06120_),
    .Y(_06122_));
 sky130_fd_sc_hd__a21bo_1 _16630_ (.A1(_05760_),
    .A2(_05793_),
    .B1_N(_05761_),
    .X(_06123_));
 sky130_fd_sc_hd__a21oi_2 _16631_ (.A1(_06121_),
    .A2(_06122_),
    .B1(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__a21o_1 _16632_ (.A1(_06121_),
    .A2(_06122_),
    .B1(_06123_),
    .X(_06125_));
 sky130_fd_sc_hd__nand2_1 _16633_ (.A(_06121_),
    .B(_06123_),
    .Y(_06127_));
 sky130_fd_sc_hd__nand3_1 _16634_ (.A(_06121_),
    .B(_06122_),
    .C(_06123_),
    .Y(_06128_));
 sky130_fd_sc_hd__inv_2 _16635_ (.A(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__nor2_1 _16636_ (.A(_06124_),
    .B(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__nand2_1 _16637_ (.A(_06125_),
    .B(_06128_),
    .Y(_06131_));
 sky130_fd_sc_hd__o22ai_4 _16638_ (.A1(_05969_),
    .A2(_05974_),
    .B1(_05857_),
    .B2(_05977_),
    .Y(_06132_));
 sky130_fd_sc_hd__nand2_1 _16639_ (.A(_05827_),
    .B(_05846_),
    .Y(_06133_));
 sky130_fd_sc_hd__a21o_1 _16640_ (.A1(_05529_),
    .A2(_05878_),
    .B1(_05876_),
    .X(_06134_));
 sky130_fd_sc_hd__a21oi_2 _16641_ (.A1(_05529_),
    .A2(_05878_),
    .B1(_05876_),
    .Y(_06135_));
 sky130_fd_sc_hd__a32o_4 _16642_ (.A1(net255),
    .A2(_09698_),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net2),
    .X(_06136_));
 sky130_fd_sc_hd__o2111ai_4 _16643_ (.A1(_11387_),
    .A2(_12988_),
    .B1(net36),
    .C1(net235),
    .D1(_03993_),
    .Y(_06138_));
 sky130_fd_sc_hd__or3_2 _16644_ (.A(net36),
    .B(_04004_),
    .C(_03993_),
    .X(_06139_));
 sky130_fd_sc_hd__or3b_2 _16645_ (.A(_03982_),
    .B(net37),
    .C_N(net36),
    .X(_06140_));
 sky130_fd_sc_hd__o211ai_4 _16646_ (.A1(net261),
    .A2(_11387_),
    .B1(_01293_),
    .C1(_11354_),
    .Y(_06141_));
 sky130_fd_sc_hd__nand4_4 _16647_ (.A(_06138_),
    .B(_06139_),
    .C(_06140_),
    .D(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__a22oi_4 _16648_ (.A1(_06138_),
    .A2(_06139_),
    .B1(_06140_),
    .B2(_06141_),
    .Y(_06143_));
 sky130_fd_sc_hd__a21o_1 _16649_ (.A1(_06136_),
    .A2(_06142_),
    .B1(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__a21oi_4 _16650_ (.A1(_06136_),
    .A2(_06142_),
    .B1(_06143_),
    .Y(_06145_));
 sky130_fd_sc_hd__and2_2 _16651_ (.A(_06143_),
    .B(_06136_),
    .X(_06146_));
 sky130_fd_sc_hd__o22ai_4 _16652_ (.A1(_06136_),
    .A2(_06142_),
    .B1(_06145_),
    .B2(_06146_),
    .Y(_06147_));
 sky130_fd_sc_hd__a21oi_2 _16653_ (.A1(_05810_),
    .A2(_05818_),
    .B1(_05820_),
    .Y(_06149_));
 sky130_fd_sc_hd__a32o_2 _16654_ (.A1(_00625_),
    .A2(net250),
    .A3(net252),
    .B1(_11793_),
    .B2(net5),
    .X(_06150_));
 sky130_fd_sc_hd__o211ai_4 _16655_ (.A1(net254),
    .A2(_02442_),
    .B1(net289),
    .C1(_02421_),
    .Y(_06151_));
 sky130_fd_sc_hd__or3b_2 _16656_ (.A(net34),
    .B(_04026_),
    .C_N(net64),
    .X(_06152_));
 sky130_fd_sc_hd__o21ai_1 _16657_ (.A1(net263),
    .A2(net246),
    .B1(net291),
    .Y(_06153_));
 sky130_fd_sc_hd__a21oi_1 _16658_ (.A1(net7),
    .A2(net249),
    .B1(_06153_),
    .Y(_06154_));
 sky130_fd_sc_hd__a211o_1 _16659_ (.A1(_11420_),
    .A2(net282),
    .B1(_08261_),
    .C1(net247),
    .X(_06155_));
 sky130_fd_sc_hd__nor2_1 _16660_ (.A(_04048_),
    .B(_08283_),
    .Y(_06156_));
 sky130_fd_sc_hd__o2bb2a_2 _16661_ (.A1_N(_06151_),
    .A2_N(_06152_),
    .B1(_06154_),
    .B2(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__o2bb2ai_2 _16662_ (.A1_N(_06151_),
    .A2_N(_06152_),
    .B1(_06154_),
    .B2(_06156_),
    .Y(_06158_));
 sky130_fd_sc_hd__o211ai_1 _16663_ (.A1(net247),
    .A2(_06153_),
    .B1(_06152_),
    .C1(_06151_),
    .Y(_06160_));
 sky130_fd_sc_hd__o2111ai_4 _16664_ (.A1(_04048_),
    .A2(_08283_),
    .B1(_06151_),
    .C1(_06152_),
    .D1(_06155_),
    .Y(_06161_));
 sky130_fd_sc_hd__o211a_4 _16665_ (.A1(_06160_),
    .A2(_06156_),
    .B1(_06150_),
    .C1(_06158_),
    .X(_06162_));
 sky130_fd_sc_hd__a21oi_4 _16666_ (.A1(_06158_),
    .A2(_06161_),
    .B1(_06150_),
    .Y(_06163_));
 sky130_fd_sc_hd__nor3_4 _16667_ (.A(_06149_),
    .B(_06162_),
    .C(_06163_),
    .Y(_06164_));
 sky130_fd_sc_hd__a211o_1 _16668_ (.A1(_05821_),
    .A2(_05823_),
    .B1(_06162_),
    .C1(_06163_),
    .X(_06165_));
 sky130_fd_sc_hd__o21a_1 _16669_ (.A1(_06162_),
    .A2(_06163_),
    .B1(_06149_),
    .X(_06166_));
 sky130_fd_sc_hd__o21ai_2 _16670_ (.A1(_06162_),
    .A2(_06163_),
    .B1(_06149_),
    .Y(_06167_));
 sky130_fd_sc_hd__o221a_1 _16671_ (.A1(_06136_),
    .A2(_06142_),
    .B1(_06145_),
    .B2(_06146_),
    .C1(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__o221ai_4 _16672_ (.A1(_06136_),
    .A2(_06142_),
    .B1(_06145_),
    .B2(_06146_),
    .C1(_06167_),
    .Y(_06169_));
 sky130_fd_sc_hd__nand3b_1 _16673_ (.A_N(_06147_),
    .B(_06165_),
    .C(_06167_),
    .Y(_06171_));
 sky130_fd_sc_hd__o21ai_4 _16674_ (.A1(_06164_),
    .A2(_06166_),
    .B1(_06147_),
    .Y(_06172_));
 sky130_fd_sc_hd__o21ai_2 _16675_ (.A1(_06164_),
    .A2(_06169_),
    .B1(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__o211a_1 _16676_ (.A1(_06164_),
    .A2(_06169_),
    .B1(_06172_),
    .C1(_06135_),
    .X(_06174_));
 sky130_fd_sc_hd__o211ai_2 _16677_ (.A1(_06164_),
    .A2(_06169_),
    .B1(_06172_),
    .C1(_06135_),
    .Y(_06175_));
 sky130_fd_sc_hd__a21oi_1 _16678_ (.A1(_06171_),
    .A2(_06172_),
    .B1(_06135_),
    .Y(_06176_));
 sky130_fd_sc_hd__a21o_2 _16679_ (.A1(_06171_),
    .A2(_06172_),
    .B1(_06135_),
    .X(_06177_));
 sky130_fd_sc_hd__o211a_4 _16680_ (.A1(_05828_),
    .A2(_05845_),
    .B1(_06175_),
    .C1(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__o211a_1 _16681_ (.A1(_06174_),
    .A2(_06176_),
    .B1(_05827_),
    .C1(_05846_),
    .X(_06179_));
 sky130_fd_sc_hd__nand4_2 _16682_ (.A(_05827_),
    .B(_05846_),
    .C(_06175_),
    .D(_06177_),
    .Y(_06180_));
 sky130_fd_sc_hd__o22ai_2 _16683_ (.A1(_05828_),
    .A2(_05845_),
    .B1(_06174_),
    .B2(_06176_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_1 _16684_ (.A(_06180_),
    .B(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__a21boi_4 _16685_ (.A1(_05862_),
    .A2(_05869_),
    .B1_N(_05870_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _16686_ (.A(_05870_),
    .B(_05872_),
    .Y(_06185_));
 sky130_fd_sc_hd__and3_1 _16687_ (.A(_04132_),
    .B(_07658_),
    .C(net230),
    .X(_06186_));
 sky130_fd_sc_hd__nor2_1 _16688_ (.A(_04059_),
    .B(_07691_),
    .Y(_06187_));
 sky130_fd_sc_hd__o22a_2 _16689_ (.A1(_04059_),
    .A2(_07691_),
    .B1(_04133_),
    .B2(_07669_),
    .X(_06188_));
 sky130_fd_sc_hd__nand3_4 _16690_ (.A(net224),
    .B(net292),
    .C(net188),
    .Y(_06189_));
 sky130_fd_sc_hd__or3b_4 _16691_ (.A(net62),
    .B(_04069_),
    .C_N(net61),
    .X(_06190_));
 sky130_fd_sc_hd__or3b_2 _16692_ (.A(net61),
    .B(_04080_),
    .C_N(net60),
    .X(_06191_));
 sky130_fd_sc_hd__o211ai_4 _16693_ (.A1(net232),
    .A2(_04557_),
    .B1(net299),
    .C1(net219),
    .Y(_06193_));
 sky130_fd_sc_hd__o2111a_2 _16694_ (.A1(_04080_),
    .A2(net298),
    .B1(_06189_),
    .C1(_06190_),
    .D1(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__o2111ai_4 _16695_ (.A1(_04080_),
    .A2(net298),
    .B1(_06189_),
    .C1(_06190_),
    .D1(_06193_),
    .Y(_06195_));
 sky130_fd_sc_hd__a22oi_4 _16696_ (.A1(_06189_),
    .A2(_06190_),
    .B1(_06191_),
    .B2(_06193_),
    .Y(_06196_));
 sky130_fd_sc_hd__a22o_1 _16697_ (.A1(_06189_),
    .A2(_06190_),
    .B1(_06191_),
    .B2(_06193_),
    .X(_06197_));
 sky130_fd_sc_hd__o21ai_1 _16698_ (.A1(_06188_),
    .A2(_06194_),
    .B1(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__o21a_1 _16699_ (.A1(_06188_),
    .A2(_06194_),
    .B1(_06197_),
    .X(_06199_));
 sky130_fd_sc_hd__o22ai_4 _16700_ (.A1(_06186_),
    .A2(_06187_),
    .B1(_06194_),
    .B2(_06196_),
    .Y(_06200_));
 sky130_fd_sc_hd__nand3_4 _16701_ (.A(_06197_),
    .B(_06188_),
    .C(_06195_),
    .Y(_06201_));
 sky130_fd_sc_hd__o211ai_1 _16702_ (.A1(_06186_),
    .A2(_06187_),
    .B1(_06195_),
    .C1(_06197_),
    .Y(_06202_));
 sky130_fd_sc_hd__o21ai_1 _16703_ (.A1(_06194_),
    .A2(_06196_),
    .B1(_06188_),
    .Y(_06204_));
 sky130_fd_sc_hd__a21oi_2 _16704_ (.A1(_06200_),
    .A2(_06201_),
    .B1(_05908_),
    .Y(_06205_));
 sky130_fd_sc_hd__nand3_2 _16705_ (.A(_06204_),
    .B(_05906_),
    .C(_06202_),
    .Y(_06206_));
 sky130_fd_sc_hd__nand3_2 _16706_ (.A(_05908_),
    .B(_06200_),
    .C(_06201_),
    .Y(_06207_));
 sky130_fd_sc_hd__a21oi_2 _16707_ (.A1(_06206_),
    .A2(_06207_),
    .B1(_06184_),
    .Y(_06208_));
 sky130_fd_sc_hd__and3_1 _16708_ (.A(_06206_),
    .B(_06207_),
    .C(_06184_),
    .X(_06209_));
 sky130_fd_sc_hd__a21oi_1 _16709_ (.A1(_06206_),
    .A2(_06207_),
    .B1(_06185_),
    .Y(_06210_));
 sky130_fd_sc_hd__a21o_1 _16710_ (.A1(_06206_),
    .A2(_06207_),
    .B1(_06185_),
    .X(_06211_));
 sky130_fd_sc_hd__and3_1 _16711_ (.A(_06185_),
    .B(_06206_),
    .C(_06207_),
    .X(_06212_));
 sky130_fd_sc_hd__nand3_1 _16712_ (.A(_06185_),
    .B(_06206_),
    .C(_06207_),
    .Y(_06213_));
 sky130_fd_sc_hd__nand2_1 _16713_ (.A(_06211_),
    .B(_06213_),
    .Y(_06215_));
 sky130_fd_sc_hd__nor2_2 _16714_ (.A(_04146_),
    .B(_04375_),
    .Y(_06216_));
 sky130_fd_sc_hd__o311a_1 _16715_ (.A1(net232),
    .A2(_04787_),
    .A3(_05551_),
    .B1(_05549_),
    .C1(_04342_),
    .X(_06217_));
 sky130_fd_sc_hd__a31oi_4 _16716_ (.A1(_05549_),
    .A2(_05553_),
    .A3(_04342_),
    .B1(_06216_),
    .Y(_06218_));
 sky130_fd_sc_hd__o21ai_4 _16717_ (.A1(net245),
    .A2(net241),
    .B1(net17),
    .Y(_06219_));
 sky130_fd_sc_hd__nand4b_4 _16718_ (.A_N(_11409_),
    .B(_04168_),
    .C(net308),
    .D(_03953_),
    .Y(_06220_));
 sky130_fd_sc_hd__nand4_4 _16719_ (.A(_06519_),
    .B(_03955_),
    .C(_05926_),
    .D(_04168_),
    .Y(_06221_));
 sky130_fd_sc_hd__o21ai_4 _16720_ (.A1(_05927_),
    .A2(_06220_),
    .B1(net201),
    .Y(_06222_));
 sky130_fd_sc_hd__o211ai_2 _16721_ (.A1(_05927_),
    .A2(_06220_),
    .B1(net33),
    .C1(_06219_),
    .Y(_06223_));
 sky130_fd_sc_hd__o211ai_4 _16722_ (.A1(net232),
    .A2(_05927_),
    .B1(_04484_),
    .C1(_05933_),
    .Y(_06224_));
 sky130_fd_sc_hd__nor2_1 _16723_ (.A(_04157_),
    .B(_04331_),
    .Y(_06226_));
 sky130_fd_sc_hd__or3_1 _16724_ (.A(net44),
    .B(_04157_),
    .C(_03286_),
    .X(_06227_));
 sky130_fd_sc_hd__and4_1 _16725_ (.A(_06219_),
    .B(_06221_),
    .C(_06226_),
    .D(net33),
    .X(_06228_));
 sky130_fd_sc_hd__nand4_4 _16726_ (.A(_06219_),
    .B(_06221_),
    .C(_06226_),
    .D(net33),
    .Y(_06229_));
 sky130_fd_sc_hd__o311a_2 _16727_ (.A1(_03286_),
    .A2(net44),
    .A3(_04157_),
    .B1(_06223_),
    .C1(_06224_),
    .X(_06230_));
 sky130_fd_sc_hd__o221ai_2 _16728_ (.A1(_04157_),
    .A2(_04331_),
    .B1(_06222_),
    .B2(_03286_),
    .C1(_06224_),
    .Y(_06231_));
 sky130_fd_sc_hd__o21ai_2 _16729_ (.A1(_06228_),
    .A2(_06230_),
    .B1(_06218_),
    .Y(_06232_));
 sky130_fd_sc_hd__o211ai_2 _16730_ (.A1(_06216_),
    .A2(_06217_),
    .B1(_06229_),
    .C1(_06231_),
    .Y(_06233_));
 sky130_fd_sc_hd__o22ai_2 _16731_ (.A1(_06216_),
    .A2(_06217_),
    .B1(_06228_),
    .B2(_06230_),
    .Y(_06234_));
 sky130_fd_sc_hd__nand3_1 _16732_ (.A(_06231_),
    .B(_06218_),
    .C(_06229_),
    .Y(_06235_));
 sky130_fd_sc_hd__a32oi_4 _16733_ (.A1(_05921_),
    .A2(_05923_),
    .A3(_05936_),
    .B1(_05938_),
    .B2(_05919_),
    .Y(_06237_));
 sky130_fd_sc_hd__a32o_1 _16734_ (.A1(_05921_),
    .A2(_05923_),
    .A3(_05936_),
    .B1(_05919_),
    .B2(_05938_),
    .X(_06238_));
 sky130_fd_sc_hd__nand3_4 _16735_ (.A(_06234_),
    .B(_06235_),
    .C(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__and3_1 _16736_ (.A(_06232_),
    .B(_06233_),
    .C(_06237_),
    .X(_06240_));
 sky130_fd_sc_hd__nand3_4 _16737_ (.A(_06232_),
    .B(_06233_),
    .C(_06237_),
    .Y(_06241_));
 sky130_fd_sc_hd__a22oi_2 _16738_ (.A1(net11),
    .A2(_05249_),
    .B1(_04792_),
    .B2(_05227_),
    .Y(_06242_));
 sky130_fd_sc_hd__a32o_1 _16739_ (.A1(net215),
    .A2(_05227_),
    .A3(net185),
    .B1(_05249_),
    .B2(net11),
    .X(_06243_));
 sky130_fd_sc_hd__a32oi_4 _16740_ (.A1(net212),
    .A2(net183),
    .A3(net305),
    .B1(_04911_),
    .B2(net13),
    .Y(_06244_));
 sky130_fd_sc_hd__nand3_2 _16741_ (.A(net181),
    .B(net180),
    .C(net317),
    .Y(_06245_));
 sky130_fd_sc_hd__or3b_2 _16742_ (.A(net58),
    .B(_04135_),
    .C_N(net55),
    .X(_06246_));
 sky130_fd_sc_hd__a21oi_2 _16743_ (.A1(_06245_),
    .A2(_06246_),
    .B1(_06244_),
    .Y(_06248_));
 sky130_fd_sc_hd__a21o_1 _16744_ (.A1(_06245_),
    .A2(_06246_),
    .B1(_06244_),
    .X(_06249_));
 sky130_fd_sc_hd__o221ai_4 _16745_ (.A1(_04135_),
    .A2(net316),
    .B1(_05294_),
    .B2(_04638_),
    .C1(_06244_),
    .Y(_06250_));
 sky130_fd_sc_hd__a21oi_1 _16746_ (.A1(_06249_),
    .A2(_06250_),
    .B1(_06243_),
    .Y(_06251_));
 sky130_fd_sc_hd__a21o_1 _16747_ (.A1(_06249_),
    .A2(_06250_),
    .B1(_06243_),
    .X(_06252_));
 sky130_fd_sc_hd__a31oi_4 _16748_ (.A1(_06244_),
    .A2(_06245_),
    .A3(_06246_),
    .B1(_06242_),
    .Y(_06253_));
 sky130_fd_sc_hd__and3_1 _16749_ (.A(_06243_),
    .B(_06249_),
    .C(_06250_),
    .X(_06254_));
 sky130_fd_sc_hd__nand2_1 _16750_ (.A(_06253_),
    .B(_06249_),
    .Y(_06255_));
 sky130_fd_sc_hd__nand3_2 _16751_ (.A(_06239_),
    .B(_06252_),
    .C(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__nand4_2 _16752_ (.A(_06239_),
    .B(_06241_),
    .C(_06252_),
    .D(_06255_),
    .Y(_06257_));
 sky130_fd_sc_hd__o2bb2ai_4 _16753_ (.A1_N(_06239_),
    .A2_N(_06241_),
    .B1(_06251_),
    .B2(_06254_),
    .Y(_06259_));
 sky130_fd_sc_hd__a2bb2oi_4 _16754_ (.A1_N(_05948_),
    .A2_N(_05952_),
    .B1(_06257_),
    .B2(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__a21o_1 _16755_ (.A1(_06257_),
    .A2(_06259_),
    .B1(_05953_),
    .X(_06261_));
 sky130_fd_sc_hd__o211a_1 _16756_ (.A1(_06240_),
    .A2(_06256_),
    .B1(_06259_),
    .C1(_05953_),
    .X(_06262_));
 sky130_fd_sc_hd__o211ai_4 _16757_ (.A1(_06240_),
    .A2(_06256_),
    .B1(_06259_),
    .C1(_05953_),
    .Y(_06263_));
 sky130_fd_sc_hd__nand3_2 _16758_ (.A(_06261_),
    .B(_06263_),
    .C(_06215_),
    .Y(_06264_));
 sky130_fd_sc_hd__o22ai_4 _16759_ (.A1(_06208_),
    .A2(_06209_),
    .B1(_06260_),
    .B2(_06262_),
    .Y(_06265_));
 sky130_fd_sc_hd__o21a_1 _16760_ (.A1(_06210_),
    .A2(_06212_),
    .B1(_06263_),
    .X(_06266_));
 sky130_fd_sc_hd__o21ai_4 _16761_ (.A1(_06215_),
    .A2(_06260_),
    .B1(_06263_),
    .Y(_06267_));
 sky130_fd_sc_hd__inv_2 _16762_ (.A(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__o211ai_2 _16763_ (.A1(_06208_),
    .A2(_06209_),
    .B1(_06261_),
    .C1(_06263_),
    .Y(_06270_));
 sky130_fd_sc_hd__o22ai_2 _16764_ (.A1(_06210_),
    .A2(_06212_),
    .B1(_06260_),
    .B2(_06262_),
    .Y(_06271_));
 sky130_fd_sc_hd__nand2_1 _16765_ (.A(_06270_),
    .B(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__a2bb2oi_4 _16766_ (.A1_N(_05964_),
    .A2_N(_05966_),
    .B1(_06264_),
    .B2(_06265_),
    .Y(_06273_));
 sky130_fd_sc_hd__a21oi_2 _16767_ (.A1(_06270_),
    .A2(_06271_),
    .B1(_05968_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand3_2 _16768_ (.A(_05967_),
    .B(_06264_),
    .C(_06265_),
    .Y(_06275_));
 sky130_fd_sc_hd__a22oi_4 _16769_ (.A1(_06180_),
    .A2(_06182_),
    .B1(_06272_),
    .B2(_05967_),
    .Y(_06276_));
 sky130_fd_sc_hd__nand2_1 _16770_ (.A(_06275_),
    .B(_06183_),
    .Y(_06277_));
 sky130_fd_sc_hd__nand3b_2 _16771_ (.A_N(_06273_),
    .B(_06275_),
    .C(_06183_),
    .Y(_06278_));
 sky130_fd_sc_hd__o22ai_4 _16772_ (.A1(_06178_),
    .A2(_06179_),
    .B1(_06273_),
    .B2(_06274_),
    .Y(_06279_));
 sky130_fd_sc_hd__o211a_1 _16773_ (.A1(_06273_),
    .A2(_06277_),
    .B1(_06279_),
    .C1(_06132_),
    .X(_06280_));
 sky130_fd_sc_hd__o211ai_4 _16774_ (.A1(_06273_),
    .A2(_06277_),
    .B1(_06279_),
    .C1(_06132_),
    .Y(_06281_));
 sky130_fd_sc_hd__a21oi_4 _16775_ (.A1(_06278_),
    .A2(_06279_),
    .B1(_06132_),
    .Y(_06282_));
 sky130_fd_sc_hd__a21o_1 _16776_ (.A1(_06278_),
    .A2(_06279_),
    .B1(_06132_),
    .X(_06283_));
 sky130_fd_sc_hd__o211ai_1 _16777_ (.A1(_06124_),
    .A2(_06129_),
    .B1(_06281_),
    .C1(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__o21ai_1 _16778_ (.A1(_06280_),
    .A2(_06282_),
    .B1(_06130_),
    .Y(_06285_));
 sky130_fd_sc_hd__nand3_4 _16779_ (.A(_06130_),
    .B(_06281_),
    .C(_06283_),
    .Y(_06286_));
 sky130_fd_sc_hd__o22ai_4 _16780_ (.A1(_06124_),
    .A2(_06129_),
    .B1(_06280_),
    .B2(_06282_),
    .Y(_06287_));
 sky130_fd_sc_hd__o211a_2 _16781_ (.A1(_05983_),
    .A2(_05987_),
    .B1(_06286_),
    .C1(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__o211ai_2 _16782_ (.A1(_05983_),
    .A2(_05987_),
    .B1(_06286_),
    .C1(_06287_),
    .Y(_06289_));
 sky130_fd_sc_hd__a22oi_4 _16783_ (.A1(_05986_),
    .A2(_06050_),
    .B1(_06286_),
    .B2(_06287_),
    .Y(_06291_));
 sky130_fd_sc_hd__a22o_1 _16784_ (.A1(_05986_),
    .A2(_06050_),
    .B1(_06286_),
    .B2(_06287_),
    .X(_06292_));
 sky130_fd_sc_hd__o22ai_4 _16785_ (.A1(_06045_),
    .A2(_06046_),
    .B1(_06288_),
    .B2(_06291_),
    .Y(_06293_));
 sky130_fd_sc_hd__o211ai_4 _16786_ (.A1(_06043_),
    .A2(_06044_),
    .B1(_06289_),
    .C1(_06292_),
    .Y(_06294_));
 sky130_fd_sc_hd__a31o_1 _16787_ (.A1(_06051_),
    .A2(_06284_),
    .A3(_06285_),
    .B1(_06048_),
    .X(_06295_));
 sky130_fd_sc_hd__o22ai_2 _16788_ (.A1(_06043_),
    .A2(_06044_),
    .B1(_06288_),
    .B2(_06291_),
    .Y(_06296_));
 sky130_fd_sc_hd__o211a_2 _16789_ (.A1(_06288_),
    .A2(_06295_),
    .B1(_06024_),
    .C1(_06296_),
    .X(_06297_));
 sky130_fd_sc_hd__o211ai_4 _16790_ (.A1(_06288_),
    .A2(_06295_),
    .B1(_06024_),
    .C1(_06296_),
    .Y(_06298_));
 sky130_fd_sc_hd__nand3_2 _16791_ (.A(_06025_),
    .B(_06293_),
    .C(_06294_),
    .Y(_06299_));
 sky130_fd_sc_hd__o2bb2ai_4 _16792_ (.A1_N(_06298_),
    .A2_N(_06299_),
    .B1(_05717_),
    .B2(_05718_),
    .Y(_06300_));
 sky130_fd_sc_hd__a31oi_4 _16793_ (.A1(_06025_),
    .A2(_06293_),
    .A3(_06294_),
    .B1(_05721_),
    .Y(_06302_));
 sky130_fd_sc_hd__a31o_1 _16794_ (.A1(_06025_),
    .A2(_06293_),
    .A3(_06294_),
    .B1(_05721_),
    .X(_06303_));
 sky130_fd_sc_hd__nand3_2 _16795_ (.A(_06299_),
    .B(_05719_),
    .C(_06298_),
    .Y(_06304_));
 sky130_fd_sc_hd__a21o_2 _16796_ (.A1(_06008_),
    .A2(_05687_),
    .B1(_06004_),
    .X(_06305_));
 sky130_fd_sc_hd__a21o_1 _16797_ (.A1(_06300_),
    .A2(_06304_),
    .B1(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__o211ai_1 _16798_ (.A1(_06297_),
    .A2(_06303_),
    .B1(_06300_),
    .C1(_06305_),
    .Y(_06307_));
 sky130_fd_sc_hd__a21oi_1 _16799_ (.A1(_06306_),
    .A2(_06307_),
    .B1(_06016_),
    .Y(_06308_));
 sky130_fd_sc_hd__nand2_1 _16800_ (.A(_06306_),
    .B(_06016_),
    .Y(_06309_));
 sky130_fd_sc_hd__a21oi_2 _16801_ (.A1(_06016_),
    .A2(_06306_),
    .B1(_06308_),
    .Y(_06310_));
 sky130_fd_sc_hd__nand3_1 _16802_ (.A(_05712_),
    .B(_06019_),
    .C(_06020_),
    .Y(_06311_));
 sky130_fd_sc_hd__a31oi_2 _16803_ (.A1(_05445_),
    .A2(_04942_),
    .A3(_04934_),
    .B1(_05444_),
    .Y(_06313_));
 sky130_fd_sc_hd__a22o_1 _16804_ (.A1(_05439_),
    .A2(_05705_),
    .B1(_05707_),
    .B2(_06015_),
    .X(_06314_));
 sky130_fd_sc_hd__o2bb2ai_4 _16805_ (.A1_N(_06019_),
    .A2_N(_06314_),
    .B1(_06311_),
    .B2(_06313_),
    .Y(_06315_));
 sky130_fd_sc_hd__and4_1 _16806_ (.A(_05445_),
    .B(_05712_),
    .C(_06019_),
    .D(_06020_),
    .X(_06316_));
 sky130_fd_sc_hd__nand4_2 _16807_ (.A(_05445_),
    .B(_05712_),
    .C(_06019_),
    .D(_06020_),
    .Y(_06317_));
 sky130_fd_sc_hd__a211oi_4 _16808_ (.A1(_04066_),
    .A2(_04259_),
    .B1(_04938_),
    .C1(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__a21oi_4 _16809_ (.A1(_04939_),
    .A2(_06316_),
    .B1(_06315_),
    .Y(_06319_));
 sky130_fd_sc_hd__a21o_1 _16810_ (.A1(_04939_),
    .A2(_06316_),
    .B1(_06315_),
    .X(_06320_));
 sky130_fd_sc_hd__xnor2_1 _16811_ (.A(_06310_),
    .B(_06319_),
    .Y(net81));
 sky130_fd_sc_hd__a21oi_1 _16812_ (.A1(_06299_),
    .A2(_05719_),
    .B1(_06297_),
    .Y(_06321_));
 sky130_fd_sc_hd__a41oi_4 _16813_ (.A1(_05986_),
    .A2(_06050_),
    .A3(_06286_),
    .A4(_06287_),
    .B1(_06047_),
    .Y(_06322_));
 sky130_fd_sc_hd__o21ai_1 _16814_ (.A1(_06048_),
    .A2(_06291_),
    .B1(_06289_),
    .Y(_06323_));
 sky130_fd_sc_hd__and2b_4 _16815_ (.A_N(net49),
    .B(net50),
    .X(_06324_));
 sky130_fd_sc_hd__nand2b_4 _16816_ (.A_N(net49),
    .B(net50),
    .Y(_06325_));
 sky130_fd_sc_hd__and2b_4 _16817_ (.A_N(net50),
    .B(net49),
    .X(_06326_));
 sky130_fd_sc_hd__o21a_1 _16818_ (.A1(_06324_),
    .A2(_06326_),
    .B1(net1),
    .X(_06327_));
 sky130_fd_sc_hd__o21ai_1 _16819_ (.A1(_06324_),
    .A2(_06326_),
    .B1(net1),
    .Y(_06328_));
 sky130_fd_sc_hd__a21oi_1 _16820_ (.A1(_04309_),
    .A2(_04517_),
    .B1(_06028_),
    .Y(_06329_));
 sky130_fd_sc_hd__and3b_1 _16821_ (.A_N(net49),
    .B(net48),
    .C(net12),
    .X(_06330_));
 sky130_fd_sc_hd__o2bb2a_1 _16822_ (.A1_N(net12),
    .A2_N(_06029_),
    .B1(_06028_),
    .B2(_04528_),
    .X(_06331_));
 sky130_fd_sc_hd__a22o_1 _16823_ (.A1(net12),
    .A2(_06029_),
    .B1(_04539_),
    .B2(_06026_),
    .X(_06333_));
 sky130_fd_sc_hd__o221a_1 _16824_ (.A1(_06324_),
    .A2(_06326_),
    .B1(_06329_),
    .B2(_06330_),
    .C1(net1),
    .X(_06334_));
 sky130_fd_sc_hd__o21ai_1 _16825_ (.A1(_06329_),
    .A2(_06330_),
    .B1(_06327_),
    .Y(_06335_));
 sky130_fd_sc_hd__a211o_1 _16826_ (.A1(_06026_),
    .A2(_04539_),
    .B1(_06330_),
    .C1(_06327_),
    .X(_06336_));
 sky130_fd_sc_hd__nand2_2 _16827_ (.A(_06335_),
    .B(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__a21oi_2 _16828_ (.A1(_06052_),
    .A2(_06059_),
    .B1(_06057_),
    .Y(_06338_));
 sky130_fd_sc_hd__a21oi_1 _16829_ (.A1(_06058_),
    .A2(_06061_),
    .B1(_06337_),
    .Y(_06339_));
 sky130_fd_sc_hd__xnor2_1 _16830_ (.A(_06337_),
    .B(_06338_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand3_2 _16831_ (.A(_06078_),
    .B(_06081_),
    .C(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__o21bai_4 _16832_ (.A1(_06077_),
    .A2(_06080_),
    .B1_N(_06340_),
    .Y(_06342_));
 sky130_fd_sc_hd__nand2_1 _16833_ (.A(_06341_),
    .B(_06342_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand3_1 _16834_ (.A(_06341_),
    .B(_06342_),
    .C(_06033_),
    .Y(_06345_));
 sky130_fd_sc_hd__a21o_1 _16835_ (.A1(_06341_),
    .A2(_06342_),
    .B1(_06033_),
    .X(_06346_));
 sky130_fd_sc_hd__and3_1 _16836_ (.A(_06037_),
    .B(_06341_),
    .C(_06342_),
    .X(_06347_));
 sky130_fd_sc_hd__o2bb2a_1 _16837_ (.A1_N(_06345_),
    .A2_N(_06346_),
    .B1(_06035_),
    .B2(_06036_),
    .X(_06348_));
 sky130_fd_sc_hd__a31o_1 _16838_ (.A1(_06037_),
    .A2(_06341_),
    .A3(_06342_),
    .B1(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__a21oi_2 _16839_ (.A1(_06122_),
    .A2(_06127_),
    .B1(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__a21o_1 _16840_ (.A1(_06122_),
    .A2(_06127_),
    .B1(_06349_),
    .X(_06351_));
 sky130_fd_sc_hd__o211ai_1 _16841_ (.A1(_06347_),
    .A2(_06348_),
    .B1(_06122_),
    .C1(_06128_),
    .Y(_06352_));
 sky130_fd_sc_hd__nand2_1 _16842_ (.A(_06351_),
    .B(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__a2bb2o_1 _16843_ (.A1_N(_05716_),
    .A2_N(_06040_),
    .B1(_06351_),
    .B2(_06352_),
    .X(_06355_));
 sky130_fd_sc_hd__and4bb_1 _16844_ (.A_N(_05716_),
    .B_N(_06040_),
    .C(_06351_),
    .D(_06352_),
    .X(_06356_));
 sky130_fd_sc_hd__o41a_1 _16845_ (.A1(_05716_),
    .A2(_06037_),
    .A3(_06039_),
    .A4(_06353_),
    .B1(_06355_),
    .X(_06357_));
 sky130_fd_sc_hd__o41ai_2 _16846_ (.A1(_05716_),
    .A2(_06037_),
    .A3(_06039_),
    .A4(_06353_),
    .B1(_06355_),
    .Y(_06358_));
 sky130_fd_sc_hd__o21ai_1 _16847_ (.A1(_06131_),
    .A2(_06282_),
    .B1(_06281_),
    .Y(_06359_));
 sky130_fd_sc_hd__a21oi_1 _16848_ (.A1(_06068_),
    .A2(_06070_),
    .B1(_06065_),
    .Y(_06360_));
 sky130_fd_sc_hd__a31o_1 _16849_ (.A1(_06066_),
    .A2(_06067_),
    .A3(_06070_),
    .B1(_06065_),
    .X(_06361_));
 sky130_fd_sc_hd__o22a_1 _16850_ (.A1(_05457_),
    .A2(_04986_),
    .B1(_04989_),
    .B2(_03725_),
    .X(_06362_));
 sky130_fd_sc_hd__or3b_1 _16851_ (.A(_03835_),
    .B(net43),
    .C_N(net42),
    .X(_06363_));
 sky130_fd_sc_hd__nand3_2 _16852_ (.A(_05841_),
    .B(net265),
    .C(net243),
    .Y(_06364_));
 sky130_fd_sc_hd__nor2_1 _16853_ (.A(_03916_),
    .B(_04483_),
    .Y(_06366_));
 sky130_fd_sc_hd__or3b_1 _16854_ (.A(_03916_),
    .B(net42),
    .C_N(net41),
    .X(_06367_));
 sky130_fd_sc_hd__a221oi_2 _16855_ (.A1(net306),
    .A2(_06497_),
    .B1(net265),
    .B2(net30),
    .C1(_04481_),
    .Y(_06368_));
 sky130_fd_sc_hd__o211ai_2 _16856_ (.A1(_04747_),
    .A2(net264),
    .B1(net279),
    .C1(_06486_),
    .Y(_06369_));
 sky130_fd_sc_hd__o2bb2ai_2 _16857_ (.A1_N(_06363_),
    .A2_N(_06364_),
    .B1(_06366_),
    .B2(_06368_),
    .Y(_06370_));
 sky130_fd_sc_hd__and4_1 _16858_ (.A(_06363_),
    .B(_06364_),
    .C(_06367_),
    .D(_06369_),
    .X(_06371_));
 sky130_fd_sc_hd__o2111ai_4 _16859_ (.A1(_03835_),
    .A2(_04898_),
    .B1(_06364_),
    .C1(_06367_),
    .D1(_06369_),
    .Y(_06372_));
 sky130_fd_sc_hd__nand2_1 _16860_ (.A(_06370_),
    .B(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__nor2_1 _16861_ (.A(_06362_),
    .B(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand3_1 _16862_ (.A(_06362_),
    .B(_06370_),
    .C(_06372_),
    .Y(_06375_));
 sky130_fd_sc_hd__a21o_1 _16863_ (.A1(_06370_),
    .A2(_06372_),
    .B1(_06362_),
    .X(_06377_));
 sky130_fd_sc_hd__o2111ai_2 _16864_ (.A1(_06068_),
    .A2(_06070_),
    .B1(_06361_),
    .C1(_06375_),
    .D1(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__o2bb2ai_1 _16865_ (.A1_N(_06362_),
    .A2_N(_06373_),
    .B1(_06072_),
    .B2(_06360_),
    .Y(_06379_));
 sky130_fd_sc_hd__o21ai_1 _16866_ (.A1(_06374_),
    .A2(_06379_),
    .B1(_06378_),
    .Y(_06380_));
 sky130_fd_sc_hd__a32o_1 _16867_ (.A1(net318),
    .A2(_04452_),
    .A3(net275),
    .B1(_05765_),
    .B2(net23),
    .X(_06381_));
 sky130_fd_sc_hd__or3_1 _16868_ (.A(net46),
    .B(_04124_),
    .C(_03616_),
    .X(_06382_));
 sky130_fd_sc_hd__nand3_2 _16869_ (.A(net266),
    .B(net303),
    .C(net276),
    .Y(_06383_));
 sky130_fd_sc_hd__nor2_2 _16870_ (.A(_03506_),
    .B(_05465_),
    .Y(_06384_));
 sky130_fd_sc_hd__a31oi_2 _16871_ (.A1(net313),
    .A2(_04747_),
    .A3(_05462_),
    .B1(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__o221ai_4 _16872_ (.A1(_03616_),
    .A2(_05229_),
    .B1(_05463_),
    .B2(_04758_),
    .C1(_06383_),
    .Y(_06386_));
 sky130_fd_sc_hd__and3_1 _16873_ (.A(_06385_),
    .B(_06383_),
    .C(_06382_),
    .X(_06388_));
 sky130_fd_sc_hd__o211ai_1 _16874_ (.A1(_03616_),
    .A2(_05229_),
    .B1(_06383_),
    .C1(_06385_),
    .Y(_06389_));
 sky130_fd_sc_hd__a21oi_1 _16875_ (.A1(_06382_),
    .A2(_06383_),
    .B1(_06385_),
    .Y(_06390_));
 sky130_fd_sc_hd__a21o_1 _16876_ (.A1(_06382_),
    .A2(_06383_),
    .B1(_06385_),
    .X(_06391_));
 sky130_fd_sc_hd__o211a_1 _16877_ (.A1(_06386_),
    .A2(_06384_),
    .B1(_06381_),
    .C1(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__a21oi_1 _16878_ (.A1(_06389_),
    .A2(_06391_),
    .B1(_06381_),
    .Y(_06393_));
 sky130_fd_sc_hd__nor2_1 _16879_ (.A(_06392_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__xnor2_2 _16880_ (.A(_06380_),
    .B(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__a21o_1 _16881_ (.A1(_06088_),
    .A2(_06095_),
    .B1(_06096_),
    .X(_06396_));
 sky130_fd_sc_hd__and3_1 _16882_ (.A(_07242_),
    .B(net257),
    .C(net280),
    .X(_06397_));
 sky130_fd_sc_hd__nor2_2 _16883_ (.A(_03938_),
    .B(_04270_),
    .Y(_06399_));
 sky130_fd_sc_hd__a31oi_4 _16884_ (.A1(_07242_),
    .A2(net257),
    .A3(net280),
    .B1(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__o211ai_4 _16885_ (.A1(net261),
    .A2(_08656_),
    .B1(_04215_),
    .C1(_08700_),
    .Y(_06401_));
 sky130_fd_sc_hd__or3b_2 _16886_ (.A(_03949_),
    .B(net40),
    .C_N(net39),
    .X(_06402_));
 sky130_fd_sc_hd__o31a_1 _16887_ (.A1(_04216_),
    .A2(_08689_),
    .A3(_08667_),
    .B1(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__o21ai_1 _16888_ (.A1(_03949_),
    .A2(_04218_),
    .B1(_06401_),
    .Y(_06404_));
 sky130_fd_sc_hd__nor2_2 _16889_ (.A(_03960_),
    .B(_03737_),
    .Y(_06405_));
 sky130_fd_sc_hd__o311a_1 _16890_ (.A1(_04747_),
    .A2(net264),
    .A3(_09665_),
    .B1(net285),
    .C1(_09698_),
    .X(_06406_));
 sky130_fd_sc_hd__o211ai_2 _16891_ (.A1(net261),
    .A2(_09665_),
    .B1(net285),
    .C1(_09698_),
    .Y(_06407_));
 sky130_fd_sc_hd__o31a_1 _16892_ (.A1(_03960_),
    .A2(_04037_),
    .A3(net39),
    .B1(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__a31o_1 _16893_ (.A1(net255),
    .A2(_09698_),
    .A3(net285),
    .B1(_06405_),
    .X(_06410_));
 sky130_fd_sc_hd__o211ai_2 _16894_ (.A1(_03949_),
    .A2(_04218_),
    .B1(_06401_),
    .C1(_06407_),
    .Y(_06411_));
 sky130_fd_sc_hd__o2bb2ai_4 _16895_ (.A1_N(_06401_),
    .A2_N(_06402_),
    .B1(_06405_),
    .B2(_06406_),
    .Y(_06412_));
 sky130_fd_sc_hd__o21ai_1 _16896_ (.A1(_06405_),
    .A2(_06411_),
    .B1(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__o2111ai_1 _16897_ (.A1(_03960_),
    .A2(_03737_),
    .B1(_06400_),
    .C1(_06407_),
    .D1(_06403_),
    .Y(_06414_));
 sky130_fd_sc_hd__o22ai_1 _16898_ (.A1(_06397_),
    .A2(_06399_),
    .B1(_06404_),
    .B2(_06410_),
    .Y(_06415_));
 sky130_fd_sc_hd__o21ai_1 _16899_ (.A1(_06403_),
    .A2(_06408_),
    .B1(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__o211ai_2 _16900_ (.A1(_06403_),
    .A2(_06408_),
    .B1(_06414_),
    .C1(_06415_),
    .Y(_06417_));
 sky130_fd_sc_hd__nand2_1 _16901_ (.A(_06413_),
    .B(_06400_),
    .Y(_06418_));
 sky130_fd_sc_hd__o221ai_4 _16902_ (.A1(_06397_),
    .A2(_06399_),
    .B1(_06405_),
    .B2(_06411_),
    .C1(_06412_),
    .Y(_06419_));
 sky130_fd_sc_hd__o211ai_4 _16903_ (.A1(_06412_),
    .A2(_06400_),
    .B1(_06145_),
    .C1(_06417_),
    .Y(_06421_));
 sky130_fd_sc_hd__nand3_4 _16904_ (.A(_06418_),
    .B(_06419_),
    .C(_06144_),
    .Y(_06422_));
 sky130_fd_sc_hd__o2111ai_4 _16905_ (.A1(_06099_),
    .A2(_06094_),
    .B1(_06097_),
    .C1(_06421_),
    .D1(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__a22o_1 _16906_ (.A1(_06097_),
    .A2(_06101_),
    .B1(_06421_),
    .B2(_06422_),
    .X(_06424_));
 sky130_fd_sc_hd__a21o_1 _16907_ (.A1(_06421_),
    .A2(_06422_),
    .B1(_06396_),
    .X(_06425_));
 sky130_fd_sc_hd__o211ai_4 _16908_ (.A1(_06096_),
    .A2(_06100_),
    .B1(_06421_),
    .C1(_06422_),
    .Y(_06426_));
 sky130_fd_sc_hd__o2111ai_4 _16909_ (.A1(_06105_),
    .A2(_05749_),
    .B1(_06103_),
    .C1(_06423_),
    .D1(_06424_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand3_2 _16910_ (.A(_06425_),
    .B(_06426_),
    .C(_06110_),
    .Y(_06428_));
 sky130_fd_sc_hd__a21o_2 _16911_ (.A1(_06427_),
    .A2(_06428_),
    .B1(_06395_),
    .X(_06429_));
 sky130_fd_sc_hd__nand3_4 _16912_ (.A(_06395_),
    .B(_06427_),
    .C(_06428_),
    .Y(_06430_));
 sky130_fd_sc_hd__a31o_2 _16913_ (.A1(_06135_),
    .A2(_06171_),
    .A3(_06172_),
    .B1(_06133_),
    .X(_06432_));
 sky130_fd_sc_hd__o2bb2ai_4 _16914_ (.A1_N(_06429_),
    .A2_N(_06430_),
    .B1(_06134_),
    .B2(_06173_),
    .Y(_06433_));
 sky130_fd_sc_hd__a22oi_4 _16915_ (.A1(_06429_),
    .A2(_06430_),
    .B1(_06432_),
    .B2(_06177_),
    .Y(_06434_));
 sky130_fd_sc_hd__and4_1 _16916_ (.A(_06177_),
    .B(_06429_),
    .C(_06430_),
    .D(_06432_),
    .X(_06435_));
 sky130_fd_sc_hd__nand4_4 _16917_ (.A(_06177_),
    .B(_06429_),
    .C(_06430_),
    .D(_06432_),
    .Y(_06436_));
 sky130_fd_sc_hd__o21ai_2 _16918_ (.A1(_06084_),
    .A2(_06112_),
    .B1(_06114_),
    .Y(_06437_));
 sky130_fd_sc_hd__o21a_1 _16919_ (.A1(_06084_),
    .A2(_06112_),
    .B1(_06114_),
    .X(_06438_));
 sky130_fd_sc_hd__o21ai_4 _16920_ (.A1(_06434_),
    .A2(_06435_),
    .B1(_06437_),
    .Y(_06439_));
 sky130_fd_sc_hd__o211ai_4 _16921_ (.A1(_06178_),
    .A2(_06433_),
    .B1(_06436_),
    .C1(_06438_),
    .Y(_06440_));
 sky130_fd_sc_hd__o21ai_1 _16922_ (.A1(_06434_),
    .A2(_06435_),
    .B1(_06438_),
    .Y(_06441_));
 sky130_fd_sc_hd__o211ai_2 _16923_ (.A1(_06178_),
    .A2(_06433_),
    .B1(_06436_),
    .C1(_06437_),
    .Y(_06443_));
 sky130_fd_sc_hd__nand2_1 _16924_ (.A(_06439_),
    .B(_06440_),
    .Y(_06444_));
 sky130_fd_sc_hd__o32a_1 _16925_ (.A1(_04353_),
    .A2(net205),
    .A3(_05932_),
    .B1(_04375_),
    .B2(_04157_),
    .X(_06445_));
 sky130_fd_sc_hd__o32ai_4 _16926_ (.A1(_04353_),
    .A2(net205),
    .A3(_05932_),
    .B1(_04375_),
    .B2(_04157_),
    .Y(_06446_));
 sky130_fd_sc_hd__nor2_1 _16927_ (.A(_04168_),
    .B(_04331_),
    .Y(_06447_));
 sky130_fd_sc_hd__or3_2 _16928_ (.A(net44),
    .B(_04168_),
    .C(_03286_),
    .X(_06448_));
 sky130_fd_sc_hd__o31ai_4 _16929_ (.A1(net17),
    .A2(net245),
    .A3(net241),
    .B1(net18),
    .Y(_06449_));
 sky130_fd_sc_hd__nor2_2 _16930_ (.A(net17),
    .B(net18),
    .Y(_06450_));
 sky130_fd_sc_hd__or2_4 _16931_ (.A(net17),
    .B(net18),
    .X(_06451_));
 sky130_fd_sc_hd__nand4_4 _16932_ (.A(_06519_),
    .B(_03955_),
    .C(_05926_),
    .D(_06450_),
    .Y(_06452_));
 sky130_fd_sc_hd__o21ai_4 _16933_ (.A1(_05931_),
    .A2(_06451_),
    .B1(net200),
    .Y(_06454_));
 sky130_fd_sc_hd__o211ai_2 _16934_ (.A1(net175),
    .A2(_06451_),
    .B1(net33),
    .C1(net200),
    .Y(_06455_));
 sky130_fd_sc_hd__a31oi_1 _16935_ (.A1(_06219_),
    .A2(_06221_),
    .A3(_04484_),
    .B1(_06447_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand2_2 _16936_ (.A(_06456_),
    .B(_06455_),
    .Y(_06457_));
 sky130_fd_sc_hd__o2bb2ai_1 _16937_ (.A1_N(_06456_),
    .A2_N(_06455_),
    .B1(_06448_),
    .B2(net18),
    .Y(_06458_));
 sky130_fd_sc_hd__nand2_2 _16938_ (.A(_06458_),
    .B(_06445_),
    .Y(_06459_));
 sky130_fd_sc_hd__o211ai_4 _16939_ (.A1(_06448_),
    .A2(net18),
    .B1(_06446_),
    .C1(_06457_),
    .Y(_06460_));
 sky130_fd_sc_hd__o221a_1 _16940_ (.A1(_04146_),
    .A2(_04375_),
    .B1(_05554_),
    .B2(_04353_),
    .C1(_06229_),
    .X(_06461_));
 sky130_fd_sc_hd__a32oi_4 _16941_ (.A1(_06223_),
    .A2(_06224_),
    .A3(_06227_),
    .B1(_06218_),
    .B2(_06229_),
    .Y(_06462_));
 sky130_fd_sc_hd__o2bb2a_2 _16942_ (.A1_N(_06459_),
    .A2_N(_06460_),
    .B1(_06461_),
    .B2(_06230_),
    .X(_06463_));
 sky130_fd_sc_hd__o2bb2ai_4 _16943_ (.A1_N(_06459_),
    .A2_N(_06460_),
    .B1(_06461_),
    .B2(_06230_),
    .Y(_06465_));
 sky130_fd_sc_hd__nand3_4 _16944_ (.A(_06459_),
    .B(_06460_),
    .C(_06462_),
    .Y(_06466_));
 sky130_fd_sc_hd__o22a_1 _16945_ (.A1(_04113_),
    .A2(_05260_),
    .B1(_05077_),
    .B2(_05238_),
    .X(_06467_));
 sky130_fd_sc_hd__a32o_1 _16946_ (.A1(net212),
    .A2(net183),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net13),
    .X(_06468_));
 sky130_fd_sc_hd__nand3_2 _16947_ (.A(net181),
    .B(net180),
    .C(net305),
    .Y(_06469_));
 sky130_fd_sc_hd__or3b_2 _16948_ (.A(net59),
    .B(_04135_),
    .C_N(net58),
    .X(_06470_));
 sky130_fd_sc_hd__o211ai_4 _16949_ (.A1(net185),
    .A2(_05551_),
    .B1(net317),
    .C1(_05549_),
    .Y(_06471_));
 sky130_fd_sc_hd__or3b_1 _16950_ (.A(net58),
    .B(_04146_),
    .C_N(net55),
    .X(_06472_));
 sky130_fd_sc_hd__a22oi_2 _16951_ (.A1(_06469_),
    .A2(_06470_),
    .B1(_06471_),
    .B2(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__a22o_1 _16952_ (.A1(_06469_),
    .A2(_06470_),
    .B1(_06471_),
    .B2(_06472_),
    .X(_06474_));
 sky130_fd_sc_hd__o2111a_2 _16953_ (.A1(_04146_),
    .A2(net316),
    .B1(_06469_),
    .C1(_06470_),
    .D1(_06471_),
    .X(_06476_));
 sky130_fd_sc_hd__o2111ai_4 _16954_ (.A1(_04146_),
    .A2(net316),
    .B1(_06469_),
    .C1(_06470_),
    .D1(_06471_),
    .Y(_06477_));
 sky130_fd_sc_hd__a21oi_1 _16955_ (.A1(_06474_),
    .A2(_06477_),
    .B1(_06468_),
    .Y(_06478_));
 sky130_fd_sc_hd__o21ai_1 _16956_ (.A1(_06473_),
    .A2(_06476_),
    .B1(_06467_),
    .Y(_06479_));
 sky130_fd_sc_hd__and3_1 _16957_ (.A(_06468_),
    .B(_06474_),
    .C(_06477_),
    .X(_06480_));
 sky130_fd_sc_hd__nand3_1 _16958_ (.A(_06468_),
    .B(_06474_),
    .C(_06477_),
    .Y(_06481_));
 sky130_fd_sc_hd__nand3_1 _16959_ (.A(_06474_),
    .B(_06477_),
    .C(_06467_),
    .Y(_06482_));
 sky130_fd_sc_hd__o21ai_1 _16960_ (.A1(_06473_),
    .A2(_06476_),
    .B1(_06468_),
    .Y(_06483_));
 sky130_fd_sc_hd__nand2_1 _16961_ (.A(_06482_),
    .B(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__o2bb2ai_4 _16962_ (.A1_N(_06465_),
    .A2_N(_06466_),
    .B1(_06478_),
    .B2(_06480_),
    .Y(_06485_));
 sky130_fd_sc_hd__a32o_1 _16963_ (.A1(_06459_),
    .A2(_06462_),
    .A3(_06460_),
    .B1(_06483_),
    .B2(_06482_),
    .X(_06487_));
 sky130_fd_sc_hd__nand4_4 _16964_ (.A(_06465_),
    .B(_06466_),
    .C(_06479_),
    .D(_06481_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand2_2 _16965_ (.A(_06241_),
    .B(_06256_),
    .Y(_06489_));
 sky130_fd_sc_hd__a21oi_4 _16966_ (.A1(_06485_),
    .A2(_06488_),
    .B1(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__a21o_1 _16967_ (.A1(_06485_),
    .A2(_06488_),
    .B1(_06489_),
    .X(_06491_));
 sky130_fd_sc_hd__o211a_2 _16968_ (.A1(_06463_),
    .A2(_06487_),
    .B1(_06485_),
    .C1(_06489_),
    .X(_06492_));
 sky130_fd_sc_hd__o211ai_4 _16969_ (.A1(_06463_),
    .A2(_06487_),
    .B1(_06485_),
    .C1(_06489_),
    .Y(_06493_));
 sky130_fd_sc_hd__nor2_2 _16970_ (.A(_04069_),
    .B(_07691_),
    .Y(_06494_));
 sky130_fd_sc_hd__o311a_2 _16971_ (.A1(net7),
    .A2(net249),
    .A3(_04407_),
    .B1(_07658_),
    .C1(net224),
    .X(_06495_));
 sky130_fd_sc_hd__o22a_1 _16972_ (.A1(_04069_),
    .A2(_07691_),
    .B1(net187),
    .B2(_07669_),
    .X(_06496_));
 sky130_fd_sc_hd__o211ai_4 _16973_ (.A1(net232),
    .A2(_04787_),
    .B1(_05688_),
    .C1(net215),
    .Y(_06498_));
 sky130_fd_sc_hd__or3b_2 _16974_ (.A(net61),
    .B(_04091_),
    .C_N(net60),
    .X(_06499_));
 sky130_fd_sc_hd__or3b_2 _16975_ (.A(net62),
    .B(_04080_),
    .C_N(net61),
    .X(_06500_));
 sky130_fd_sc_hd__nand3_2 _16976_ (.A(net219),
    .B(_04559_),
    .C(net292),
    .Y(_06501_));
 sky130_fd_sc_hd__a22oi_4 _16977_ (.A1(_06498_),
    .A2(_06499_),
    .B1(_06500_),
    .B2(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__a22o_1 _16978_ (.A1(_06498_),
    .A2(_06499_),
    .B1(_06500_),
    .B2(_06501_),
    .X(_06503_));
 sky130_fd_sc_hd__and4_2 _16979_ (.A(_06498_),
    .B(_06499_),
    .C(_06500_),
    .D(_06501_),
    .X(_06504_));
 sky130_fd_sc_hd__o2111ai_2 _16980_ (.A1(_04091_),
    .A2(_05720_),
    .B1(_06498_),
    .C1(_06500_),
    .D1(_06501_),
    .Y(_06505_));
 sky130_fd_sc_hd__o21ai_2 _16981_ (.A1(_06502_),
    .A2(_06504_),
    .B1(_06496_),
    .Y(_06506_));
 sky130_fd_sc_hd__o21ai_2 _16982_ (.A1(_06494_),
    .A2(_06495_),
    .B1(_06503_),
    .Y(_06507_));
 sky130_fd_sc_hd__nand3_2 _16983_ (.A(_06503_),
    .B(_06505_),
    .C(_06496_),
    .Y(_06509_));
 sky130_fd_sc_hd__o22ai_4 _16984_ (.A1(_06494_),
    .A2(_06495_),
    .B1(_06502_),
    .B2(_06504_),
    .Y(_06510_));
 sky130_fd_sc_hd__a21oi_2 _16985_ (.A1(_06243_),
    .A2(_06250_),
    .B1(_06248_),
    .Y(_06511_));
 sky130_fd_sc_hd__nand4_1 _16986_ (.A(_06249_),
    .B(_06255_),
    .C(_06509_),
    .D(_06510_),
    .Y(_06512_));
 sky130_fd_sc_hd__o221a_2 _16987_ (.A1(_06248_),
    .A2(_06253_),
    .B1(_06504_),
    .B2(_06507_),
    .C1(_06506_),
    .X(_06513_));
 sky130_fd_sc_hd__o221ai_4 _16988_ (.A1(_06248_),
    .A2(_06253_),
    .B1(_06504_),
    .B2(_06507_),
    .C1(_06506_),
    .Y(_06514_));
 sky130_fd_sc_hd__a31o_2 _16989_ (.A1(_06511_),
    .A2(_06510_),
    .A3(_06509_),
    .B1(_06199_),
    .X(_06515_));
 sky130_fd_sc_hd__a21o_1 _16990_ (.A1(_06512_),
    .A2(_06514_),
    .B1(_06198_),
    .X(_06516_));
 sky130_fd_sc_hd__o21ai_4 _16991_ (.A1(_06513_),
    .A2(_06515_),
    .B1(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__nand3_4 _16992_ (.A(_06491_),
    .B(_06493_),
    .C(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__o21bai_4 _16993_ (.A1(_06490_),
    .A2(_06492_),
    .B1_N(_06517_),
    .Y(_06520_));
 sky130_fd_sc_hd__o21ai_4 _16994_ (.A1(_06490_),
    .A2(_06492_),
    .B1(_06517_),
    .Y(_06521_));
 sky130_fd_sc_hd__o2111ai_4 _16995_ (.A1(_06513_),
    .A2(_06515_),
    .B1(_06516_),
    .C1(_06493_),
    .D1(_06491_),
    .Y(_06522_));
 sky130_fd_sc_hd__o211a_1 _16996_ (.A1(_06260_),
    .A2(_06266_),
    .B1(_06518_),
    .C1(_06520_),
    .X(_06523_));
 sky130_fd_sc_hd__o211ai_4 _16997_ (.A1(_06260_),
    .A2(_06266_),
    .B1(_06518_),
    .C1(_06520_),
    .Y(_06524_));
 sky130_fd_sc_hd__nand3_4 _16998_ (.A(_06521_),
    .B(_06522_),
    .C(_06267_),
    .Y(_06525_));
 sky130_fd_sc_hd__o32a_2 _16999_ (.A1(_06149_),
    .A2(_06162_),
    .A3(_06163_),
    .B1(_06147_),
    .B2(_06166_),
    .X(_06526_));
 sky130_fd_sc_hd__a31oi_4 _17000_ (.A1(_05908_),
    .A2(_06200_),
    .A3(_06201_),
    .B1(_06184_),
    .Y(_06527_));
 sky130_fd_sc_hd__a32o_2 _17001_ (.A1(_05908_),
    .A2(_06200_),
    .A3(_06201_),
    .B1(_06206_),
    .B2(_06184_),
    .X(_06528_));
 sky130_fd_sc_hd__o32a_2 _17002_ (.A1(_02869_),
    .A2(_11420_),
    .A3(_11343_),
    .B1(_03982_),
    .B2(_02891_),
    .X(_06529_));
 sky130_fd_sc_hd__o211ai_2 _17003_ (.A1(_11387_),
    .A2(_12988_),
    .B1(_01293_),
    .C1(net235),
    .Y(_06531_));
 sky130_fd_sc_hd__or3b_1 _17004_ (.A(_04004_),
    .B(net37),
    .C_N(net36),
    .X(_06532_));
 sky130_fd_sc_hd__or3_1 _17005_ (.A(net36),
    .B(_04015_),
    .C(_03993_),
    .X(_06533_));
 sky130_fd_sc_hd__o211ai_2 _17006_ (.A1(net254),
    .A2(_00646_),
    .B1(_12330_),
    .C1(_00625_),
    .Y(_06534_));
 sky130_fd_sc_hd__a22oi_2 _17007_ (.A1(_06531_),
    .A2(_06532_),
    .B1(_06533_),
    .B2(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__a22o_1 _17008_ (.A1(_06531_),
    .A2(_06532_),
    .B1(_06533_),
    .B2(_06534_),
    .X(_06536_));
 sky130_fd_sc_hd__o2111a_1 _17009_ (.A1(_04015_),
    .A2(_12363_),
    .B1(_06531_),
    .C1(_06532_),
    .D1(_06534_),
    .X(_06537_));
 sky130_fd_sc_hd__o21a_1 _17010_ (.A1(_06535_),
    .A2(_06537_),
    .B1(_06529_),
    .X(_06538_));
 sky130_fd_sc_hd__nor3_2 _17011_ (.A(_06529_),
    .B(_06535_),
    .C(_06537_),
    .Y(_06539_));
 sky130_fd_sc_hd__nor2_1 _17012_ (.A(_06538_),
    .B(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__a21oi_2 _17013_ (.A1(_06150_),
    .A2(_06161_),
    .B1(_06157_),
    .Y(_06542_));
 sky130_fd_sc_hd__and3_1 _17014_ (.A(_03993_),
    .B(net6),
    .C(net34),
    .X(_06543_));
 sky130_fd_sc_hd__o311a_1 _17015_ (.A1(net263),
    .A2(_11387_),
    .A3(_02442_),
    .B1(net252),
    .C1(_02421_),
    .X(_06544_));
 sky130_fd_sc_hd__a31o_1 _17016_ (.A1(_02421_),
    .A2(net249),
    .A3(net252),
    .B1(_06543_),
    .X(_06545_));
 sky130_fd_sc_hd__nand3_2 _17017_ (.A(_04132_),
    .B(net291),
    .C(net230),
    .Y(_06546_));
 sky130_fd_sc_hd__or3b_1 _17018_ (.A(net64),
    .B(_04059_),
    .C_N(net63),
    .X(_06547_));
 sky130_fd_sc_hd__and3_1 _17019_ (.A(_03971_),
    .B(net7),
    .C(net64),
    .X(_06548_));
 sky130_fd_sc_hd__o21a_1 _17020_ (.A1(net263),
    .A2(net246),
    .B1(net289),
    .X(_06549_));
 sky130_fd_sc_hd__o311a_1 _17021_ (.A1(net263),
    .A2(_11387_),
    .A3(_03954_),
    .B1(net289),
    .C1(_03952_),
    .X(_06550_));
 sky130_fd_sc_hd__a22oi_4 _17022_ (.A1(net7),
    .A2(_10335_),
    .B1(_06549_),
    .B2(_03952_),
    .Y(_06551_));
 sky130_fd_sc_hd__o211ai_4 _17023_ (.A1(_04059_),
    .A2(_08283_),
    .B1(_06546_),
    .C1(_06551_),
    .Y(_06553_));
 sky130_fd_sc_hd__a21oi_2 _17024_ (.A1(_06546_),
    .A2(_06547_),
    .B1(_06551_),
    .Y(_06554_));
 sky130_fd_sc_hd__o2bb2ai_2 _17025_ (.A1_N(_06546_),
    .A2_N(_06547_),
    .B1(_06548_),
    .B2(_06550_),
    .Y(_06555_));
 sky130_fd_sc_hd__o211a_2 _17026_ (.A1(_06543_),
    .A2(_06544_),
    .B1(_06553_),
    .C1(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__o211ai_2 _17027_ (.A1(_06543_),
    .A2(_06544_),
    .B1(_06553_),
    .C1(_06555_),
    .Y(_06557_));
 sky130_fd_sc_hd__a21oi_2 _17028_ (.A1(_06553_),
    .A2(_06555_),
    .B1(_06545_),
    .Y(_06558_));
 sky130_fd_sc_hd__a21o_1 _17029_ (.A1(_06553_),
    .A2(_06555_),
    .B1(_06545_),
    .X(_06559_));
 sky130_fd_sc_hd__o211a_1 _17030_ (.A1(_06157_),
    .A2(_06162_),
    .B1(_06557_),
    .C1(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__o211ai_4 _17031_ (.A1(_06157_),
    .A2(_06162_),
    .B1(_06557_),
    .C1(_06559_),
    .Y(_06561_));
 sky130_fd_sc_hd__o21ai_4 _17032_ (.A1(_06556_),
    .A2(_06558_),
    .B1(_06542_),
    .Y(_06562_));
 sky130_fd_sc_hd__nand2_1 _17033_ (.A(_06561_),
    .B(_06562_),
    .Y(_06564_));
 sky130_fd_sc_hd__o211ai_4 _17034_ (.A1(_06538_),
    .A2(_06539_),
    .B1(_06561_),
    .C1(_06562_),
    .Y(_06565_));
 sky130_fd_sc_hd__nand2_2 _17035_ (.A(_06564_),
    .B(_06540_),
    .Y(_06566_));
 sky130_fd_sc_hd__nand2_2 _17036_ (.A(_06562_),
    .B(_06540_),
    .Y(_06567_));
 sky130_fd_sc_hd__a21o_1 _17037_ (.A1(_06561_),
    .A2(_06562_),
    .B1(_06540_),
    .X(_06568_));
 sky130_fd_sc_hd__o221a_1 _17038_ (.A1(_06205_),
    .A2(_06527_),
    .B1(_06560_),
    .B2(_06567_),
    .C1(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__o221ai_4 _17039_ (.A1(_06205_),
    .A2(_06527_),
    .B1(_06560_),
    .B2(_06567_),
    .C1(_06568_),
    .Y(_06570_));
 sky130_fd_sc_hd__nand3_2 _17040_ (.A(_06528_),
    .B(_06565_),
    .C(_06566_),
    .Y(_06571_));
 sky130_fd_sc_hd__nand2_1 _17041_ (.A(_06570_),
    .B(_06571_),
    .Y(_06572_));
 sky130_fd_sc_hd__a21oi_1 _17042_ (.A1(_06570_),
    .A2(_06571_),
    .B1(_06526_),
    .Y(_06573_));
 sky130_fd_sc_hd__and3_1 _17043_ (.A(_06571_),
    .B(_06526_),
    .C(_06570_),
    .X(_06575_));
 sky130_fd_sc_hd__o211a_1 _17044_ (.A1(_06166_),
    .A2(_06147_),
    .B1(_06165_),
    .C1(_06572_),
    .X(_06576_));
 sky130_fd_sc_hd__nand2_2 _17045_ (.A(_06572_),
    .B(_06526_),
    .Y(_06577_));
 sky130_fd_sc_hd__a31o_1 _17046_ (.A1(_06528_),
    .A2(_06565_),
    .A3(_06566_),
    .B1(_06526_),
    .X(_06578_));
 sky130_fd_sc_hd__o211a_1 _17047_ (.A1(_06164_),
    .A2(_06168_),
    .B1(_06570_),
    .C1(_06571_),
    .X(_06579_));
 sky130_fd_sc_hd__o211ai_2 _17048_ (.A1(_06164_),
    .A2(_06168_),
    .B1(_06570_),
    .C1(_06571_),
    .Y(_06580_));
 sky130_fd_sc_hd__o21ai_1 _17049_ (.A1(_06569_),
    .A2(_06578_),
    .B1(_06577_),
    .Y(_06581_));
 sky130_fd_sc_hd__o2111ai_4 _17050_ (.A1(_06569_),
    .A2(_06578_),
    .B1(_06577_),
    .C1(_06524_),
    .D1(_06525_),
    .Y(_06582_));
 sky130_fd_sc_hd__o2bb2ai_2 _17051_ (.A1_N(_06524_),
    .A2_N(_06525_),
    .B1(_06576_),
    .B2(_06579_),
    .Y(_06583_));
 sky130_fd_sc_hd__o211ai_4 _17052_ (.A1(_06576_),
    .A2(_06579_),
    .B1(_06524_),
    .C1(_06525_),
    .Y(_06584_));
 sky130_fd_sc_hd__o2bb2ai_4 _17053_ (.A1_N(_06524_),
    .A2_N(_06525_),
    .B1(_06573_),
    .B2(_06575_),
    .Y(_06586_));
 sky130_fd_sc_hd__a21oi_2 _17054_ (.A1(_06275_),
    .A2(_06183_),
    .B1(_06273_),
    .Y(_06587_));
 sky130_fd_sc_hd__nand3_2 _17055_ (.A(_06584_),
    .B(_06587_),
    .C(_06586_),
    .Y(_06588_));
 sky130_fd_sc_hd__o211a_2 _17056_ (.A1(_06273_),
    .A2(_06276_),
    .B1(_06582_),
    .C1(_06583_),
    .X(_06589_));
 sky130_fd_sc_hd__o211ai_4 _17057_ (.A1(_06273_),
    .A2(_06276_),
    .B1(_06582_),
    .C1(_06583_),
    .Y(_06590_));
 sky130_fd_sc_hd__nand4_2 _17058_ (.A(_06439_),
    .B(_06440_),
    .C(_06588_),
    .D(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__a22o_1 _17059_ (.A1(_06439_),
    .A2(_06440_),
    .B1(_06588_),
    .B2(_06590_),
    .X(_06592_));
 sky130_fd_sc_hd__a32oi_4 _17060_ (.A1(_06584_),
    .A2(_06587_),
    .A3(_06586_),
    .B1(_06439_),
    .B2(_06440_),
    .Y(_06593_));
 sky130_fd_sc_hd__a32o_1 _17061_ (.A1(_06584_),
    .A2(_06587_),
    .A3(_06586_),
    .B1(_06439_),
    .B2(_06440_),
    .X(_06594_));
 sky130_fd_sc_hd__a22o_1 _17062_ (.A1(_06441_),
    .A2(_06443_),
    .B1(_06588_),
    .B2(_06590_),
    .X(_06595_));
 sky130_fd_sc_hd__o211ai_4 _17063_ (.A1(_06589_),
    .A2(_06594_),
    .B1(_06359_),
    .C1(_06595_),
    .Y(_06597_));
 sky130_fd_sc_hd__o2111ai_4 _17064_ (.A1(_06282_),
    .A2(_06131_),
    .B1(_06281_),
    .C1(_06591_),
    .D1(_06592_),
    .Y(_06598_));
 sky130_fd_sc_hd__nand3_1 _17065_ (.A(_06358_),
    .B(_06597_),
    .C(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__a21o_1 _17066_ (.A1(_06597_),
    .A2(_06598_),
    .B1(_06358_),
    .X(_06600_));
 sky130_fd_sc_hd__nand2_1 _17067_ (.A(_06357_),
    .B(_06598_),
    .Y(_06601_));
 sky130_fd_sc_hd__and3_1 _17068_ (.A(_06357_),
    .B(_06597_),
    .C(_06598_),
    .X(_06602_));
 sky130_fd_sc_hd__nand3_1 _17069_ (.A(_06357_),
    .B(_06597_),
    .C(_06598_),
    .Y(_06603_));
 sky130_fd_sc_hd__a21o_1 _17070_ (.A1(_06597_),
    .A2(_06598_),
    .B1(_06357_),
    .X(_06604_));
 sky130_fd_sc_hd__nand2_1 _17071_ (.A(_06323_),
    .B(_06604_),
    .Y(_06605_));
 sky130_fd_sc_hd__nand3_1 _17072_ (.A(_06323_),
    .B(_06603_),
    .C(_06604_),
    .Y(_06606_));
 sky130_fd_sc_hd__o211ai_4 _17073_ (.A1(_06291_),
    .A2(_06322_),
    .B1(_06599_),
    .C1(_06600_),
    .Y(_06608_));
 sky130_fd_sc_hd__o211ai_2 _17074_ (.A1(_06602_),
    .A2(_06605_),
    .B1(_06608_),
    .C1(_06043_),
    .Y(_06609_));
 sky130_fd_sc_hd__a21o_1 _17075_ (.A1(_06606_),
    .A2(_06608_),
    .B1(_06043_),
    .X(_06610_));
 sky130_fd_sc_hd__a21bo_1 _17076_ (.A1(_06606_),
    .A2(_06608_),
    .B1_N(_06043_),
    .X(_06611_));
 sky130_fd_sc_hd__nand3b_1 _17077_ (.A_N(_06043_),
    .B(_06606_),
    .C(_06608_),
    .Y(_06612_));
 sky130_fd_sc_hd__and3_1 _17078_ (.A(_06321_),
    .B(_06611_),
    .C(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__nand3_2 _17079_ (.A(_06321_),
    .B(_06611_),
    .C(_06612_),
    .Y(_06614_));
 sky130_fd_sc_hd__o211a_1 _17080_ (.A1(_06297_),
    .A2(_06302_),
    .B1(_06609_),
    .C1(_06610_),
    .X(_06615_));
 sky130_fd_sc_hd__o211ai_4 _17081_ (.A1(_06297_),
    .A2(_06302_),
    .B1(_06609_),
    .C1(_06610_),
    .Y(_06616_));
 sky130_fd_sc_hd__a32oi_4 _17082_ (.A1(_06300_),
    .A2(_06304_),
    .A3(_06305_),
    .B1(_06614_),
    .B2(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__o2111a_1 _17083_ (.A1(_06303_),
    .A2(_06297_),
    .B1(_06300_),
    .C1(_06305_),
    .D1(_06616_),
    .X(_06619_));
 sky130_fd_sc_hd__o2111ai_1 _17084_ (.A1(_06303_),
    .A2(_06297_),
    .B1(_06300_),
    .C1(_06305_),
    .D1(_06616_),
    .Y(_06620_));
 sky130_fd_sc_hd__a21oi_2 _17085_ (.A1(_06619_),
    .A2(_06614_),
    .B1(_06617_),
    .Y(_06621_));
 sky130_fd_sc_hd__o2bb2a_1 _17086_ (.A1_N(_06016_),
    .A2_N(_06306_),
    .B1(_06308_),
    .B2(_06319_),
    .X(_06622_));
 sky130_fd_sc_hd__xnor2_1 _17087_ (.A(_06621_),
    .B(_06622_),
    .Y(net82));
 sky130_fd_sc_hd__o31a_1 _17088_ (.A1(_05716_),
    .A2(_06040_),
    .A3(_06353_),
    .B1(_06351_),
    .X(_06623_));
 sky130_fd_sc_hd__nand2_2 _17089_ (.A(_06358_),
    .B(_06597_),
    .Y(_06624_));
 sky130_fd_sc_hd__nand2_1 _17090_ (.A(_06598_),
    .B(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__a21oi_2 _17091_ (.A1(_06444_),
    .A2(_06588_),
    .B1(_06589_),
    .Y(_06626_));
 sky130_fd_sc_hd__nand2_1 _17092_ (.A(_06428_),
    .B(_06430_),
    .Y(_06627_));
 sky130_fd_sc_hd__a32oi_4 _17093_ (.A1(_06528_),
    .A2(_06565_),
    .A3(_06566_),
    .B1(_06570_),
    .B2(_06526_),
    .Y(_06629_));
 sky130_fd_sc_hd__or3b_1 _17094_ (.A(_03916_),
    .B(net43),
    .C_N(net42),
    .X(_06630_));
 sky130_fd_sc_hd__o211ai_2 _17095_ (.A1(_04747_),
    .A2(net264),
    .B1(net243),
    .C1(_06486_),
    .Y(_06631_));
 sky130_fd_sc_hd__or3b_1 _17096_ (.A(_03938_),
    .B(net42),
    .C_N(net41),
    .X(_06632_));
 sky130_fd_sc_hd__nand3_1 _17097_ (.A(_07242_),
    .B(net257),
    .C(net279),
    .Y(_06633_));
 sky130_fd_sc_hd__a22oi_2 _17098_ (.A1(_06630_),
    .A2(_06631_),
    .B1(_06632_),
    .B2(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__o2111a_1 _17099_ (.A1(_03916_),
    .A2(_04898_),
    .B1(_06631_),
    .C1(_06632_),
    .D1(_06633_),
    .X(_06635_));
 sky130_fd_sc_hd__o2111ai_1 _17100_ (.A1(_03916_),
    .A2(_04898_),
    .B1(_06631_),
    .C1(_06632_),
    .D1(_06633_),
    .Y(_06636_));
 sky130_fd_sc_hd__a32o_1 _17101_ (.A1(_05841_),
    .A2(net265),
    .A3(_04985_),
    .B1(_04988_),
    .B2(net29),
    .X(_06637_));
 sky130_fd_sc_hd__nand3b_1 _17102_ (.A_N(_06634_),
    .B(_06636_),
    .C(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__o21bai_1 _17103_ (.A1(_06634_),
    .A2(_06635_),
    .B1_N(_06637_),
    .Y(_06640_));
 sky130_fd_sc_hd__o221a_1 _17104_ (.A1(_05457_),
    .A2(_04986_),
    .B1(_04989_),
    .B2(_03725_),
    .C1(_06370_),
    .X(_06641_));
 sky130_fd_sc_hd__nand2_1 _17105_ (.A(_06362_),
    .B(_06370_),
    .Y(_06642_));
 sky130_fd_sc_hd__o2bb2ai_1 _17106_ (.A1_N(_06638_),
    .A2_N(_06640_),
    .B1(_06641_),
    .B2(_06371_),
    .Y(_06643_));
 sky130_fd_sc_hd__nand4_2 _17107_ (.A(_06372_),
    .B(_06638_),
    .C(_06640_),
    .D(_06642_),
    .Y(_06644_));
 sky130_fd_sc_hd__o32a_1 _17108_ (.A1(_05763_),
    .A2(net306),
    .A3(_04703_),
    .B1(_03506_),
    .B2(_05766_),
    .X(_06645_));
 sky130_fd_sc_hd__a32o_1 _17109_ (.A1(net313),
    .A2(_04747_),
    .A3(net275),
    .B1(_05765_),
    .B2(net26),
    .X(_06646_));
 sky130_fd_sc_hd__or3b_1 _17110_ (.A(_03616_),
    .B(net47),
    .C_N(net46),
    .X(_06647_));
 sky130_fd_sc_hd__nand3_1 _17111_ (.A(net266),
    .B(net302),
    .C(_05462_),
    .Y(_06648_));
 sky130_fd_sc_hd__or3_1 _17112_ (.A(net46),
    .B(_04124_),
    .C(_03725_),
    .X(_06649_));
 sky130_fd_sc_hd__o211ai_2 _17113_ (.A1(_04747_),
    .A2(_05436_),
    .B1(net276),
    .C1(_05414_),
    .Y(_06651_));
 sky130_fd_sc_hd__a22oi_2 _17114_ (.A1(_06647_),
    .A2(_06648_),
    .B1(_06649_),
    .B2(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__o2111a_1 _17115_ (.A1(_03616_),
    .A2(_05465_),
    .B1(_06648_),
    .C1(_06649_),
    .D1(_06651_),
    .X(_06653_));
 sky130_fd_sc_hd__o2111ai_1 _17116_ (.A1(_03616_),
    .A2(_05465_),
    .B1(_06648_),
    .C1(_06649_),
    .D1(_06651_),
    .Y(_06654_));
 sky130_fd_sc_hd__o21a_1 _17117_ (.A1(_06652_),
    .A2(_06653_),
    .B1(_06645_),
    .X(_06655_));
 sky130_fd_sc_hd__nor3_1 _17118_ (.A(_06645_),
    .B(_06652_),
    .C(_06653_),
    .Y(_06656_));
 sky130_fd_sc_hd__nor2_1 _17119_ (.A(_06655_),
    .B(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__a21oi_1 _17120_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__nand3_1 _17121_ (.A(_06643_),
    .B(_06644_),
    .C(_06657_),
    .Y(_06659_));
 sky130_fd_sc_hd__and2b_1 _17122_ (.A_N(_06658_),
    .B(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__o21ai_1 _17123_ (.A1(_06529_),
    .A2(_06537_),
    .B1(_06536_),
    .Y(_06662_));
 sky130_fd_sc_hd__o21a_1 _17124_ (.A1(_06529_),
    .A2(_06537_),
    .B1(_06536_),
    .X(_06663_));
 sky130_fd_sc_hd__o32a_1 _17125_ (.A1(_04268_),
    .A2(_08689_),
    .A3(_08667_),
    .B1(_03949_),
    .B2(_04270_),
    .X(_06664_));
 sky130_fd_sc_hd__o211ai_2 _17126_ (.A1(net261),
    .A2(_09665_),
    .B1(_04215_),
    .C1(_09698_),
    .Y(_06665_));
 sky130_fd_sc_hd__or3b_1 _17127_ (.A(_03960_),
    .B(net40),
    .C_N(net39),
    .X(_06666_));
 sky130_fd_sc_hd__o211ai_2 _17128_ (.A1(net261),
    .A2(_11387_),
    .B1(net285),
    .C1(_11354_),
    .Y(_06667_));
 sky130_fd_sc_hd__or3_1 _17129_ (.A(net39),
    .B(_04037_),
    .C(_03982_),
    .X(_06668_));
 sky130_fd_sc_hd__a22oi_1 _17130_ (.A1(_06665_),
    .A2(_06666_),
    .B1(_06667_),
    .B2(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__a22o_1 _17131_ (.A1(_06665_),
    .A2(_06666_),
    .B1(_06667_),
    .B2(_06668_),
    .X(_06670_));
 sky130_fd_sc_hd__and4_1 _17132_ (.A(_06665_),
    .B(_06666_),
    .C(_06667_),
    .D(_06668_),
    .X(_06671_));
 sky130_fd_sc_hd__nand4_1 _17133_ (.A(_06665_),
    .B(_06666_),
    .C(_06667_),
    .D(_06668_),
    .Y(_06673_));
 sky130_fd_sc_hd__o21ai_1 _17134_ (.A1(_06669_),
    .A2(_06671_),
    .B1(_06664_),
    .Y(_06674_));
 sky130_fd_sc_hd__nand3b_1 _17135_ (.A_N(_06664_),
    .B(_06670_),
    .C(_06673_),
    .Y(_06675_));
 sky130_fd_sc_hd__o21bai_1 _17136_ (.A1(_06669_),
    .A2(_06671_),
    .B1_N(_06664_),
    .Y(_06676_));
 sky130_fd_sc_hd__nand3_1 _17137_ (.A(_06670_),
    .B(_06673_),
    .C(_06664_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand3_1 _17138_ (.A(_06663_),
    .B(_06676_),
    .C(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__nand3_2 _17139_ (.A(_06674_),
    .B(_06675_),
    .C(_06662_),
    .Y(_06679_));
 sky130_fd_sc_hd__a21oi_1 _17140_ (.A1(_06678_),
    .A2(_06679_),
    .B1(_06416_),
    .Y(_06680_));
 sky130_fd_sc_hd__a21o_1 _17141_ (.A1(_06678_),
    .A2(_06679_),
    .B1(_06416_),
    .X(_06681_));
 sky130_fd_sc_hd__and3_1 _17142_ (.A(_06678_),
    .B(_06679_),
    .C(_06416_),
    .X(_06682_));
 sky130_fd_sc_hd__nand3_1 _17143_ (.A(_06678_),
    .B(_06679_),
    .C(_06416_),
    .Y(_06684_));
 sky130_fd_sc_hd__nand2_1 _17144_ (.A(_06422_),
    .B(_06426_),
    .Y(_06685_));
 sky130_fd_sc_hd__a21oi_1 _17145_ (.A1(_06681_),
    .A2(_06684_),
    .B1(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__a21o_1 _17146_ (.A1(_06681_),
    .A2(_06684_),
    .B1(_06685_),
    .X(_06687_));
 sky130_fd_sc_hd__a211oi_1 _17147_ (.A1(_06422_),
    .A2(_06426_),
    .B1(_06680_),
    .C1(_06682_),
    .Y(_06688_));
 sky130_fd_sc_hd__a211o_1 _17148_ (.A1(_06422_),
    .A2(_06426_),
    .B1(_06680_),
    .C1(_06682_),
    .X(_06689_));
 sky130_fd_sc_hd__o21bai_2 _17149_ (.A1(_06686_),
    .A2(_06688_),
    .B1_N(_06660_),
    .Y(_06690_));
 sky130_fd_sc_hd__nand3_1 _17150_ (.A(_06689_),
    .B(_06660_),
    .C(_06687_),
    .Y(_06691_));
 sky130_fd_sc_hd__a21oi_1 _17151_ (.A1(_06690_),
    .A2(_06691_),
    .B1(_06629_),
    .Y(_06692_));
 sky130_fd_sc_hd__a21o_1 _17152_ (.A1(_06690_),
    .A2(_06691_),
    .B1(_06629_),
    .X(_06693_));
 sky130_fd_sc_hd__nand3_2 _17153_ (.A(_06629_),
    .B(_06690_),
    .C(_06691_),
    .Y(_06695_));
 sky130_fd_sc_hd__inv_2 _17154_ (.A(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__a21oi_1 _17155_ (.A1(_06693_),
    .A2(_06695_),
    .B1(_06627_),
    .Y(_06697_));
 sky130_fd_sc_hd__a21o_1 _17156_ (.A1(_06693_),
    .A2(_06695_),
    .B1(_06627_),
    .X(_06698_));
 sky130_fd_sc_hd__a21oi_1 _17157_ (.A1(_06428_),
    .A2(_06430_),
    .B1(_06692_),
    .Y(_06699_));
 sky130_fd_sc_hd__a211o_1 _17158_ (.A1(_06428_),
    .A2(_06430_),
    .B1(_06692_),
    .C1(_06696_),
    .X(_06700_));
 sky130_fd_sc_hd__a21o_1 _17159_ (.A1(_06695_),
    .A2(_06699_),
    .B1(_06697_),
    .X(_06701_));
 sky130_fd_sc_hd__a32oi_4 _17160_ (.A1(_06521_),
    .A2(_06522_),
    .A3(_06267_),
    .B1(_06577_),
    .B2(_06580_),
    .Y(_06702_));
 sky130_fd_sc_hd__a32oi_4 _17161_ (.A1(_06268_),
    .A2(_06518_),
    .A3(_06520_),
    .B1(_06525_),
    .B2(_06581_),
    .Y(_06703_));
 sky130_fd_sc_hd__o21ai_4 _17162_ (.A1(_06517_),
    .A2(_06490_),
    .B1(_06493_),
    .Y(_06704_));
 sky130_fd_sc_hd__o21a_1 _17163_ (.A1(_06517_),
    .A2(_06490_),
    .B1(_06493_),
    .X(_06706_));
 sky130_fd_sc_hd__a32o_1 _17164_ (.A1(net219),
    .A2(_04559_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net10),
    .X(_06707_));
 sky130_fd_sc_hd__o211ai_4 _17165_ (.A1(_04787_),
    .A2(net208),
    .B1(_05688_),
    .C1(net212),
    .Y(_06708_));
 sky130_fd_sc_hd__or3b_2 _17166_ (.A(net61),
    .B(_04113_),
    .C_N(net60),
    .X(_06709_));
 sky130_fd_sc_hd__o221ai_4 _17167_ (.A1(net232),
    .A2(_04787_),
    .B1(_04091_),
    .B2(_04558_),
    .C1(net292),
    .Y(_06710_));
 sky130_fd_sc_hd__or3b_2 _17168_ (.A(net62),
    .B(_04091_),
    .C_N(net61),
    .X(_06711_));
 sky130_fd_sc_hd__a22oi_4 _17169_ (.A1(_06708_),
    .A2(_06709_),
    .B1(_06710_),
    .B2(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__a22o_1 _17170_ (.A1(_06708_),
    .A2(_06709_),
    .B1(_06710_),
    .B2(_06711_),
    .X(_06713_));
 sky130_fd_sc_hd__o2111a_1 _17171_ (.A1(_04091_),
    .A2(_06859_),
    .B1(_06708_),
    .C1(_06709_),
    .D1(_06710_),
    .X(_06714_));
 sky130_fd_sc_hd__o2111ai_2 _17172_ (.A1(_04091_),
    .A2(_06859_),
    .B1(_06708_),
    .C1(_06709_),
    .D1(_06710_),
    .Y(_06715_));
 sky130_fd_sc_hd__o21bai_2 _17173_ (.A1(_06712_),
    .A2(_06714_),
    .B1_N(_06707_),
    .Y(_06717_));
 sky130_fd_sc_hd__and3_2 _17174_ (.A(_06707_),
    .B(_06713_),
    .C(_06715_),
    .X(_06718_));
 sky130_fd_sc_hd__nand3_1 _17175_ (.A(_06707_),
    .B(_06713_),
    .C(_06715_),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_1 _17176_ (.A(_06717_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__nor2_1 _17177_ (.A(_06468_),
    .B(_06473_),
    .Y(_06721_));
 sky130_fd_sc_hd__o21ai_1 _17178_ (.A1(_06467_),
    .A2(_06476_),
    .B1(_06474_),
    .Y(_06722_));
 sky130_fd_sc_hd__a21oi_1 _17179_ (.A1(_06468_),
    .A2(_06477_),
    .B1(_06473_),
    .Y(_06723_));
 sky130_fd_sc_hd__o2bb2ai_2 _17180_ (.A1_N(_06717_),
    .A2_N(_06719_),
    .B1(_06721_),
    .B2(_06476_),
    .Y(_06724_));
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(_06722_),
    .B(_06717_),
    .Y(_06725_));
 sky130_fd_sc_hd__nand3_1 _17182_ (.A(_06722_),
    .B(_06719_),
    .C(_06717_),
    .Y(_06726_));
 sky130_fd_sc_hd__o31a_2 _17183_ (.A1(_06494_),
    .A2(_06495_),
    .A3(_06502_),
    .B1(_06505_),
    .X(_06728_));
 sky130_fd_sc_hd__a21oi_1 _17184_ (.A1(_06724_),
    .A2(_06726_),
    .B1(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__a21o_1 _17185_ (.A1(_06724_),
    .A2(_06726_),
    .B1(_06728_),
    .X(_06730_));
 sky130_fd_sc_hd__a21boi_2 _17186_ (.A1(_06720_),
    .A2(_06723_),
    .B1_N(_06728_),
    .Y(_06731_));
 sky130_fd_sc_hd__o21ai_2 _17187_ (.A1(_06718_),
    .A2(_06725_),
    .B1(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__a21oi_2 _17188_ (.A1(_06726_),
    .A2(_06731_),
    .B1(_06729_),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_1 _17189_ (.A(_06730_),
    .B(_06732_),
    .Y(_06734_));
 sky130_fd_sc_hd__a21boi_1 _17190_ (.A1(_06484_),
    .A2(_06465_),
    .B1_N(_06466_),
    .Y(_06735_));
 sky130_fd_sc_hd__nand2_1 _17191_ (.A(_06466_),
    .B(_06488_),
    .Y(_06736_));
 sky130_fd_sc_hd__nor2_1 _17192_ (.A(_04135_),
    .B(_05260_),
    .Y(_06737_));
 sky130_fd_sc_hd__and3_1 _17193_ (.A(net181),
    .B(net180),
    .C(_05227_),
    .X(_06739_));
 sky130_fd_sc_hd__o22a_1 _17194_ (.A1(_04135_),
    .A2(_05260_),
    .B1(_05294_),
    .B2(_05238_),
    .X(_06740_));
 sky130_fd_sc_hd__or3b_1 _17195_ (.A(net58),
    .B(_04157_),
    .C_N(net55),
    .X(_06741_));
 sky130_fd_sc_hd__o221ai_4 _17196_ (.A1(net232),
    .A2(_05927_),
    .B1(_04157_),
    .B2(_05552_),
    .C1(_04627_),
    .Y(_06742_));
 sky130_fd_sc_hd__a211oi_2 _17197_ (.A1(_04788_),
    .A2(_05550_),
    .B1(_04900_),
    .C1(_05548_),
    .Y(_06743_));
 sky130_fd_sc_hd__o211ai_2 _17198_ (.A1(net185),
    .A2(_05551_),
    .B1(_04889_),
    .C1(_05549_),
    .Y(_06744_));
 sky130_fd_sc_hd__and3b_1 _17199_ (.A_N(net59),
    .B(net15),
    .C(net58),
    .X(_06745_));
 sky130_fd_sc_hd__or3b_1 _17200_ (.A(net59),
    .B(_04146_),
    .C_N(net58),
    .X(_06746_));
 sky130_fd_sc_hd__o2111a_1 _17201_ (.A1(_04157_),
    .A2(net316),
    .B1(_06742_),
    .C1(_06744_),
    .D1(_06746_),
    .X(_06747_));
 sky130_fd_sc_hd__o2111ai_4 _17202_ (.A1(_04157_),
    .A2(net316),
    .B1(_06742_),
    .C1(_06744_),
    .D1(_06746_),
    .Y(_06748_));
 sky130_fd_sc_hd__o2bb2ai_4 _17203_ (.A1_N(_06741_),
    .A2_N(_06742_),
    .B1(_06743_),
    .B2(_06745_),
    .Y(_06750_));
 sky130_fd_sc_hd__a21boi_4 _17204_ (.A1(_06748_),
    .A2(_06750_),
    .B1_N(_06740_),
    .Y(_06751_));
 sky130_fd_sc_hd__o211a_2 _17205_ (.A1(_06737_),
    .A2(_06739_),
    .B1(_06748_),
    .C1(_06750_),
    .X(_06752_));
 sky130_fd_sc_hd__nor2_1 _17206_ (.A(_06751_),
    .B(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__a22oi_4 _17207_ (.A1(_04179_),
    .A2(_06447_),
    .B1(_06457_),
    .B2(_06446_),
    .Y(_06754_));
 sky130_fd_sc_hd__a32o_2 _17208_ (.A1(_06219_),
    .A2(_06221_),
    .A3(_04342_),
    .B1(_04364_),
    .B2(net17),
    .X(_06755_));
 sky130_fd_sc_hd__a41oi_4 _17209_ (.A1(_11420_),
    .A2(net284),
    .A3(_05926_),
    .A4(_06450_),
    .B1(_04201_),
    .Y(_06756_));
 sky130_fd_sc_hd__o41ai_4 _17210_ (.A1(net17),
    .A2(net18),
    .A3(net245),
    .A4(net241),
    .B1(net19),
    .Y(_06757_));
 sky130_fd_sc_hd__nor3_2 _17211_ (.A(net17),
    .B(net18),
    .C(net19),
    .Y(_06758_));
 sky130_fd_sc_hd__or3_4 _17212_ (.A(net17),
    .B(net18),
    .C(net19),
    .X(_06759_));
 sky130_fd_sc_hd__nor4_4 _17213_ (.A(net262),
    .B(net244),
    .C(_05927_),
    .D(_06759_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand4_4 _17214_ (.A(_06519_),
    .B(_03955_),
    .C(_05926_),
    .D(_06758_),
    .Y(_06762_));
 sky130_fd_sc_hd__o31a_2 _17215_ (.A1(net245),
    .A2(net241),
    .A3(_06759_),
    .B1(_06757_),
    .X(_06763_));
 sky130_fd_sc_hd__o21ai_4 _17216_ (.A1(_05931_),
    .A2(_06759_),
    .B1(_06757_),
    .Y(_06764_));
 sky130_fd_sc_hd__nand3_1 _17217_ (.A(net196),
    .B(net171),
    .C(net33),
    .Y(_06765_));
 sky130_fd_sc_hd__o211ai_2 _17218_ (.A1(net175),
    .A2(_06451_),
    .B1(_04484_),
    .C1(net200),
    .Y(_06766_));
 sky130_fd_sc_hd__nor2_1 _17219_ (.A(_04179_),
    .B(_04331_),
    .Y(_06767_));
 sky130_fd_sc_hd__or3_2 _17220_ (.A(net44),
    .B(_04179_),
    .C(_03286_),
    .X(_06768_));
 sky130_fd_sc_hd__or4_1 _17221_ (.A(net44),
    .B(net19),
    .C(_04179_),
    .D(_03286_),
    .X(_06769_));
 sky130_fd_sc_hd__nand3_4 _17222_ (.A(_06765_),
    .B(_06766_),
    .C(_06768_),
    .Y(_06770_));
 sky130_fd_sc_hd__a21oi_4 _17223_ (.A1(_06769_),
    .A2(_06770_),
    .B1(_06755_),
    .Y(_06772_));
 sky130_fd_sc_hd__o41a_1 _17224_ (.A1(_03286_),
    .A2(net44),
    .A3(_04179_),
    .A4(net19),
    .B1(_06755_),
    .X(_06773_));
 sky130_fd_sc_hd__o311a_2 _17225_ (.A1(_03286_),
    .A2(_06764_),
    .A3(_06768_),
    .B1(_06770_),
    .C1(_06755_),
    .X(_06774_));
 sky130_fd_sc_hd__a211oi_2 _17226_ (.A1(_06773_),
    .A2(_06770_),
    .B1(_06754_),
    .C1(_06772_),
    .Y(_06775_));
 sky130_fd_sc_hd__a211o_1 _17227_ (.A1(_06773_),
    .A2(_06770_),
    .B1(_06754_),
    .C1(_06772_),
    .X(_06776_));
 sky130_fd_sc_hd__o21a_2 _17228_ (.A1(_06772_),
    .A2(_06774_),
    .B1(_06754_),
    .X(_06777_));
 sky130_fd_sc_hd__o21ai_4 _17229_ (.A1(_06772_),
    .A2(_06774_),
    .B1(_06754_),
    .Y(_06778_));
 sky130_fd_sc_hd__and3_1 _17230_ (.A(_06753_),
    .B(_06776_),
    .C(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__nand3_1 _17231_ (.A(_06753_),
    .B(_06776_),
    .C(_06778_),
    .Y(_06780_));
 sky130_fd_sc_hd__o22ai_4 _17232_ (.A1(_06751_),
    .A2(_06752_),
    .B1(_06775_),
    .B2(_06777_),
    .Y(_06781_));
 sky130_fd_sc_hd__o211ai_2 _17233_ (.A1(_06751_),
    .A2(_06752_),
    .B1(_06776_),
    .C1(_06778_),
    .Y(_06783_));
 sky130_fd_sc_hd__o21ai_1 _17234_ (.A1(_06775_),
    .A2(_06777_),
    .B1(_06753_),
    .Y(_06784_));
 sky130_fd_sc_hd__nand2_1 _17235_ (.A(_06736_),
    .B(_06781_),
    .Y(_06785_));
 sky130_fd_sc_hd__nand3_4 _17236_ (.A(_06736_),
    .B(_06780_),
    .C(_06781_),
    .Y(_06786_));
 sky130_fd_sc_hd__nand3_4 _17237_ (.A(_06784_),
    .B(_06735_),
    .C(_06783_),
    .Y(_06787_));
 sky130_fd_sc_hd__a21o_1 _17238_ (.A1(_06786_),
    .A2(_06787_),
    .B1(_06734_),
    .X(_06788_));
 sky130_fd_sc_hd__o211ai_2 _17239_ (.A1(_06779_),
    .A2(_06785_),
    .B1(_06787_),
    .C1(_06734_),
    .Y(_06789_));
 sky130_fd_sc_hd__nand4_4 _17240_ (.A(_06730_),
    .B(_06732_),
    .C(_06786_),
    .D(_06787_),
    .Y(_06790_));
 sky130_fd_sc_hd__a22o_2 _17241_ (.A1(_06730_),
    .A2(_06732_),
    .B1(_06786_),
    .B2(_06787_),
    .X(_06791_));
 sky130_fd_sc_hd__nand3_4 _17242_ (.A(_06791_),
    .B(_06704_),
    .C(_06790_),
    .Y(_06792_));
 sky130_fd_sc_hd__a21oi_2 _17243_ (.A1(_06790_),
    .A2(_06791_),
    .B1(_06704_),
    .Y(_06794_));
 sky130_fd_sc_hd__nand3_4 _17244_ (.A(_06706_),
    .B(_06788_),
    .C(_06789_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand3_2 _17245_ (.A(net223),
    .B(net291),
    .C(net188),
    .Y(_06796_));
 sky130_fd_sc_hd__or3b_1 _17246_ (.A(net64),
    .B(_04069_),
    .C_N(net63),
    .X(_06797_));
 sky130_fd_sc_hd__and3_1 _17247_ (.A(_03971_),
    .B(net8),
    .C(net64),
    .X(_06798_));
 sky130_fd_sc_hd__a31oi_4 _17248_ (.A1(_04132_),
    .A2(net289),
    .A3(net230),
    .B1(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__a21oi_4 _17249_ (.A1(_06796_),
    .A2(_06797_),
    .B1(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__o211a_1 _17250_ (.A1(_04069_),
    .A2(_08283_),
    .B1(_06796_),
    .C1(_06799_),
    .X(_06801_));
 sky130_fd_sc_hd__o211ai_2 _17251_ (.A1(_04069_),
    .A2(_08283_),
    .B1(_06796_),
    .C1(_06799_),
    .Y(_06802_));
 sky130_fd_sc_hd__a32o_1 _17252_ (.A1(_03952_),
    .A2(net232),
    .A3(net252),
    .B1(_11793_),
    .B2(net7),
    .X(_06803_));
 sky130_fd_sc_hd__o21bai_4 _17253_ (.A1(_06800_),
    .A2(_06801_),
    .B1_N(_06803_),
    .Y(_06805_));
 sky130_fd_sc_hd__and2_1 _17254_ (.A(_06802_),
    .B(_06803_),
    .X(_06806_));
 sky130_fd_sc_hd__nand2_1 _17255_ (.A(_06802_),
    .B(_06803_),
    .Y(_06807_));
 sky130_fd_sc_hd__nand3b_1 _17256_ (.A_N(_06800_),
    .B(_06802_),
    .C(_06803_),
    .Y(_06808_));
 sky130_fd_sc_hd__a21o_1 _17257_ (.A1(_06545_),
    .A2(_06553_),
    .B1(_06554_),
    .X(_06809_));
 sky130_fd_sc_hd__o211a_1 _17258_ (.A1(_06800_),
    .A2(_06807_),
    .B1(_06809_),
    .C1(_06805_),
    .X(_06810_));
 sky130_fd_sc_hd__o221ai_4 _17259_ (.A1(_06800_),
    .A2(_06807_),
    .B1(_06554_),
    .B2(_06556_),
    .C1(_06805_),
    .Y(_06811_));
 sky130_fd_sc_hd__a21oi_2 _17260_ (.A1(_06805_),
    .A2(_06808_),
    .B1(_06809_),
    .Y(_06812_));
 sky130_fd_sc_hd__a21o_1 _17261_ (.A1(_06805_),
    .A2(_06808_),
    .B1(_06809_),
    .X(_06813_));
 sky130_fd_sc_hd__o22a_1 _17262_ (.A1(_13021_),
    .A2(_02869_),
    .B1(_02891_),
    .B2(_04004_),
    .X(_06814_));
 sky130_fd_sc_hd__a32o_1 _17263_ (.A1(net235),
    .A2(net251),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net4),
    .X(_06816_));
 sky130_fd_sc_hd__a32oi_4 _17264_ (.A1(_00625_),
    .A2(net250),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net5),
    .Y(_06817_));
 sky130_fd_sc_hd__or3_1 _17265_ (.A(net36),
    .B(_04026_),
    .C(_03993_),
    .X(_06818_));
 sky130_fd_sc_hd__a311o_2 _17266_ (.A1(_06519_),
    .A2(net286),
    .A3(_02432_),
    .B1(_12341_),
    .C1(_02410_),
    .X(_06819_));
 sky130_fd_sc_hd__o211ai_1 _17267_ (.A1(_04026_),
    .A2(_12363_),
    .B1(_06819_),
    .C1(_06817_),
    .Y(_06820_));
 sky130_fd_sc_hd__a21oi_1 _17268_ (.A1(_06818_),
    .A2(_06819_),
    .B1(_06817_),
    .Y(_06821_));
 sky130_fd_sc_hd__a21o_1 _17269_ (.A1(_06818_),
    .A2(_06819_),
    .B1(_06817_),
    .X(_06822_));
 sky130_fd_sc_hd__a31oi_1 _17270_ (.A1(_06817_),
    .A2(_06818_),
    .A3(_06819_),
    .B1(_06814_),
    .Y(_06823_));
 sky130_fd_sc_hd__a21oi_1 _17271_ (.A1(_06816_),
    .A2(_06820_),
    .B1(_06821_),
    .Y(_06824_));
 sky130_fd_sc_hd__o21ai_1 _17272_ (.A1(_06816_),
    .A2(_06820_),
    .B1(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__o21a_1 _17273_ (.A1(_06814_),
    .A2(_06822_),
    .B1(_06825_),
    .X(_06827_));
 sky130_fd_sc_hd__o21ai_2 _17274_ (.A1(_06814_),
    .A2(_06822_),
    .B1(_06825_),
    .Y(_06828_));
 sky130_fd_sc_hd__o21ai_4 _17275_ (.A1(_06810_),
    .A2(_06812_),
    .B1(_06827_),
    .Y(_06829_));
 sky130_fd_sc_hd__nand3_2 _17276_ (.A(_06811_),
    .B(_06813_),
    .C(_06828_),
    .Y(_06830_));
 sky130_fd_sc_hd__a32oi_4 _17277_ (.A1(_06509_),
    .A2(_06510_),
    .A3(_06511_),
    .B1(_06514_),
    .B2(_06199_),
    .Y(_06831_));
 sky130_fd_sc_hd__a21oi_4 _17278_ (.A1(_06829_),
    .A2(_06830_),
    .B1(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__a221o_1 _17279_ (.A1(_06198_),
    .A2(_06512_),
    .B1(_06829_),
    .B2(_06830_),
    .C1(_06513_),
    .X(_06833_));
 sky130_fd_sc_hd__and3_2 _17280_ (.A(_06829_),
    .B(_06831_),
    .C(_06830_),
    .X(_06834_));
 sky130_fd_sc_hd__nand3_2 _17281_ (.A(_06829_),
    .B(_06831_),
    .C(_06830_),
    .Y(_06835_));
 sky130_fd_sc_hd__o31a_2 _17282_ (.A1(_06542_),
    .A2(_06556_),
    .A3(_06558_),
    .B1(_06567_),
    .X(_06836_));
 sky130_fd_sc_hd__a21o_2 _17283_ (.A1(_06561_),
    .A2(_06567_),
    .B1(_06832_),
    .X(_06838_));
 sky130_fd_sc_hd__nor2_1 _17284_ (.A(_06834_),
    .B(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__a211o_1 _17285_ (.A1(_06561_),
    .A2(_06567_),
    .B1(_06832_),
    .C1(_06834_),
    .X(_06840_));
 sky130_fd_sc_hd__o21ai_4 _17286_ (.A1(_06832_),
    .A2(_06834_),
    .B1(_06836_),
    .Y(_06841_));
 sky130_fd_sc_hd__inv_2 _17287_ (.A(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__o2bb2a_1 _17288_ (.A1_N(_06561_),
    .A2_N(_06567_),
    .B1(_06832_),
    .B2(_06834_),
    .X(_06843_));
 sky130_fd_sc_hd__and3_1 _17289_ (.A(_06833_),
    .B(_06835_),
    .C(_06836_),
    .X(_06844_));
 sky130_fd_sc_hd__o21ai_1 _17290_ (.A1(_06834_),
    .A2(_06838_),
    .B1(_06841_),
    .Y(_06845_));
 sky130_fd_sc_hd__o2111ai_4 _17291_ (.A1(_06834_),
    .A2(_06838_),
    .B1(_06841_),
    .C1(_06795_),
    .D1(_06792_),
    .Y(_06846_));
 sky130_fd_sc_hd__o2bb2ai_2 _17292_ (.A1_N(_06792_),
    .A2_N(_06795_),
    .B1(_06839_),
    .B2(_06842_),
    .Y(_06847_));
 sky130_fd_sc_hd__nand3_2 _17293_ (.A(_06792_),
    .B(_06795_),
    .C(_06845_),
    .Y(_06849_));
 sky130_fd_sc_hd__o2bb2ai_2 _17294_ (.A1_N(_06792_),
    .A2_N(_06795_),
    .B1(_06843_),
    .B2(_06844_),
    .Y(_06850_));
 sky130_fd_sc_hd__nand3_2 _17295_ (.A(_06847_),
    .B(_06703_),
    .C(_06846_),
    .Y(_06851_));
 sky130_fd_sc_hd__o211a_2 _17296_ (.A1(_06523_),
    .A2(_06702_),
    .B1(_06849_),
    .C1(_06850_),
    .X(_06852_));
 sky130_fd_sc_hd__o211ai_4 _17297_ (.A1(_06523_),
    .A2(_06702_),
    .B1(_06849_),
    .C1(_06850_),
    .Y(_06853_));
 sky130_fd_sc_hd__a21o_1 _17298_ (.A1(_06851_),
    .A2(_06853_),
    .B1(_06701_),
    .X(_06854_));
 sky130_fd_sc_hd__nand3_2 _17299_ (.A(_06701_),
    .B(_06851_),
    .C(_06853_),
    .Y(_06855_));
 sky130_fd_sc_hd__nand4_2 _17300_ (.A(_06698_),
    .B(_06700_),
    .C(_06851_),
    .D(_06853_),
    .Y(_06856_));
 sky130_fd_sc_hd__a22o_1 _17301_ (.A1(_06698_),
    .A2(_06700_),
    .B1(_06851_),
    .B2(_06853_),
    .X(_06857_));
 sky130_fd_sc_hd__o211a_2 _17302_ (.A1(_06589_),
    .A2(_06593_),
    .B1(_06856_),
    .C1(_06857_),
    .X(_06858_));
 sky130_fd_sc_hd__o211ai_4 _17303_ (.A1(_06589_),
    .A2(_06593_),
    .B1(_06856_),
    .C1(_06857_),
    .Y(_06860_));
 sky130_fd_sc_hd__nand3_2 _17304_ (.A(_06854_),
    .B(_06855_),
    .C(_06626_),
    .Y(_06861_));
 sky130_fd_sc_hd__nand2_1 _17305_ (.A(_06342_),
    .B(_06345_),
    .Y(_06862_));
 sky130_fd_sc_hd__and2_4 _17306_ (.A(_04190_),
    .B(net51),
    .X(_06863_));
 sky130_fd_sc_hd__nand2_8 _17307_ (.A(_04190_),
    .B(net51),
    .Y(_06864_));
 sky130_fd_sc_hd__nor2_8 _17308_ (.A(net51),
    .B(_04190_),
    .Y(_06865_));
 sky130_fd_sc_hd__or2_4 _17309_ (.A(net51),
    .B(_04190_),
    .X(_06866_));
 sky130_fd_sc_hd__o21a_1 _17310_ (.A1(_06863_),
    .A2(_06865_),
    .B1(net1),
    .X(_06867_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(net23),
    .B(_06029_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand3_2 _17312_ (.A(net318),
    .B(_04452_),
    .C(_06026_),
    .Y(_06869_));
 sky130_fd_sc_hd__a21oi_1 _17313_ (.A1(_04309_),
    .A2(_04517_),
    .B1(_06325_),
    .Y(_06871_));
 sky130_fd_sc_hd__o21ai_4 _17314_ (.A1(_04298_),
    .A2(_04506_),
    .B1(_06324_),
    .Y(_06872_));
 sky130_fd_sc_hd__and3_1 _17315_ (.A(_04190_),
    .B(net49),
    .C(net12),
    .X(_06873_));
 sky130_fd_sc_hd__nand2_1 _17316_ (.A(net12),
    .B(_06326_),
    .Y(_06874_));
 sky130_fd_sc_hd__o2bb2a_1 _17317_ (.A1_N(_06868_),
    .A2_N(_06869_),
    .B1(_06871_),
    .B2(_06873_),
    .X(_06875_));
 sky130_fd_sc_hd__o2bb2ai_2 _17318_ (.A1_N(_06868_),
    .A2_N(_06869_),
    .B1(_06871_),
    .B2(_06873_),
    .Y(_06876_));
 sky130_fd_sc_hd__nand4_4 _17319_ (.A(_06868_),
    .B(_06869_),
    .C(_06872_),
    .D(_06874_),
    .Y(_06877_));
 sky130_fd_sc_hd__o2111ai_4 _17320_ (.A1(_06863_),
    .A2(_06865_),
    .B1(_06877_),
    .C1(net1),
    .D1(_06876_),
    .Y(_06878_));
 sky130_fd_sc_hd__a21o_1 _17321_ (.A1(_06876_),
    .A2(_06877_),
    .B1(_06867_),
    .X(_06879_));
 sky130_fd_sc_hd__nor2_1 _17322_ (.A(_06381_),
    .B(_06390_),
    .Y(_06880_));
 sky130_fd_sc_hd__o221ai_4 _17323_ (.A1(_04474_),
    .A2(_05763_),
    .B1(_05766_),
    .B2(_03396_),
    .C1(_06391_),
    .Y(_06882_));
 sky130_fd_sc_hd__o2111ai_4 _17324_ (.A1(_06384_),
    .A2(_06386_),
    .B1(_06878_),
    .C1(_06879_),
    .D1(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__o2bb2ai_2 _17325_ (.A1_N(_06878_),
    .A2_N(_06879_),
    .B1(_06880_),
    .B2(_06388_),
    .Y(_06884_));
 sky130_fd_sc_hd__a22oi_1 _17326_ (.A1(_06333_),
    .A2(_06327_),
    .B1(_06884_),
    .B2(_06883_),
    .Y(_06885_));
 sky130_fd_sc_hd__o2111a_1 _17327_ (.A1(_06329_),
    .A2(_06330_),
    .B1(_06327_),
    .C1(_06883_),
    .D1(_06884_),
    .X(_06886_));
 sky130_fd_sc_hd__o211a_1 _17328_ (.A1(_06328_),
    .A2(_06331_),
    .B1(_06883_),
    .C1(_06884_),
    .X(_06887_));
 sky130_fd_sc_hd__a21oi_1 _17329_ (.A1(_06883_),
    .A2(_06884_),
    .B1(_06335_),
    .Y(_06888_));
 sky130_fd_sc_hd__a2bb2oi_1 _17330_ (.A1_N(_06374_),
    .A2_N(_06379_),
    .B1(_06394_),
    .B2(_06378_),
    .Y(_06889_));
 sky130_fd_sc_hd__o2bb2ai_1 _17331_ (.A1_N(_06394_),
    .A2_N(_06378_),
    .B1(_06374_),
    .B2(_06379_),
    .Y(_06890_));
 sky130_fd_sc_hd__o21a_1 _17332_ (.A1(_06885_),
    .A2(_06886_),
    .B1(_06889_),
    .X(_06891_));
 sky130_fd_sc_hd__o21ai_1 _17333_ (.A1(_06885_),
    .A2(_06886_),
    .B1(_06889_),
    .Y(_06893_));
 sky130_fd_sc_hd__o21ai_2 _17334_ (.A1(_06887_),
    .A2(_06888_),
    .B1(_06890_),
    .Y(_06894_));
 sky130_fd_sc_hd__o2bb2ai_1 _17335_ (.A1_N(_06893_),
    .A2_N(_06894_),
    .B1(_06337_),
    .B2(_06338_),
    .Y(_06895_));
 sky130_fd_sc_hd__nand2_1 _17336_ (.A(_06894_),
    .B(_06339_),
    .Y(_06896_));
 sky130_fd_sc_hd__o21ai_2 _17337_ (.A1(_06891_),
    .A2(_06896_),
    .B1(_06895_),
    .Y(_06897_));
 sky130_fd_sc_hd__o211a_1 _17338_ (.A1(_06891_),
    .A2(_06896_),
    .B1(_06895_),
    .C1(_06862_),
    .X(_06898_));
 sky130_fd_sc_hd__xnor2_1 _17339_ (.A(_06862_),
    .B(_06897_),
    .Y(_06899_));
 sky130_fd_sc_hd__xor2_1 _17340_ (.A(_06862_),
    .B(_06897_),
    .X(_06900_));
 sky130_fd_sc_hd__nand2_1 _17341_ (.A(_06436_),
    .B(_06438_),
    .Y(_06901_));
 sky130_fd_sc_hd__and3_1 _17342_ (.A(_06436_),
    .B(_06443_),
    .C(_06900_),
    .X(_06902_));
 sky130_fd_sc_hd__o211ai_1 _17343_ (.A1(_06438_),
    .A2(_06434_),
    .B1(_06436_),
    .C1(_06900_),
    .Y(_06904_));
 sky130_fd_sc_hd__o221a_1 _17344_ (.A1(_06433_),
    .A2(_06178_),
    .B1(_06437_),
    .B2(_06435_),
    .C1(_06899_),
    .X(_06905_));
 sky130_fd_sc_hd__o211ai_2 _17345_ (.A1(_06178_),
    .A2(_06433_),
    .B1(_06899_),
    .C1(_06901_),
    .Y(_06906_));
 sky130_fd_sc_hd__nand2_1 _17346_ (.A(_06904_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__o31a_1 _17347_ (.A1(_06035_),
    .A2(_06036_),
    .A3(_06344_),
    .B1(_06907_),
    .X(_06908_));
 sky130_fd_sc_hd__and3_1 _17348_ (.A(_06904_),
    .B(_06906_),
    .C(_06347_),
    .X(_06909_));
 sky130_fd_sc_hd__nor2_1 _17349_ (.A(_06908_),
    .B(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__xor2_1 _17350_ (.A(_06347_),
    .B(_06907_),
    .X(_06911_));
 sky130_fd_sc_hd__a21oi_1 _17351_ (.A1(_06860_),
    .A2(_06861_),
    .B1(_06910_),
    .Y(_06912_));
 sky130_fd_sc_hd__o2bb2ai_2 _17352_ (.A1_N(_06860_),
    .A2_N(_06861_),
    .B1(_06908_),
    .B2(_06909_),
    .Y(_06913_));
 sky130_fd_sc_hd__a31oi_4 _17353_ (.A1(_06626_),
    .A2(_06854_),
    .A3(_06855_),
    .B1(_06911_),
    .Y(_06915_));
 sky130_fd_sc_hd__nand2_1 _17354_ (.A(_06861_),
    .B(_06910_),
    .Y(_06916_));
 sky130_fd_sc_hd__nand3_1 _17355_ (.A(_06860_),
    .B(_06861_),
    .C(_06910_),
    .Y(_06917_));
 sky130_fd_sc_hd__o21ai_1 _17356_ (.A1(_06858_),
    .A2(_06916_),
    .B1(_06913_),
    .Y(_06918_));
 sky130_fd_sc_hd__a22oi_2 _17357_ (.A1(_06598_),
    .A2(_06624_),
    .B1(_06913_),
    .B2(_06917_),
    .Y(_06919_));
 sky130_fd_sc_hd__a221oi_4 _17358_ (.A1(_06915_),
    .A2(_06860_),
    .B1(_06601_),
    .B2(_06597_),
    .C1(_06912_),
    .Y(_06920_));
 sky130_fd_sc_hd__o2111ai_4 _17359_ (.A1(_06916_),
    .A2(_06858_),
    .B1(_06624_),
    .C1(_06598_),
    .D1(_06913_),
    .Y(_06921_));
 sky130_fd_sc_hd__o2bb2ai_2 _17360_ (.A1_N(_06625_),
    .A2_N(_06918_),
    .B1(_06350_),
    .B2(_06356_),
    .Y(_06922_));
 sky130_fd_sc_hd__o21ai_1 _17361_ (.A1(_06919_),
    .A2(_06920_),
    .B1(_06623_),
    .Y(_06923_));
 sky130_fd_sc_hd__o22ai_2 _17362_ (.A1(_06350_),
    .A2(_06356_),
    .B1(_06919_),
    .B2(_06920_),
    .Y(_06924_));
 sky130_fd_sc_hd__nand3b_1 _17363_ (.A_N(_06919_),
    .B(_06921_),
    .C(_06623_),
    .Y(_06926_));
 sky130_fd_sc_hd__o2bb2ai_1 _17364_ (.A1_N(_06043_),
    .A2_N(_06608_),
    .B1(_06602_),
    .B2(_06605_),
    .Y(_06927_));
 sky130_fd_sc_hd__o2bb2a_1 _17365_ (.A1_N(_06043_),
    .A2_N(_06608_),
    .B1(_06605_),
    .B2(_06602_),
    .X(_06928_));
 sky130_fd_sc_hd__nand3_1 _17366_ (.A(_06924_),
    .B(_06926_),
    .C(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__o211ai_4 _17367_ (.A1(_06920_),
    .A2(_06922_),
    .B1(_06927_),
    .C1(_06923_),
    .Y(_06930_));
 sky130_fd_sc_hd__a21oi_1 _17368_ (.A1(_06929_),
    .A2(_06930_),
    .B1(_06615_),
    .Y(_06931_));
 sky130_fd_sc_hd__a31oi_2 _17369_ (.A1(_06924_),
    .A2(_06926_),
    .A3(_06928_),
    .B1(_06616_),
    .Y(_06932_));
 sky130_fd_sc_hd__nand3_1 _17370_ (.A(_06615_),
    .B(_06929_),
    .C(_06930_),
    .Y(_06933_));
 sky130_fd_sc_hd__a21oi_2 _17371_ (.A1(_06930_),
    .A2(_06932_),
    .B1(_06931_),
    .Y(_06934_));
 sky130_fd_sc_hd__o22ai_2 _17372_ (.A1(_06613_),
    .A2(_06620_),
    .B1(_06309_),
    .B2(_06617_),
    .Y(_06935_));
 sky130_fd_sc_hd__a31o_1 _17373_ (.A1(_06320_),
    .A2(_06621_),
    .A3(_06310_),
    .B1(_06935_),
    .X(_06937_));
 sky130_fd_sc_hd__xor2_1 _17374_ (.A(_06934_),
    .B(_06937_),
    .X(net83));
 sky130_fd_sc_hd__o21ai_1 _17375_ (.A1(_06623_),
    .A2(_06919_),
    .B1(_06921_),
    .Y(_06938_));
 sky130_fd_sc_hd__a32o_1 _17376_ (.A1(_06597_),
    .A2(_06918_),
    .A3(_06601_),
    .B1(_06921_),
    .B2(_06623_),
    .X(_06939_));
 sky130_fd_sc_hd__o31a_1 _17377_ (.A1(_06035_),
    .A2(_06036_),
    .A3(_06344_),
    .B1(_06906_),
    .X(_06940_));
 sky130_fd_sc_hd__and3_1 _17378_ (.A(_06904_),
    .B(_06037_),
    .C(_06346_),
    .X(_06941_));
 sky130_fd_sc_hd__a31o_1 _17379_ (.A1(_06436_),
    .A2(_06443_),
    .A3(_06900_),
    .B1(_06940_),
    .X(_06942_));
 sky130_fd_sc_hd__nand2_1 _17380_ (.A(_06860_),
    .B(_06916_),
    .Y(_06943_));
 sky130_fd_sc_hd__a32oi_4 _17381_ (.A1(_06703_),
    .A2(_06846_),
    .A3(_06847_),
    .B1(_06700_),
    .B2(_06698_),
    .Y(_06944_));
 sky130_fd_sc_hd__o21ai_1 _17382_ (.A1(_06701_),
    .A2(_06852_),
    .B1(_06851_),
    .Y(_06945_));
 sky130_fd_sc_hd__o21ai_2 _17383_ (.A1(_06836_),
    .A2(_06832_),
    .B1(_06835_),
    .Y(_06947_));
 sky130_fd_sc_hd__nand2_1 _17384_ (.A(_06679_),
    .B(_06684_),
    .Y(_06948_));
 sky130_fd_sc_hd__o22a_1 _17385_ (.A1(_09720_),
    .A2(_04268_),
    .B1(_04270_),
    .B2(_03960_),
    .X(_06949_));
 sky130_fd_sc_hd__a32o_1 _17386_ (.A1(net255),
    .A2(_09698_),
    .A3(net280),
    .B1(_04269_),
    .B2(net2),
    .X(_06950_));
 sky130_fd_sc_hd__o2111ai_4 _17387_ (.A1(_11387_),
    .A2(_12988_),
    .B1(net39),
    .C1(net235),
    .D1(_04037_),
    .Y(_06951_));
 sky130_fd_sc_hd__or3_1 _17388_ (.A(net39),
    .B(_04037_),
    .C(_04004_),
    .X(_06952_));
 sky130_fd_sc_hd__nor2_2 _17389_ (.A(_03982_),
    .B(_04218_),
    .Y(_06953_));
 sky130_fd_sc_hd__o311a_1 _17390_ (.A1(_04747_),
    .A2(net264),
    .A3(_11387_),
    .B1(net281),
    .C1(_11354_),
    .X(_06954_));
 sky130_fd_sc_hd__a21oi_1 _17391_ (.A1(_11442_),
    .A2(net281),
    .B1(_06953_),
    .Y(_06955_));
 sky130_fd_sc_hd__o221ai_4 _17392_ (.A1(_04004_),
    .A2(_03737_),
    .B1(_04216_),
    .B2(net236),
    .C1(_06951_),
    .Y(_06956_));
 sky130_fd_sc_hd__o211ai_1 _17393_ (.A1(_04004_),
    .A2(_03737_),
    .B1(_06951_),
    .C1(_06955_),
    .Y(_06958_));
 sky130_fd_sc_hd__o2bb2ai_4 _17394_ (.A1_N(_06951_),
    .A2_N(_06952_),
    .B1(_06953_),
    .B2(_06954_),
    .Y(_06959_));
 sky130_fd_sc_hd__o21ai_1 _17395_ (.A1(_06953_),
    .A2(_06956_),
    .B1(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__o211a_1 _17396_ (.A1(_06953_),
    .A2(_06956_),
    .B1(_06959_),
    .C1(_06950_),
    .X(_06961_));
 sky130_fd_sc_hd__o211ai_2 _17397_ (.A1(_06953_),
    .A2(_06956_),
    .B1(_06959_),
    .C1(_06950_),
    .Y(_06962_));
 sky130_fd_sc_hd__a21oi_1 _17398_ (.A1(_06958_),
    .A2(_06959_),
    .B1(_06950_),
    .Y(_06963_));
 sky130_fd_sc_hd__a21o_1 _17399_ (.A1(_06958_),
    .A2(_06959_),
    .B1(_06950_),
    .X(_06964_));
 sky130_fd_sc_hd__o211ai_2 _17400_ (.A1(_06821_),
    .A2(_06823_),
    .B1(_06962_),
    .C1(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__o21ai_2 _17401_ (.A1(_06961_),
    .A2(_06963_),
    .B1(_06824_),
    .Y(_06966_));
 sky130_fd_sc_hd__o21ai_2 _17402_ (.A1(_06664_),
    .A2(_06671_),
    .B1(_06670_),
    .Y(_06967_));
 sky130_fd_sc_hd__a21oi_1 _17403_ (.A1(_06965_),
    .A2(_06966_),
    .B1(_06967_),
    .Y(_06969_));
 sky130_fd_sc_hd__a21o_1 _17404_ (.A1(_06965_),
    .A2(_06966_),
    .B1(_06967_),
    .X(_06970_));
 sky130_fd_sc_hd__and3_1 _17405_ (.A(_06965_),
    .B(_06966_),
    .C(_06967_),
    .X(_06971_));
 sky130_fd_sc_hd__nand3_1 _17406_ (.A(_06965_),
    .B(_06966_),
    .C(_06967_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand3_2 _17407_ (.A(_06948_),
    .B(_06970_),
    .C(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__a21oi_2 _17408_ (.A1(_06970_),
    .A2(_06972_),
    .B1(_06948_),
    .Y(_06974_));
 sky130_fd_sc_hd__o21bai_1 _17409_ (.A1(_06969_),
    .A2(_06971_),
    .B1_N(_06948_),
    .Y(_06975_));
 sky130_fd_sc_hd__nand2_1 _17410_ (.A(_06973_),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__a32oi_4 _17411_ (.A1(net266),
    .A2(net302),
    .A3(net275),
    .B1(_05765_),
    .B2(net27),
    .Y(_06977_));
 sky130_fd_sc_hd__a31oi_4 _17412_ (.A1(_04397_),
    .A2(_04725_),
    .A3(_05425_),
    .B1(_05463_),
    .Y(_06978_));
 sky130_fd_sc_hd__a22oi_4 _17413_ (.A1(net28),
    .A2(_05464_),
    .B1(_05414_),
    .B2(_06978_),
    .Y(_06980_));
 sky130_fd_sc_hd__or3_1 _17414_ (.A(net46),
    .B(_04124_),
    .C(_03835_),
    .X(_06981_));
 sky130_fd_sc_hd__nand4_1 _17415_ (.A(_04124_),
    .B(_05841_),
    .C(net265),
    .D(net46),
    .Y(_06982_));
 sky130_fd_sc_hd__a32oi_2 _17416_ (.A1(_05841_),
    .A2(net265),
    .A3(net276),
    .B1(_05228_),
    .B2(net29),
    .Y(_06983_));
 sky130_fd_sc_hd__a21oi_2 _17417_ (.A1(_06981_),
    .A2(_06982_),
    .B1(_06980_),
    .Y(_06984_));
 sky130_fd_sc_hd__o311a_1 _17418_ (.A1(_03835_),
    .A2(_04124_),
    .A3(net46),
    .B1(_06982_),
    .C1(_06980_),
    .X(_06985_));
 sky130_fd_sc_hd__o21ai_1 _17419_ (.A1(_06984_),
    .A2(_06985_),
    .B1(_06977_),
    .Y(_06986_));
 sky130_fd_sc_hd__or3_1 _17420_ (.A(_06977_),
    .B(_06984_),
    .C(_06985_),
    .X(_06987_));
 sky130_fd_sc_hd__nand2_1 _17421_ (.A(_06986_),
    .B(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__a21o_1 _17422_ (.A1(_06636_),
    .A2(_06637_),
    .B1(_06634_),
    .X(_06989_));
 sky130_fd_sc_hd__a32o_1 _17423_ (.A1(_06486_),
    .A2(net260),
    .A3(_04985_),
    .B1(_04988_),
    .B2(net30),
    .X(_06991_));
 sky130_fd_sc_hd__or3b_1 _17424_ (.A(_03949_),
    .B(net42),
    .C_N(net41),
    .X(_06992_));
 sky130_fd_sc_hd__o211ai_2 _17425_ (.A1(net260),
    .A2(_08656_),
    .B1(net279),
    .C1(_08700_),
    .Y(_06993_));
 sky130_fd_sc_hd__and3_1 _17426_ (.A(_04102_),
    .B(net42),
    .C(net31),
    .X(_06994_));
 sky130_fd_sc_hd__and3_1 _17427_ (.A(_07242_),
    .B(net257),
    .C(net243),
    .X(_06995_));
 sky130_fd_sc_hd__a31oi_1 _17428_ (.A1(_07242_),
    .A2(net257),
    .A3(net243),
    .B1(_06994_),
    .Y(_06996_));
 sky130_fd_sc_hd__a21oi_1 _17429_ (.A1(_06992_),
    .A2(_06993_),
    .B1(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__o2bb2ai_1 _17430_ (.A1_N(_06992_),
    .A2_N(_06993_),
    .B1(_06994_),
    .B2(_06995_),
    .Y(_06998_));
 sky130_fd_sc_hd__o211ai_2 _17431_ (.A1(_03949_),
    .A2(_04483_),
    .B1(_06993_),
    .C1(_06996_),
    .Y(_06999_));
 sky130_fd_sc_hd__nand3_2 _17432_ (.A(_06991_),
    .B(_06998_),
    .C(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__a21o_1 _17433_ (.A1(_06998_),
    .A2(_06999_),
    .B1(_06991_),
    .X(_07002_));
 sky130_fd_sc_hd__nand3_1 _17434_ (.A(_06989_),
    .B(_07000_),
    .C(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__a21oi_1 _17435_ (.A1(_07000_),
    .A2(_07002_),
    .B1(_06989_),
    .Y(_07004_));
 sky130_fd_sc_hd__a21o_1 _17436_ (.A1(_07000_),
    .A2(_07002_),
    .B1(_06989_),
    .X(_07005_));
 sky130_fd_sc_hd__and3_1 _17437_ (.A(_07005_),
    .B(_06988_),
    .C(_07003_),
    .X(_07006_));
 sky130_fd_sc_hd__a21oi_2 _17438_ (.A1(_07003_),
    .A2(_07005_),
    .B1(_06988_),
    .Y(_07007_));
 sky130_fd_sc_hd__nor2_1 _17439_ (.A(_07006_),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__nand3_1 _17440_ (.A(_06973_),
    .B(_06975_),
    .C(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__a21o_1 _17441_ (.A1(_06973_),
    .A2(_06975_),
    .B1(_07008_),
    .X(_07010_));
 sky130_fd_sc_hd__o21ai_1 _17442_ (.A1(_06974_),
    .A2(_07008_),
    .B1(_06973_),
    .Y(_07011_));
 sky130_fd_sc_hd__o21a_1 _17443_ (.A1(_06974_),
    .A2(_07008_),
    .B1(_06973_),
    .X(_07013_));
 sky130_fd_sc_hd__nand2_1 _17444_ (.A(_06976_),
    .B(_07008_),
    .Y(_07014_));
 sky130_fd_sc_hd__o21ai_1 _17445_ (.A1(_07006_),
    .A2(_07007_),
    .B1(_06973_),
    .Y(_07015_));
 sky130_fd_sc_hd__nand4_2 _17446_ (.A(_06835_),
    .B(_06838_),
    .C(_07009_),
    .D(_07010_),
    .Y(_07016_));
 sky130_fd_sc_hd__o211ai_4 _17447_ (.A1(_06974_),
    .A2(_07015_),
    .B1(_06947_),
    .C1(_07014_),
    .Y(_07017_));
 sky130_fd_sc_hd__inv_2 _17448_ (.A(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__a21o_1 _17449_ (.A1(_06687_),
    .A2(_06660_),
    .B1(_06688_),
    .X(_07019_));
 sky130_fd_sc_hd__a21o_1 _17450_ (.A1(_07016_),
    .A2(_07017_),
    .B1(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__nand2_2 _17451_ (.A(_07016_),
    .B(_07019_),
    .Y(_07021_));
 sky130_fd_sc_hd__nand3_2 _17452_ (.A(_07016_),
    .B(_07017_),
    .C(_07019_),
    .Y(_07022_));
 sky130_fd_sc_hd__o21ai_2 _17453_ (.A1(_07021_),
    .A2(_07018_),
    .B1(_07020_),
    .Y(_07024_));
 sky130_fd_sc_hd__a32oi_4 _17454_ (.A1(_06791_),
    .A2(_06704_),
    .A3(_06790_),
    .B1(_06840_),
    .B2(_06841_),
    .Y(_07025_));
 sky130_fd_sc_hd__a21oi_2 _17455_ (.A1(_06792_),
    .A2(_06845_),
    .B1(_06794_),
    .Y(_07026_));
 sky130_fd_sc_hd__a21oi_1 _17456_ (.A1(_06707_),
    .A2(_06715_),
    .B1(_06712_),
    .Y(_07027_));
 sky130_fd_sc_hd__o21ai_4 _17457_ (.A1(_06740_),
    .A2(_06747_),
    .B1(_06750_),
    .Y(_07028_));
 sky130_fd_sc_hd__and3_1 _17458_ (.A(_03927_),
    .B(net13),
    .C(net61),
    .X(_07029_));
 sky130_fd_sc_hd__a31oi_4 _17459_ (.A1(net212),
    .A2(net183),
    .A3(net292),
    .B1(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__nand3_1 _17460_ (.A(net181),
    .B(net180),
    .C(_05688_),
    .Y(_07031_));
 sky130_fd_sc_hd__or3b_1 _17461_ (.A(net61),
    .B(_04135_),
    .C_N(net60),
    .X(_07032_));
 sky130_fd_sc_hd__a21oi_1 _17462_ (.A1(_07031_),
    .A2(_07032_),
    .B1(_07030_),
    .Y(_07033_));
 sky130_fd_sc_hd__a21o_1 _17463_ (.A1(_07031_),
    .A2(_07032_),
    .B1(_07030_),
    .X(_07035_));
 sky130_fd_sc_hd__and3_2 _17464_ (.A(_07030_),
    .B(_07031_),
    .C(_07032_),
    .X(_07036_));
 sky130_fd_sc_hd__o221ai_4 _17465_ (.A1(_04135_),
    .A2(_05720_),
    .B1(_05294_),
    .B2(_05699_),
    .C1(_07030_),
    .Y(_07037_));
 sky130_fd_sc_hd__a32o_1 _17466_ (.A1(net215),
    .A2(_07658_),
    .A3(net185),
    .B1(_07680_),
    .B2(net11),
    .X(_07038_));
 sky130_fd_sc_hd__o21bai_2 _17467_ (.A1(_07033_),
    .A2(_07036_),
    .B1_N(_07038_),
    .Y(_07039_));
 sky130_fd_sc_hd__nand2_1 _17468_ (.A(_07035_),
    .B(_07038_),
    .Y(_07040_));
 sky130_fd_sc_hd__nand3_1 _17469_ (.A(_07035_),
    .B(_07037_),
    .C(_07038_),
    .Y(_07041_));
 sky130_fd_sc_hd__o21a_1 _17470_ (.A1(_07036_),
    .A2(_07040_),
    .B1(_07039_),
    .X(_07042_));
 sky130_fd_sc_hd__a21oi_1 _17471_ (.A1(_07039_),
    .A2(_07041_),
    .B1(_07028_),
    .Y(_07043_));
 sky130_fd_sc_hd__o211a_2 _17472_ (.A1(_07036_),
    .A2(_07040_),
    .B1(_07039_),
    .C1(_07028_),
    .X(_07044_));
 sky130_fd_sc_hd__o211ai_4 _17473_ (.A1(_07036_),
    .A2(_07040_),
    .B1(_07039_),
    .C1(_07028_),
    .Y(_07046_));
 sky130_fd_sc_hd__o21ai_2 _17474_ (.A1(_07043_),
    .A2(_07044_),
    .B1(_07027_),
    .Y(_07047_));
 sky130_fd_sc_hd__o22ai_4 _17475_ (.A1(_06712_),
    .A2(_06718_),
    .B1(_07028_),
    .B2(_07042_),
    .Y(_07048_));
 sky130_fd_sc_hd__o21ai_4 _17476_ (.A1(_07044_),
    .A2(_07048_),
    .B1(_07047_),
    .Y(_07049_));
 sky130_fd_sc_hd__o32a_1 _17477_ (.A1(_06754_),
    .A2(_06772_),
    .A3(_06774_),
    .B1(_06752_),
    .B2(_06751_),
    .X(_07050_));
 sky130_fd_sc_hd__o21ai_2 _17478_ (.A1(_06751_),
    .A2(_06752_),
    .B1(_06776_),
    .Y(_07051_));
 sky130_fd_sc_hd__o32a_2 _17479_ (.A1(_05238_),
    .A2(_05548_),
    .A3(net206),
    .B1(_05260_),
    .B2(_04146_),
    .X(_07052_));
 sky130_fd_sc_hd__a32o_1 _17480_ (.A1(_05549_),
    .A2(net177),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net15),
    .X(_07053_));
 sky130_fd_sc_hd__o211ai_2 _17481_ (.A1(net232),
    .A2(_05927_),
    .B1(_04889_),
    .C1(_05933_),
    .Y(_07054_));
 sky130_fd_sc_hd__or3b_2 _17482_ (.A(net59),
    .B(_04157_),
    .C_N(net58),
    .X(_07055_));
 sky130_fd_sc_hd__a32oi_4 _17483_ (.A1(_06219_),
    .A2(_06221_),
    .A3(_04627_),
    .B1(_04649_),
    .B2(net17),
    .Y(_07057_));
 sky130_fd_sc_hd__a21oi_4 _17484_ (.A1(_07054_),
    .A2(_07055_),
    .B1(_07057_),
    .Y(_07058_));
 sky130_fd_sc_hd__a21o_1 _17485_ (.A1(_07054_),
    .A2(_07055_),
    .B1(_07057_),
    .X(_07059_));
 sky130_fd_sc_hd__o211a_2 _17486_ (.A1(_04900_),
    .A2(net155),
    .B1(_07055_),
    .C1(_07057_),
    .X(_07060_));
 sky130_fd_sc_hd__o211ai_1 _17487_ (.A1(_04900_),
    .A2(net155),
    .B1(_07055_),
    .C1(_07057_),
    .Y(_07061_));
 sky130_fd_sc_hd__a21oi_1 _17488_ (.A1(_07059_),
    .A2(_07061_),
    .B1(_07053_),
    .Y(_07062_));
 sky130_fd_sc_hd__o21ai_4 _17489_ (.A1(_07058_),
    .A2(_07060_),
    .B1(_07052_),
    .Y(_07063_));
 sky130_fd_sc_hd__nand2_1 _17490_ (.A(_07053_),
    .B(_07059_),
    .Y(_07064_));
 sky130_fd_sc_hd__nor3_2 _17491_ (.A(_07052_),
    .B(_07058_),
    .C(_07060_),
    .Y(_07065_));
 sky130_fd_sc_hd__nand3_1 _17492_ (.A(_07053_),
    .B(_07059_),
    .C(_07061_),
    .Y(_07066_));
 sky130_fd_sc_hd__a32oi_4 _17493_ (.A1(net33),
    .A2(_06763_),
    .A3(_06767_),
    .B1(_06770_),
    .B2(_06755_),
    .Y(_07068_));
 sky130_fd_sc_hd__a32o_1 _17494_ (.A1(net33),
    .A2(_06763_),
    .A3(_06767_),
    .B1(_06770_),
    .B2(_06755_),
    .X(_07069_));
 sky130_fd_sc_hd__nor2_1 _17495_ (.A(_04201_),
    .B(_04331_),
    .Y(_07070_));
 sky130_fd_sc_hd__or3_1 _17496_ (.A(net44),
    .B(_04201_),
    .C(_03286_),
    .X(_07071_));
 sky130_fd_sc_hd__a41o_4 _17497_ (.A1(_06519_),
    .A2(_03955_),
    .A3(_05926_),
    .A4(_06758_),
    .B1(_04212_),
    .X(_07072_));
 sky130_fd_sc_hd__nor4_4 _17498_ (.A(net17),
    .B(net18),
    .C(net19),
    .D(net20),
    .Y(_07073_));
 sky130_fd_sc_hd__or4_4 _17499_ (.A(net17),
    .B(net18),
    .C(net19),
    .D(net20),
    .X(_07074_));
 sky130_fd_sc_hd__nor4_2 _17500_ (.A(net262),
    .B(net244),
    .C(_05927_),
    .D(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__nand4_4 _17501_ (.A(_06519_),
    .B(_03955_),
    .C(_05926_),
    .D(net271),
    .Y(_07076_));
 sky130_fd_sc_hd__a22oi_4 _17502_ (.A1(net205),
    .A2(net271),
    .B1(net171),
    .B2(net20),
    .Y(_07077_));
 sky130_fd_sc_hd__a32o_4 _17503_ (.A1(_03957_),
    .A2(_05926_),
    .A3(net272),
    .B1(net171),
    .B2(net20),
    .X(_07079_));
 sky130_fd_sc_hd__o211ai_2 _17504_ (.A1(net175),
    .A2(_07074_),
    .B1(net33),
    .C1(_07072_),
    .Y(_07080_));
 sky130_fd_sc_hd__and4_1 _17505_ (.A(_07072_),
    .B(_07076_),
    .C(net33),
    .D(_07070_),
    .X(_07081_));
 sky130_fd_sc_hd__nand4_2 _17506_ (.A(_07072_),
    .B(_07076_),
    .C(net33),
    .D(_07070_),
    .Y(_07082_));
 sky130_fd_sc_hd__o311a_2 _17507_ (.A1(_04495_),
    .A2(_06756_),
    .A3(_06761_),
    .B1(_07071_),
    .C1(_07080_),
    .X(_07083_));
 sky130_fd_sc_hd__o311ai_4 _17508_ (.A1(_04495_),
    .A2(_06756_),
    .A3(_06761_),
    .B1(_07071_),
    .C1(_07080_),
    .Y(_07084_));
 sky130_fd_sc_hd__o311a_1 _17509_ (.A1(net245),
    .A2(net241),
    .A3(_06451_),
    .B1(_04342_),
    .C1(net200),
    .X(_07085_));
 sky130_fd_sc_hd__nor2_1 _17510_ (.A(_04179_),
    .B(_04375_),
    .Y(_07086_));
 sky130_fd_sc_hd__a31o_1 _17511_ (.A1(net200),
    .A2(net172),
    .A3(_04342_),
    .B1(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__nand3b_1 _17512_ (.A_N(_07087_),
    .B(_07084_),
    .C(_07082_),
    .Y(_07088_));
 sky130_fd_sc_hd__o2bb2ai_1 _17513_ (.A1_N(_07082_),
    .A2_N(_07084_),
    .B1(_07085_),
    .B2(_07086_),
    .Y(_07090_));
 sky130_fd_sc_hd__o21bai_2 _17514_ (.A1(_07081_),
    .A2(_07083_),
    .B1_N(_07087_),
    .Y(_07091_));
 sky130_fd_sc_hd__o21ai_2 _17515_ (.A1(_07085_),
    .A2(_07086_),
    .B1(_07082_),
    .Y(_07092_));
 sky130_fd_sc_hd__nand3_4 _17516_ (.A(_07090_),
    .B(_07068_),
    .C(_07088_),
    .Y(_07093_));
 sky130_fd_sc_hd__o211a_2 _17517_ (.A1(_07092_),
    .A2(_07083_),
    .B1(_07069_),
    .C1(_07091_),
    .X(_07094_));
 sky130_fd_sc_hd__o211ai_4 _17518_ (.A1(_07092_),
    .A2(_07083_),
    .B1(_07069_),
    .C1(_07091_),
    .Y(_07095_));
 sky130_fd_sc_hd__a2bb2oi_2 _17519_ (.A1_N(_07062_),
    .A2_N(_07065_),
    .B1(_07093_),
    .B2(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__a22o_1 _17520_ (.A1(_07063_),
    .A2(_07066_),
    .B1(_07093_),
    .B2(_07095_),
    .X(_07097_));
 sky130_fd_sc_hd__o211ai_4 _17521_ (.A1(_07064_),
    .A2(_07060_),
    .B1(_07063_),
    .C1(_07093_),
    .Y(_07098_));
 sky130_fd_sc_hd__o2111a_1 _17522_ (.A1(_07064_),
    .A2(_07060_),
    .B1(_07063_),
    .C1(_07093_),
    .D1(_07095_),
    .X(_07099_));
 sky130_fd_sc_hd__o22a_2 _17523_ (.A1(_06777_),
    .A2(_07050_),
    .B1(_07096_),
    .B2(_07099_),
    .X(_07101_));
 sky130_fd_sc_hd__o22ai_4 _17524_ (.A1(_06777_),
    .A2(_07050_),
    .B1(_07096_),
    .B2(_07099_),
    .Y(_07102_));
 sky130_fd_sc_hd__o2111a_2 _17525_ (.A1(_07098_),
    .A2(_07094_),
    .B1(_07051_),
    .C1(_06778_),
    .D1(_07097_),
    .X(_07103_));
 sky130_fd_sc_hd__o2111ai_4 _17526_ (.A1(_07098_),
    .A2(_07094_),
    .B1(_07051_),
    .C1(_06778_),
    .D1(_07097_),
    .Y(_07104_));
 sky130_fd_sc_hd__o21ai_1 _17527_ (.A1(_07101_),
    .A2(_07103_),
    .B1(_07049_),
    .Y(_07105_));
 sky130_fd_sc_hd__o211a_1 _17528_ (.A1(_07048_),
    .A2(_07044_),
    .B1(_07047_),
    .C1(_07102_),
    .X(_07106_));
 sky130_fd_sc_hd__o211ai_2 _17529_ (.A1(_07048_),
    .A2(_07044_),
    .B1(_07047_),
    .C1(_07102_),
    .Y(_07107_));
 sky130_fd_sc_hd__nand3_2 _17530_ (.A(_07049_),
    .B(_07102_),
    .C(_07104_),
    .Y(_07108_));
 sky130_fd_sc_hd__a21o_1 _17531_ (.A1(_07102_),
    .A2(_07104_),
    .B1(_07049_),
    .X(_07109_));
 sky130_fd_sc_hd__a21boi_4 _17532_ (.A1(_06733_),
    .A2(_06787_),
    .B1_N(_06786_),
    .Y(_07110_));
 sky130_fd_sc_hd__o2bb2ai_2 _17533_ (.A1_N(_06733_),
    .A2_N(_06787_),
    .B1(_06785_),
    .B2(_06779_),
    .Y(_07112_));
 sky130_fd_sc_hd__nand3_4 _17534_ (.A(_07108_),
    .B(_07109_),
    .C(_07110_),
    .Y(_07113_));
 sky130_fd_sc_hd__o211ai_4 _17535_ (.A1(_07103_),
    .A2(_07107_),
    .B1(_07112_),
    .C1(_07105_),
    .Y(_07114_));
 sky130_fd_sc_hd__a21boi_2 _17536_ (.A1(_06724_),
    .A2(_06728_),
    .B1_N(_06726_),
    .Y(_07115_));
 sky130_fd_sc_hd__o2bb2ai_2 _17537_ (.A1_N(_06728_),
    .A2_N(_06724_),
    .B1(_06718_),
    .B2(_06725_),
    .Y(_07116_));
 sky130_fd_sc_hd__a21oi_1 _17538_ (.A1(_06802_),
    .A2(_06803_),
    .B1(_06800_),
    .Y(_07117_));
 sky130_fd_sc_hd__o22a_1 _17539_ (.A1(_04059_),
    .A2(_11804_),
    .B1(_04133_),
    .B2(_11782_),
    .X(_07118_));
 sky130_fd_sc_hd__a32o_1 _17540_ (.A1(net228),
    .A2(net252),
    .A3(net230),
    .B1(_11793_),
    .B2(net8),
    .X(_07119_));
 sky130_fd_sc_hd__and3_1 _17541_ (.A(_03971_),
    .B(net9),
    .C(net64),
    .X(_07120_));
 sky130_fd_sc_hd__a31oi_2 _17542_ (.A1(net223),
    .A2(net289),
    .A3(net188),
    .B1(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__a31o_1 _17543_ (.A1(net223),
    .A2(net289),
    .A3(net188),
    .B1(_07120_),
    .X(_07123_));
 sky130_fd_sc_hd__o211ai_2 _17544_ (.A1(net232),
    .A2(_04557_),
    .B1(net291),
    .C1(net219),
    .Y(_07124_));
 sky130_fd_sc_hd__or3b_1 _17545_ (.A(net64),
    .B(_04080_),
    .C_N(net63),
    .X(_07125_));
 sky130_fd_sc_hd__a32o_1 _17546_ (.A1(net219),
    .A2(_04559_),
    .A3(net291),
    .B1(_08272_),
    .B2(net10),
    .X(_07126_));
 sky130_fd_sc_hd__a21oi_2 _17547_ (.A1(_07124_),
    .A2(_07125_),
    .B1(_07121_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21o_1 _17548_ (.A1(_07124_),
    .A2(_07125_),
    .B1(_07121_),
    .X(_07128_));
 sky130_fd_sc_hd__o221a_2 _17549_ (.A1(_04080_),
    .A2(_08283_),
    .B1(_04562_),
    .B2(_08261_),
    .C1(_07121_),
    .X(_07129_));
 sky130_fd_sc_hd__o221ai_1 _17550_ (.A1(_04080_),
    .A2(_08283_),
    .B1(_04562_),
    .B2(_08261_),
    .C1(_07121_),
    .Y(_07130_));
 sky130_fd_sc_hd__o21ai_2 _17551_ (.A1(_07127_),
    .A2(_07129_),
    .B1(_07118_),
    .Y(_07131_));
 sky130_fd_sc_hd__a21o_1 _17552_ (.A1(_07123_),
    .A2(_07126_),
    .B1(_07118_),
    .X(_07132_));
 sky130_fd_sc_hd__nand3_1 _17553_ (.A(_07128_),
    .B(_07130_),
    .C(_07118_),
    .Y(_07134_));
 sky130_fd_sc_hd__o21ai_1 _17554_ (.A1(_07127_),
    .A2(_07129_),
    .B1(_07119_),
    .Y(_07135_));
 sky130_fd_sc_hd__nand3_4 _17555_ (.A(_07135_),
    .B(_07117_),
    .C(_07134_),
    .Y(_07136_));
 sky130_fd_sc_hd__o221a_1 _17556_ (.A1(_06800_),
    .A2(_06806_),
    .B1(_07129_),
    .B2(_07132_),
    .C1(_07131_),
    .X(_07137_));
 sky130_fd_sc_hd__o221ai_4 _17557_ (.A1(_06800_),
    .A2(_06806_),
    .B1(_07129_),
    .B2(_07132_),
    .C1(_07131_),
    .Y(_07138_));
 sky130_fd_sc_hd__a32o_1 _17558_ (.A1(_00625_),
    .A2(net250),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net5),
    .X(_07139_));
 sky130_fd_sc_hd__o211ai_2 _17559_ (.A1(net254),
    .A2(_02442_),
    .B1(_01293_),
    .C1(_02421_),
    .Y(_07140_));
 sky130_fd_sc_hd__or3b_1 _17560_ (.A(net37),
    .B(_04026_),
    .C_N(net36),
    .X(_07141_));
 sky130_fd_sc_hd__nor2_1 _17561_ (.A(_04048_),
    .B(_12363_),
    .Y(_07142_));
 sky130_fd_sc_hd__or3_1 _17562_ (.A(net36),
    .B(_04048_),
    .C(_03993_),
    .X(_07143_));
 sky130_fd_sc_hd__o211ai_2 _17563_ (.A1(net254),
    .A2(_03954_),
    .B1(_12330_),
    .C1(_03952_),
    .Y(_07144_));
 sky130_fd_sc_hd__o211ai_1 _17564_ (.A1(_04026_),
    .A2(_01326_),
    .B1(_07140_),
    .C1(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__o2111ai_2 _17565_ (.A1(_04048_),
    .A2(_12363_),
    .B1(_07140_),
    .C1(_07141_),
    .D1(_07144_),
    .Y(_07146_));
 sky130_fd_sc_hd__a22oi_1 _17566_ (.A1(_07140_),
    .A2(_07141_),
    .B1(_07143_),
    .B2(_07144_),
    .Y(_07147_));
 sky130_fd_sc_hd__a22o_1 _17567_ (.A1(_07140_),
    .A2(_07141_),
    .B1(_07143_),
    .B2(_07144_),
    .X(_07148_));
 sky130_fd_sc_hd__o211a_1 _17568_ (.A1(_07142_),
    .A2(_07145_),
    .B1(_07148_),
    .C1(_07139_),
    .X(_07149_));
 sky130_fd_sc_hd__a21oi_2 _17569_ (.A1(_07146_),
    .A2(_07148_),
    .B1(_07139_),
    .Y(_07150_));
 sky130_fd_sc_hd__nor2_1 _17570_ (.A(_07149_),
    .B(_07150_),
    .Y(_07151_));
 sky130_fd_sc_hd__a21bo_1 _17571_ (.A1(_07136_),
    .A2(_07138_),
    .B1_N(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__o211ai_2 _17572_ (.A1(_07149_),
    .A2(_07150_),
    .B1(_07136_),
    .C1(_07138_),
    .Y(_07153_));
 sky130_fd_sc_hd__o2bb2ai_2 _17573_ (.A1_N(_07136_),
    .A2_N(_07138_),
    .B1(_07149_),
    .B2(_07150_),
    .Y(_07155_));
 sky130_fd_sc_hd__nand3_2 _17574_ (.A(_07136_),
    .B(_07138_),
    .C(_07151_),
    .Y(_07156_));
 sky130_fd_sc_hd__a21oi_1 _17575_ (.A1(_07155_),
    .A2(_07156_),
    .B1(_07116_),
    .Y(_07157_));
 sky130_fd_sc_hd__nand3_2 _17576_ (.A(_07152_),
    .B(_07153_),
    .C(_07115_),
    .Y(_07158_));
 sky130_fd_sc_hd__nand3_4 _17577_ (.A(_07116_),
    .B(_07155_),
    .C(_07156_),
    .Y(_07159_));
 sky130_fd_sc_hd__o21ai_2 _17578_ (.A1(_06812_),
    .A2(_06827_),
    .B1(_06811_),
    .Y(_07160_));
 sky130_fd_sc_hd__a21oi_2 _17579_ (.A1(_06813_),
    .A2(_06828_),
    .B1(_06810_),
    .Y(_07161_));
 sky130_fd_sc_hd__a21oi_2 _17580_ (.A1(_07158_),
    .A2(_07159_),
    .B1(_07160_),
    .Y(_07162_));
 sky130_fd_sc_hd__a31oi_1 _17581_ (.A1(_07152_),
    .A2(_07153_),
    .A3(_07115_),
    .B1(_07161_),
    .Y(_07163_));
 sky130_fd_sc_hd__and3_1 _17582_ (.A(_07158_),
    .B(_07159_),
    .C(_07160_),
    .X(_07164_));
 sky130_fd_sc_hd__a21oi_1 _17583_ (.A1(_07158_),
    .A2(_07159_),
    .B1(_07161_),
    .Y(_07166_));
 sky130_fd_sc_hd__and3_1 _17584_ (.A(_07158_),
    .B(_07159_),
    .C(_07161_),
    .X(_07167_));
 sky130_fd_sc_hd__a21oi_1 _17585_ (.A1(_07159_),
    .A2(_07163_),
    .B1(_07162_),
    .Y(_07168_));
 sky130_fd_sc_hd__a21o_1 _17586_ (.A1(_07159_),
    .A2(_07163_),
    .B1(_07162_),
    .X(_07169_));
 sky130_fd_sc_hd__o2bb2ai_2 _17587_ (.A1_N(_07113_),
    .A2_N(_07114_),
    .B1(_07162_),
    .B2(_07164_),
    .Y(_07170_));
 sky130_fd_sc_hd__o211ai_2 _17588_ (.A1(_07166_),
    .A2(_07167_),
    .B1(_07113_),
    .C1(_07114_),
    .Y(_07171_));
 sky130_fd_sc_hd__o211ai_2 _17589_ (.A1(_07162_),
    .A2(_07164_),
    .B1(_07113_),
    .C1(_07114_),
    .Y(_07172_));
 sky130_fd_sc_hd__o2bb2ai_2 _17590_ (.A1_N(_07113_),
    .A2_N(_07114_),
    .B1(_07166_),
    .B2(_07167_),
    .Y(_07173_));
 sky130_fd_sc_hd__and3_2 _17591_ (.A(_07026_),
    .B(_07170_),
    .C(_07171_),
    .X(_07174_));
 sky130_fd_sc_hd__nand3_2 _17592_ (.A(_07026_),
    .B(_07170_),
    .C(_07171_),
    .Y(_07175_));
 sky130_fd_sc_hd__o211a_1 _17593_ (.A1(_06794_),
    .A2(_07025_),
    .B1(_07172_),
    .C1(_07173_),
    .X(_07177_));
 sky130_fd_sc_hd__o211ai_4 _17594_ (.A1(_06794_),
    .A2(_07025_),
    .B1(_07172_),
    .C1(_07173_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand3_1 _17595_ (.A(_07024_),
    .B(_07175_),
    .C(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__a21o_1 _17596_ (.A1(_07175_),
    .A2(_07178_),
    .B1(_07024_),
    .X(_07180_));
 sky130_fd_sc_hd__a22o_1 _17597_ (.A1(_07020_),
    .A2(_07022_),
    .B1(_07175_),
    .B2(_07178_),
    .X(_07181_));
 sky130_fd_sc_hd__o211a_1 _17598_ (.A1(_07021_),
    .A2(_07018_),
    .B1(_07020_),
    .C1(_07178_),
    .X(_07182_));
 sky130_fd_sc_hd__o211ai_2 _17599_ (.A1(_07021_),
    .A2(_07018_),
    .B1(_07020_),
    .C1(_07178_),
    .Y(_07183_));
 sky130_fd_sc_hd__o21ai_1 _17600_ (.A1(_07174_),
    .A2(_07183_),
    .B1(_07181_),
    .Y(_07184_));
 sky130_fd_sc_hd__o211ai_4 _17601_ (.A1(_06852_),
    .A2(_06944_),
    .B1(_07179_),
    .C1(_07180_),
    .Y(_07185_));
 sky130_fd_sc_hd__o211a_2 _17602_ (.A1(_07174_),
    .A2(_07183_),
    .B1(_06945_),
    .C1(_07181_),
    .X(_07186_));
 sky130_fd_sc_hd__o211ai_2 _17603_ (.A1(_07174_),
    .A2(_07183_),
    .B1(_06945_),
    .C1(_07181_),
    .Y(_07188_));
 sky130_fd_sc_hd__o211a_1 _17604_ (.A1(_06863_),
    .A2(_06865_),
    .B1(net1),
    .C1(_06877_),
    .X(_07189_));
 sky130_fd_sc_hd__a21oi_2 _17605_ (.A1(_06867_),
    .A2(_06877_),
    .B1(_06875_),
    .Y(_07190_));
 sky130_fd_sc_hd__a21oi_2 _17606_ (.A1(_06646_),
    .A2(_06654_),
    .B1(_06652_),
    .Y(_07191_));
 sky130_fd_sc_hd__a22o_1 _17607_ (.A1(net12),
    .A2(_06865_),
    .B1(_04539_),
    .B2(_06863_),
    .X(_07192_));
 sky130_fd_sc_hd__a32oi_4 _17608_ (.A1(net318),
    .A2(_04452_),
    .A3(_06324_),
    .B1(_06326_),
    .B2(net23),
    .Y(_07193_));
 sky130_fd_sc_hd__a32o_1 _17609_ (.A1(net318),
    .A2(_04452_),
    .A3(_06324_),
    .B1(_06326_),
    .B2(net23),
    .X(_07194_));
 sky130_fd_sc_hd__nor2_1 _17610_ (.A(_03506_),
    .B(_06030_),
    .Y(_07195_));
 sky130_fd_sc_hd__a211oi_4 _17611_ (.A1(_04397_),
    .A2(_04725_),
    .B1(_06028_),
    .C1(_04703_),
    .Y(_07196_));
 sky130_fd_sc_hd__o221ai_4 _17612_ (.A1(_04758_),
    .A2(_06028_),
    .B1(_06030_),
    .B2(_03506_),
    .C1(_07193_),
    .Y(_07197_));
 sky130_fd_sc_hd__o21a_1 _17613_ (.A1(_07195_),
    .A2(_07196_),
    .B1(_07194_),
    .X(_07199_));
 sky130_fd_sc_hd__o21ai_2 _17614_ (.A1(_07195_),
    .A2(_07196_),
    .B1(_07194_),
    .Y(_07200_));
 sky130_fd_sc_hd__nand3b_2 _17615_ (.A_N(_07192_),
    .B(_07197_),
    .C(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__a21bo_1 _17616_ (.A1(_07197_),
    .A2(_07200_),
    .B1_N(_07192_),
    .X(_07202_));
 sky130_fd_sc_hd__a221o_1 _17617_ (.A1(_04539_),
    .A2(_06863_),
    .B1(_06865_),
    .B2(net12),
    .C1(_07199_),
    .X(_07203_));
 sky130_fd_sc_hd__a21oi_1 _17618_ (.A1(_07192_),
    .A2(_07197_),
    .B1(_07199_),
    .Y(_07204_));
 sky130_fd_sc_hd__a21o_1 _17619_ (.A1(_07197_),
    .A2(_07200_),
    .B1(_07192_),
    .X(_07205_));
 sky130_fd_sc_hd__nand3_1 _17620_ (.A(_07192_),
    .B(_07197_),
    .C(_07200_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand3_1 _17621_ (.A(_07191_),
    .B(_07201_),
    .C(_07202_),
    .Y(_07207_));
 sky130_fd_sc_hd__nand3b_2 _17622_ (.A_N(_07191_),
    .B(_07205_),
    .C(_07206_),
    .Y(_07208_));
 sky130_fd_sc_hd__a21oi_1 _17623_ (.A1(_07207_),
    .A2(_07208_),
    .B1(_07190_),
    .Y(_07210_));
 sky130_fd_sc_hd__and3_1 _17624_ (.A(_07190_),
    .B(_07207_),
    .C(_07208_),
    .X(_07211_));
 sky130_fd_sc_hd__o211a_1 _17625_ (.A1(_06875_),
    .A2(_07189_),
    .B1(_07207_),
    .C1(_07208_),
    .X(_07212_));
 sky130_fd_sc_hd__a21boi_1 _17626_ (.A1(_07207_),
    .A2(_07208_),
    .B1_N(_07190_),
    .Y(_07213_));
 sky130_fd_sc_hd__o2bb2ai_1 _17627_ (.A1_N(_06644_),
    .A2_N(_06659_),
    .B1(_07210_),
    .B2(_07211_),
    .Y(_07214_));
 sky130_fd_sc_hd__o211ai_2 _17628_ (.A1(_07212_),
    .A2(_07213_),
    .B1(_06644_),
    .C1(_06659_),
    .Y(_07215_));
 sky130_fd_sc_hd__a21bo_1 _17629_ (.A1(_06334_),
    .A2(_06884_),
    .B1_N(_06883_),
    .X(_07216_));
 sky130_fd_sc_hd__a21o_1 _17630_ (.A1(_07214_),
    .A2(_07215_),
    .B1(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__nand3_1 _17631_ (.A(_07214_),
    .B(_07215_),
    .C(_07216_),
    .Y(_07218_));
 sky130_fd_sc_hd__o31ai_2 _17632_ (.A1(_06337_),
    .A2(_06338_),
    .A3(_06891_),
    .B1(_06894_),
    .Y(_07219_));
 sky130_fd_sc_hd__a21o_1 _17633_ (.A1(_07217_),
    .A2(_07218_),
    .B1(_07219_),
    .X(_07221_));
 sky130_fd_sc_hd__nand3_2 _17634_ (.A(_07217_),
    .B(_07218_),
    .C(_07219_),
    .Y(_07222_));
 sky130_fd_sc_hd__and2b_4 _17635_ (.A_N(net51),
    .B(net52),
    .X(_07223_));
 sky130_fd_sc_hd__nand2b_4 _17636_ (.A_N(net51),
    .B(net52),
    .Y(_07224_));
 sky130_fd_sc_hd__and2b_4 _17637_ (.A_N(net52),
    .B(net51),
    .X(_07225_));
 sky130_fd_sc_hd__nand2b_4 _17638_ (.A_N(net52),
    .B(net51),
    .Y(_07226_));
 sky130_fd_sc_hd__nand2_1 _17639_ (.A(_07224_),
    .B(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__o2111ai_2 _17640_ (.A1(_07223_),
    .A2(_07225_),
    .B1(_07222_),
    .C1(net1),
    .D1(_07221_),
    .Y(_07228_));
 sky130_fd_sc_hd__a22o_1 _17641_ (.A1(_07227_),
    .A2(net1),
    .B1(_07221_),
    .B2(_07222_),
    .X(_07229_));
 sky130_fd_sc_hd__a211oi_2 _17642_ (.A1(_07228_),
    .A2(_07229_),
    .B1(_06696_),
    .C1(_06699_),
    .Y(_07230_));
 sky130_fd_sc_hd__o211a_2 _17643_ (.A1(_06696_),
    .A2(_06699_),
    .B1(_07228_),
    .C1(_07229_),
    .X(_07232_));
 sky130_fd_sc_hd__nor2_1 _17644_ (.A(_07230_),
    .B(_07232_),
    .Y(_07233_));
 sky130_fd_sc_hd__o21a_1 _17645_ (.A1(_07230_),
    .A2(_07232_),
    .B1(_06898_),
    .X(_07234_));
 sky130_fd_sc_hd__nor3_1 _17646_ (.A(_06898_),
    .B(_07230_),
    .C(_07232_),
    .Y(_07235_));
 sky130_fd_sc_hd__nor2_1 _17647_ (.A(_06898_),
    .B(_07233_),
    .Y(_07236_));
 sky130_fd_sc_hd__a2111oi_2 _17648_ (.A1(_06342_),
    .A2(_06345_),
    .B1(_06897_),
    .C1(_07230_),
    .D1(_07232_),
    .Y(_07237_));
 sky130_fd_sc_hd__o2bb2ai_2 _17649_ (.A1_N(_07185_),
    .A2_N(_07188_),
    .B1(_07236_),
    .B2(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__o21a_1 _17650_ (.A1(_07234_),
    .A2(_07235_),
    .B1(_07185_),
    .X(_07239_));
 sky130_fd_sc_hd__o21ai_2 _17651_ (.A1(_07234_),
    .A2(_07235_),
    .B1(_07185_),
    .Y(_07240_));
 sky130_fd_sc_hd__o211ai_2 _17652_ (.A1(_07234_),
    .A2(_07235_),
    .B1(_07185_),
    .C1(_07188_),
    .Y(_07241_));
 sky130_fd_sc_hd__o221a_1 _17653_ (.A1(_06858_),
    .A2(_06915_),
    .B1(_07186_),
    .B2(_07240_),
    .C1(_07238_),
    .X(_07243_));
 sky130_fd_sc_hd__o221ai_4 _17654_ (.A1(_06858_),
    .A2(_06915_),
    .B1(_07186_),
    .B2(_07240_),
    .C1(_07238_),
    .Y(_07244_));
 sky130_fd_sc_hd__a21oi_2 _17655_ (.A1(_07238_),
    .A2(_07241_),
    .B1(_06943_),
    .Y(_07245_));
 sky130_fd_sc_hd__a21o_1 _17656_ (.A1(_07238_),
    .A2(_07241_),
    .B1(_06943_),
    .X(_07246_));
 sky130_fd_sc_hd__o211ai_1 _17657_ (.A1(_06905_),
    .A2(_06941_),
    .B1(_07244_),
    .C1(_07246_),
    .Y(_07247_));
 sky130_fd_sc_hd__o22ai_1 _17658_ (.A1(_06902_),
    .A2(_06940_),
    .B1(_07243_),
    .B2(_07245_),
    .Y(_07248_));
 sky130_fd_sc_hd__o22ai_2 _17659_ (.A1(_06905_),
    .A2(_06941_),
    .B1(_07243_),
    .B2(_07245_),
    .Y(_07249_));
 sky130_fd_sc_hd__o211ai_2 _17660_ (.A1(_06902_),
    .A2(_06940_),
    .B1(_07244_),
    .C1(_07246_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_1 _17661_ (.A(_07247_),
    .B(_07248_),
    .Y(_07251_));
 sky130_fd_sc_hd__nand3_1 _17662_ (.A(_06939_),
    .B(_07249_),
    .C(_07250_),
    .Y(_07252_));
 sky130_fd_sc_hd__a22oi_1 _17663_ (.A1(_06921_),
    .A2(_06922_),
    .B1(_07249_),
    .B2(_07250_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand3_1 _17664_ (.A(_07248_),
    .B(_06938_),
    .C(_07247_),
    .Y(_07255_));
 sky130_fd_sc_hd__a21boi_1 _17665_ (.A1(_07252_),
    .A2(_07255_),
    .B1_N(_06930_),
    .Y(_07256_));
 sky130_fd_sc_hd__a31oi_1 _17666_ (.A1(_06939_),
    .A2(_07249_),
    .A3(_07250_),
    .B1(_06930_),
    .Y(_07257_));
 sky130_fd_sc_hd__a21oi_1 _17667_ (.A1(_07257_),
    .A2(_07255_),
    .B1(_07256_),
    .Y(_07258_));
 sky130_fd_sc_hd__a22oi_1 _17668_ (.A1(_06930_),
    .A2(_06932_),
    .B1(_06937_),
    .B2(_06934_),
    .Y(_07259_));
 sky130_fd_sc_hd__xnor2_1 _17669_ (.A(_07258_),
    .B(_07259_),
    .Y(net84));
 sky130_fd_sc_hd__o21a_1 _17670_ (.A1(_06902_),
    .A2(_06940_),
    .B1(_07244_),
    .X(_07260_));
 sky130_fd_sc_hd__o21ai_1 _17671_ (.A1(_06942_),
    .A2(_07245_),
    .B1(_07244_),
    .Y(_07261_));
 sky130_fd_sc_hd__inv_2 _17672_ (.A(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__a21boi_1 _17673_ (.A1(_07215_),
    .A2(_07216_),
    .B1_N(_07214_),
    .Y(_07264_));
 sky130_fd_sc_hd__a32o_1 _17674_ (.A1(_06863_),
    .A2(_04452_),
    .A3(net318),
    .B1(net23),
    .B2(_06865_),
    .X(_07265_));
 sky130_fd_sc_hd__a32oi_2 _17675_ (.A1(net313),
    .A2(_04747_),
    .A3(_06324_),
    .B1(_06326_),
    .B2(net26),
    .Y(_07266_));
 sky130_fd_sc_hd__a32o_1 _17676_ (.A1(net313),
    .A2(_04747_),
    .A3(_06324_),
    .B1(_06326_),
    .B2(net26),
    .X(_07267_));
 sky130_fd_sc_hd__nor2_1 _17677_ (.A(_03616_),
    .B(_06030_),
    .Y(_07268_));
 sky130_fd_sc_hd__or3b_1 _17678_ (.A(_03616_),
    .B(net49),
    .C_N(net48),
    .X(_07269_));
 sky130_fd_sc_hd__a31o_1 _17679_ (.A1(net266),
    .A2(net302),
    .A3(_06026_),
    .B1(_07268_),
    .X(_07270_));
 sky130_fd_sc_hd__and2_1 _17680_ (.A(_07267_),
    .B(_07270_),
    .X(_07271_));
 sky130_fd_sc_hd__nand2_1 _17681_ (.A(_07267_),
    .B(_07270_),
    .Y(_07272_));
 sky130_fd_sc_hd__o221ai_2 _17682_ (.A1(_05020_),
    .A2(_06028_),
    .B1(_06030_),
    .B2(_03616_),
    .C1(_07266_),
    .Y(_07273_));
 sky130_fd_sc_hd__nand2_1 _17683_ (.A(_07270_),
    .B(_07266_),
    .Y(_07275_));
 sky130_fd_sc_hd__o211ai_1 _17684_ (.A1(_05020_),
    .A2(_06028_),
    .B1(_07267_),
    .C1(_07269_),
    .Y(_07276_));
 sky130_fd_sc_hd__nand3b_2 _17685_ (.A_N(_07265_),
    .B(_07275_),
    .C(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__nand3_2 _17686_ (.A(_07265_),
    .B(_07272_),
    .C(_07273_),
    .Y(_07278_));
 sky130_fd_sc_hd__inv_2 _17687_ (.A(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__o21a_1 _17688_ (.A1(_06980_),
    .A2(_06983_),
    .B1(_06977_),
    .X(_07280_));
 sky130_fd_sc_hd__a21oi_1 _17689_ (.A1(_06980_),
    .A2(_06983_),
    .B1(_06977_),
    .Y(_07281_));
 sky130_fd_sc_hd__o21bai_1 _17690_ (.A1(_06977_),
    .A2(_06985_),
    .B1_N(_06984_),
    .Y(_07282_));
 sky130_fd_sc_hd__o2bb2a_1 _17691_ (.A1_N(_07277_),
    .A2_N(_07278_),
    .B1(_07280_),
    .B2(_06985_),
    .X(_07283_));
 sky130_fd_sc_hd__o2bb2ai_1 _17692_ (.A1_N(_07277_),
    .A2_N(_07278_),
    .B1(_07280_),
    .B2(_06985_),
    .Y(_07284_));
 sky130_fd_sc_hd__o211ai_2 _17693_ (.A1(_06984_),
    .A2(_07281_),
    .B1(_07278_),
    .C1(_07277_),
    .Y(_07286_));
 sky130_fd_sc_hd__a31oi_1 _17694_ (.A1(_07282_),
    .A2(_07278_),
    .A3(_07277_),
    .B1(_07204_),
    .Y(_07287_));
 sky130_fd_sc_hd__a31o_1 _17695_ (.A1(_07282_),
    .A2(_07278_),
    .A3(_07277_),
    .B1(_07204_),
    .X(_07288_));
 sky130_fd_sc_hd__a22oi_1 _17696_ (.A1(_07197_),
    .A2(_07203_),
    .B1(_07284_),
    .B2(_07286_),
    .Y(_07289_));
 sky130_fd_sc_hd__a22o_1 _17697_ (.A1(_07197_),
    .A2(_07203_),
    .B1(_07284_),
    .B2(_07286_),
    .X(_07290_));
 sky130_fd_sc_hd__a21oi_1 _17698_ (.A1(_07284_),
    .A2(_07287_),
    .B1(_07289_),
    .Y(_07291_));
 sky130_fd_sc_hd__o21ai_1 _17699_ (.A1(_07283_),
    .A2(_07288_),
    .B1(_07290_),
    .Y(_07292_));
 sky130_fd_sc_hd__a32oi_2 _17700_ (.A1(_06989_),
    .A2(_07000_),
    .A3(_07002_),
    .B1(_06987_),
    .B2(_06986_),
    .Y(_07293_));
 sky130_fd_sc_hd__nand2_1 _17701_ (.A(_06988_),
    .B(_07003_),
    .Y(_07294_));
 sky130_fd_sc_hd__o21ai_1 _17702_ (.A1(_07004_),
    .A2(_07293_),
    .B1(_07292_),
    .Y(_07295_));
 sky130_fd_sc_hd__nand3_1 _17703_ (.A(_07291_),
    .B(_07294_),
    .C(_07005_),
    .Y(_07297_));
 sky130_fd_sc_hd__a32oi_4 _17704_ (.A1(_07191_),
    .A2(_07201_),
    .A3(_07202_),
    .B1(_07208_),
    .B2(_07190_),
    .Y(_07298_));
 sky130_fd_sc_hd__a21oi_1 _17705_ (.A1(_07295_),
    .A2(_07297_),
    .B1(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__a21o_1 _17706_ (.A1(_07295_),
    .A2(_07297_),
    .B1(_07298_),
    .X(_07300_));
 sky130_fd_sc_hd__and3_1 _17707_ (.A(_07295_),
    .B(_07297_),
    .C(_07298_),
    .X(_07301_));
 sky130_fd_sc_hd__nand3_1 _17708_ (.A(_07295_),
    .B(_07297_),
    .C(_07298_),
    .Y(_07302_));
 sky130_fd_sc_hd__o21ai_1 _17709_ (.A1(_07299_),
    .A2(_07301_),
    .B1(_07264_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand3b_1 _17710_ (.A_N(_07264_),
    .B(_07300_),
    .C(_07302_),
    .Y(_07304_));
 sky130_fd_sc_hd__nor2_8 _17711_ (.A(net52),
    .B(_04234_),
    .Y(_07305_));
 sky130_fd_sc_hd__nand2b_4 _17712_ (.A_N(net52),
    .B(net53),
    .Y(_07306_));
 sky130_fd_sc_hd__and2_4 _17713_ (.A(_04234_),
    .B(net52),
    .X(_07308_));
 sky130_fd_sc_hd__o21a_1 _17714_ (.A1(_07305_),
    .A2(_07308_),
    .B1(net1),
    .X(_07309_));
 sky130_fd_sc_hd__a22o_1 _17715_ (.A1(net12),
    .A2(_07225_),
    .B1(_04539_),
    .B2(_07223_),
    .X(_07310_));
 sky130_fd_sc_hd__o211a_1 _17716_ (.A1(_07305_),
    .A2(_07308_),
    .B1(net1),
    .C1(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__nor2_1 _17717_ (.A(_07310_),
    .B(_07309_),
    .Y(_07312_));
 sky130_fd_sc_hd__nor2_1 _17718_ (.A(_07311_),
    .B(_07312_),
    .Y(_07313_));
 sky130_fd_sc_hd__a21o_1 _17719_ (.A1(_07303_),
    .A2(_07304_),
    .B1(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__nand3_1 _17720_ (.A(_07303_),
    .B(_07304_),
    .C(_07313_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand2_1 _17721_ (.A(_07314_),
    .B(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__a21oi_1 _17722_ (.A1(_07017_),
    .A2(_07021_),
    .B1(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__a21o_1 _17723_ (.A1(_07017_),
    .A2(_07022_),
    .B1(_07316_),
    .X(_07319_));
 sky130_fd_sc_hd__nand3_2 _17724_ (.A(_07017_),
    .B(_07022_),
    .C(_07316_),
    .Y(_07320_));
 sky130_fd_sc_hd__o211ai_1 _17725_ (.A1(_07223_),
    .A2(_07225_),
    .B1(net1),
    .C1(_07221_),
    .Y(_07321_));
 sky130_fd_sc_hd__and2_1 _17726_ (.A(_07222_),
    .B(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__a21boi_4 _17727_ (.A1(_07319_),
    .A2(_07320_),
    .B1_N(_07322_),
    .Y(_07323_));
 sky130_fd_sc_hd__a21oi_1 _17728_ (.A1(_07222_),
    .A2(_07321_),
    .B1(_07317_),
    .Y(_07324_));
 sky130_fd_sc_hd__and3b_1 _17729_ (.A_N(_07322_),
    .B(_07320_),
    .C(_07319_),
    .X(_07325_));
 sky130_fd_sc_hd__a21oi_2 _17730_ (.A1(_07324_),
    .A2(_07320_),
    .B1(_07323_),
    .Y(_07326_));
 sky130_fd_sc_hd__a32oi_1 _17731_ (.A1(_07026_),
    .A2(_07170_),
    .A3(_07171_),
    .B1(_07022_),
    .B2(_07020_),
    .Y(_07327_));
 sky130_fd_sc_hd__a21boi_2 _17732_ (.A1(_06966_),
    .A2(_06967_),
    .B1_N(_06965_),
    .Y(_07328_));
 sky130_fd_sc_hd__o21a_1 _17733_ (.A1(_06949_),
    .A2(_06960_),
    .B1(_06959_),
    .X(_07330_));
 sky130_fd_sc_hd__o21ai_1 _17734_ (.A1(_06949_),
    .A2(_06960_),
    .B1(_06959_),
    .Y(_07331_));
 sky130_fd_sc_hd__or3_1 _17735_ (.A(net39),
    .B(_04037_),
    .C(_04015_),
    .X(_07332_));
 sky130_fd_sc_hd__o211ai_1 _17736_ (.A1(net254),
    .A2(_00646_),
    .B1(net285),
    .C1(_00625_),
    .Y(_07333_));
 sky130_fd_sc_hd__a32oi_4 _17737_ (.A1(_00625_),
    .A2(_00657_),
    .A3(net285),
    .B1(_03726_),
    .B2(net5),
    .Y(_07334_));
 sky130_fd_sc_hd__nor2_1 _17738_ (.A(_04004_),
    .B(_04218_),
    .Y(_07335_));
 sky130_fd_sc_hd__o311a_1 _17739_ (.A1(net3),
    .A2(_09665_),
    .A3(_12988_),
    .B1(net281),
    .C1(net234),
    .X(_07336_));
 sky130_fd_sc_hd__a31oi_2 _17740_ (.A1(net234),
    .A2(net251),
    .A3(net281),
    .B1(_07335_),
    .Y(_07337_));
 sky130_fd_sc_hd__nand2_1 _17741_ (.A(_07334_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__o2bb2ai_2 _17742_ (.A1_N(_07332_),
    .A2_N(_07333_),
    .B1(_07335_),
    .B2(_07336_),
    .Y(_07339_));
 sky130_fd_sc_hd__a32o_1 _17743_ (.A1(_11354_),
    .A2(net254),
    .A3(net280),
    .B1(_04269_),
    .B2(net3),
    .X(_07341_));
 sky130_fd_sc_hd__a21oi_1 _17744_ (.A1(_07338_),
    .A2(_07339_),
    .B1(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__a21o_1 _17745_ (.A1(_07338_),
    .A2(_07339_),
    .B1(_07341_),
    .X(_07343_));
 sky130_fd_sc_hd__and3_1 _17746_ (.A(_07338_),
    .B(_07339_),
    .C(_07341_),
    .X(_07344_));
 sky130_fd_sc_hd__nand3_2 _17747_ (.A(_07338_),
    .B(_07339_),
    .C(_07341_),
    .Y(_07345_));
 sky130_fd_sc_hd__a21o_1 _17748_ (.A1(_07139_),
    .A2(_07146_),
    .B1(_07147_),
    .X(_07346_));
 sky130_fd_sc_hd__a21oi_1 _17749_ (.A1(_07343_),
    .A2(_07345_),
    .B1(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__o21bai_1 _17750_ (.A1(_07342_),
    .A2(_07344_),
    .B1_N(_07346_),
    .Y(_07348_));
 sky130_fd_sc_hd__nand2_1 _17751_ (.A(_07343_),
    .B(_07346_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand3_1 _17752_ (.A(_07343_),
    .B(_07346_),
    .C(_07345_),
    .Y(_07350_));
 sky130_fd_sc_hd__a21oi_2 _17753_ (.A1(_07348_),
    .A2(_07350_),
    .B1(_07331_),
    .Y(_07352_));
 sky130_fd_sc_hd__a21oi_1 _17754_ (.A1(_06959_),
    .A2(_06962_),
    .B1(_07347_),
    .Y(_07353_));
 sky130_fd_sc_hd__and3_1 _17755_ (.A(_07331_),
    .B(_07348_),
    .C(_07350_),
    .X(_07354_));
 sky130_fd_sc_hd__o21ai_4 _17756_ (.A1(_07352_),
    .A2(_07354_),
    .B1(_07328_),
    .Y(_07355_));
 sky130_fd_sc_hd__a211o_2 _17757_ (.A1(_07353_),
    .A2(_07350_),
    .B1(_07328_),
    .C1(_07352_),
    .X(_07356_));
 sky130_fd_sc_hd__inv_2 _17758_ (.A(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__a32o_1 _17759_ (.A1(_07242_),
    .A2(net257),
    .A3(_04985_),
    .B1(_04988_),
    .B2(net31),
    .X(_07358_));
 sky130_fd_sc_hd__or3b_1 _17760_ (.A(_03960_),
    .B(net42),
    .C_N(net41),
    .X(_07359_));
 sky130_fd_sc_hd__o211ai_4 _17761_ (.A1(net260),
    .A2(_09665_),
    .B1(net279),
    .C1(_09698_),
    .Y(_07360_));
 sky130_fd_sc_hd__or3b_2 _17762_ (.A(_03949_),
    .B(net43),
    .C_N(net42),
    .X(_07361_));
 sky130_fd_sc_hd__o211ai_4 _17763_ (.A1(net260),
    .A2(_08656_),
    .B1(net243),
    .C1(_08700_),
    .Y(_07363_));
 sky130_fd_sc_hd__o2111a_1 _17764_ (.A1(_03960_),
    .A2(_04483_),
    .B1(_07360_),
    .C1(_07361_),
    .D1(_07363_),
    .X(_07364_));
 sky130_fd_sc_hd__o2111ai_2 _17765_ (.A1(_03960_),
    .A2(_04483_),
    .B1(_07360_),
    .C1(_07361_),
    .D1(_07363_),
    .Y(_07365_));
 sky130_fd_sc_hd__a22oi_2 _17766_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07361_),
    .B2(_07363_),
    .Y(_07366_));
 sky130_fd_sc_hd__a22o_1 _17767_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07361_),
    .B2(_07363_),
    .X(_07367_));
 sky130_fd_sc_hd__o21bai_2 _17768_ (.A1(_07364_),
    .A2(_07366_),
    .B1_N(_07358_),
    .Y(_07368_));
 sky130_fd_sc_hd__nand3_2 _17769_ (.A(_07358_),
    .B(_07365_),
    .C(_07367_),
    .Y(_07369_));
 sky130_fd_sc_hd__a21o_1 _17770_ (.A1(_06991_),
    .A2(_06999_),
    .B1(_06997_),
    .X(_07370_));
 sky130_fd_sc_hd__a21oi_1 _17771_ (.A1(_07368_),
    .A2(_07369_),
    .B1(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__a21o_1 _17772_ (.A1(_07368_),
    .A2(_07369_),
    .B1(_07370_),
    .X(_07372_));
 sky130_fd_sc_hd__nand3_1 _17773_ (.A(_07368_),
    .B(_07369_),
    .C(_07370_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand2_1 _17774_ (.A(_07372_),
    .B(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__a32o_1 _17775_ (.A1(_05414_),
    .A2(_05446_),
    .A3(net275),
    .B1(_05765_),
    .B2(net28),
    .X(_07376_));
 sky130_fd_sc_hd__a32oi_4 _17776_ (.A1(_05841_),
    .A2(net265),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net29),
    .Y(_07377_));
 sky130_fd_sc_hd__a32o_1 _17777_ (.A1(_05841_),
    .A2(net265),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net29),
    .X(_07378_));
 sky130_fd_sc_hd__or3_1 _17778_ (.A(net46),
    .B(_04124_),
    .C(_03916_),
    .X(_07379_));
 sky130_fd_sc_hd__o2111ai_4 _17779_ (.A1(_04747_),
    .A2(net264),
    .B1(net46),
    .C1(_06486_),
    .D1(_04124_),
    .Y(_07380_));
 sky130_fd_sc_hd__a32o_1 _17780_ (.A1(_06486_),
    .A2(net260),
    .A3(net276),
    .B1(_05228_),
    .B2(net30),
    .X(_07381_));
 sky130_fd_sc_hd__a21oi_1 _17781_ (.A1(_07379_),
    .A2(_07380_),
    .B1(_07377_),
    .Y(_07382_));
 sky130_fd_sc_hd__a21o_1 _17782_ (.A1(_07379_),
    .A2(_07380_),
    .B1(_07377_),
    .X(_07383_));
 sky130_fd_sc_hd__o311a_1 _17783_ (.A1(_03916_),
    .A2(_04124_),
    .A3(net46),
    .B1(_07380_),
    .C1(_07377_),
    .X(_07385_));
 sky130_fd_sc_hd__o211ai_2 _17784_ (.A1(_03916_),
    .A2(_05229_),
    .B1(_07380_),
    .C1(_07377_),
    .Y(_07386_));
 sky130_fd_sc_hd__a21o_1 _17785_ (.A1(_07383_),
    .A2(_07386_),
    .B1(_07376_),
    .X(_07387_));
 sky130_fd_sc_hd__nand3_1 _17786_ (.A(_07376_),
    .B(_07383_),
    .C(_07386_),
    .Y(_07388_));
 sky130_fd_sc_hd__o21ai_1 _17787_ (.A1(_07382_),
    .A2(_07385_),
    .B1(_07376_),
    .Y(_07389_));
 sky130_fd_sc_hd__nand3b_1 _17788_ (.A_N(_07376_),
    .B(_07383_),
    .C(_07386_),
    .Y(_07390_));
 sky130_fd_sc_hd__nand2_1 _17789_ (.A(_07389_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__and3_1 _17790_ (.A(_07372_),
    .B(_07374_),
    .C(_07391_),
    .X(_07392_));
 sky130_fd_sc_hd__and3_1 _17791_ (.A(_07375_),
    .B(_07389_),
    .C(_07390_),
    .X(_07393_));
 sky130_fd_sc_hd__and4_1 _17792_ (.A(_07372_),
    .B(_07374_),
    .C(_07389_),
    .D(_07390_),
    .X(_07394_));
 sky130_fd_sc_hd__and3_1 _17793_ (.A(_07375_),
    .B(_07387_),
    .C(_07388_),
    .X(_07396_));
 sky130_fd_sc_hd__nor2_1 _17794_ (.A(_07392_),
    .B(_07393_),
    .Y(_07397_));
 sky130_fd_sc_hd__o211ai_2 _17795_ (.A1(_07392_),
    .A2(_07393_),
    .B1(_07355_),
    .C1(_07356_),
    .Y(_07398_));
 sky130_fd_sc_hd__o2bb2ai_1 _17796_ (.A1_N(_07355_),
    .A2_N(_07356_),
    .B1(_07394_),
    .B2(_07396_),
    .Y(_07399_));
 sky130_fd_sc_hd__o2bb2ai_2 _17797_ (.A1_N(_07355_),
    .A2_N(_07356_),
    .B1(_07392_),
    .B2(_07393_),
    .Y(_07400_));
 sky130_fd_sc_hd__o21a_1 _17798_ (.A1(_07394_),
    .A2(_07396_),
    .B1(_07355_),
    .X(_07401_));
 sky130_fd_sc_hd__o211ai_2 _17799_ (.A1(_07394_),
    .A2(_07396_),
    .B1(_07355_),
    .C1(_07356_),
    .Y(_07402_));
 sky130_fd_sc_hd__o21ai_2 _17800_ (.A1(_07161_),
    .A2(_07157_),
    .B1(_07159_),
    .Y(_07403_));
 sky130_fd_sc_hd__a21boi_2 _17801_ (.A1(_07158_),
    .A2(_07160_),
    .B1_N(_07159_),
    .Y(_07404_));
 sky130_fd_sc_hd__nand3_1 _17802_ (.A(_07398_),
    .B(_07399_),
    .C(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__nand3_4 _17803_ (.A(_07400_),
    .B(_07403_),
    .C(_07402_),
    .Y(_07407_));
 sky130_fd_sc_hd__a21oi_1 _17804_ (.A1(_07405_),
    .A2(_07407_),
    .B1(_07011_),
    .Y(_07408_));
 sky130_fd_sc_hd__a31oi_2 _17805_ (.A1(_07398_),
    .A2(_07399_),
    .A3(_07404_),
    .B1(_07013_),
    .Y(_07409_));
 sky130_fd_sc_hd__nand3_1 _17806_ (.A(_07405_),
    .B(_07407_),
    .C(_07011_),
    .Y(_07410_));
 sky130_fd_sc_hd__a21oi_2 _17807_ (.A1(_07407_),
    .A2(_07409_),
    .B1(_07408_),
    .Y(_07411_));
 sky130_fd_sc_hd__a21o_1 _17808_ (.A1(_07407_),
    .A2(_07409_),
    .B1(_07408_),
    .X(_07412_));
 sky130_fd_sc_hd__o21ai_1 _17809_ (.A1(_07027_),
    .A2(_07043_),
    .B1(_07046_),
    .Y(_07413_));
 sky130_fd_sc_hd__a32o_2 _17810_ (.A1(net223),
    .A2(net252),
    .A3(net188),
    .B1(_11793_),
    .B2(net9),
    .X(_07414_));
 sky130_fd_sc_hd__a31oi_2 _17811_ (.A1(_11420_),
    .A2(net282),
    .A3(_04556_),
    .B1(_10324_),
    .Y(_07415_));
 sky130_fd_sc_hd__a22oi_4 _17812_ (.A1(net10),
    .A2(_10335_),
    .B1(_07415_),
    .B2(net219),
    .Y(_07416_));
 sky130_fd_sc_hd__o221ai_2 _17813_ (.A1(net232),
    .A2(_04787_),
    .B1(_04091_),
    .B2(_04558_),
    .C1(net291),
    .Y(_07418_));
 sky130_fd_sc_hd__or3b_1 _17814_ (.A(net64),
    .B(_04091_),
    .C_N(net63),
    .X(_07419_));
 sky130_fd_sc_hd__a21oi_2 _17815_ (.A1(_07418_),
    .A2(_07419_),
    .B1(_07416_),
    .Y(_07420_));
 sky130_fd_sc_hd__a21o_1 _17816_ (.A1(_07418_),
    .A2(_07419_),
    .B1(_07416_),
    .X(_07421_));
 sky130_fd_sc_hd__o221a_1 _17817_ (.A1(_04091_),
    .A2(_08283_),
    .B1(_04793_),
    .B2(_08261_),
    .C1(_07416_),
    .X(_07422_));
 sky130_fd_sc_hd__o221ai_4 _17818_ (.A1(_04091_),
    .A2(_08283_),
    .B1(_04793_),
    .B2(_08261_),
    .C1(_07416_),
    .Y(_07423_));
 sky130_fd_sc_hd__o21bai_4 _17819_ (.A1(_07420_),
    .A2(_07422_),
    .B1_N(_07414_),
    .Y(_07424_));
 sky130_fd_sc_hd__nand3_4 _17820_ (.A(_07414_),
    .B(_07421_),
    .C(_07423_),
    .Y(_07425_));
 sky130_fd_sc_hd__o21a_1 _17821_ (.A1(_07123_),
    .A2(_07126_),
    .B1(_07119_),
    .X(_07426_));
 sky130_fd_sc_hd__o21ai_1 _17822_ (.A1(_07118_),
    .A2(_07129_),
    .B1(_07128_),
    .Y(_07427_));
 sky130_fd_sc_hd__a21oi_4 _17823_ (.A1(_07424_),
    .A2(_07425_),
    .B1(_07427_),
    .Y(_07429_));
 sky130_fd_sc_hd__o211a_1 _17824_ (.A1(_07127_),
    .A2(_07426_),
    .B1(_07425_),
    .C1(_07424_),
    .X(_07430_));
 sky130_fd_sc_hd__o211ai_4 _17825_ (.A1(_07127_),
    .A2(_07426_),
    .B1(_07425_),
    .C1(_07424_),
    .Y(_07431_));
 sky130_fd_sc_hd__a32o_1 _17826_ (.A1(_02421_),
    .A2(net249),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net6),
    .X(_07432_));
 sky130_fd_sc_hd__nor2_1 _17827_ (.A(_04059_),
    .B(_12363_),
    .Y(_07433_));
 sky130_fd_sc_hd__a31oi_1 _17828_ (.A1(net228),
    .A2(_12330_),
    .A3(net230),
    .B1(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__a31o_1 _17829_ (.A1(net228),
    .A2(_12330_),
    .A3(net230),
    .B1(_07433_),
    .X(_07435_));
 sky130_fd_sc_hd__o31a_1 _17830_ (.A1(_04747_),
    .A2(net264),
    .A3(_03956_),
    .B1(_01293_),
    .X(_07436_));
 sky130_fd_sc_hd__a22oi_1 _17831_ (.A1(net7),
    .A2(_01315_),
    .B1(_07436_),
    .B2(_03952_),
    .Y(_07437_));
 sky130_fd_sc_hd__o2bb2ai_1 _17832_ (.A1_N(_03952_),
    .A2_N(_07436_),
    .B1(_04048_),
    .B2(_01326_),
    .Y(_07438_));
 sky130_fd_sc_hd__nor2_1 _17833_ (.A(_07434_),
    .B(_07437_),
    .Y(_07440_));
 sky130_fd_sc_hd__nand2_1 _17834_ (.A(_07435_),
    .B(_07438_),
    .Y(_07441_));
 sky130_fd_sc_hd__nand2_1 _17835_ (.A(_07434_),
    .B(_07437_),
    .Y(_07442_));
 sky130_fd_sc_hd__nand2_1 _17836_ (.A(_07441_),
    .B(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__a221o_1 _17837_ (.A1(_02464_),
    .A2(_02858_),
    .B1(_02880_),
    .B2(net6),
    .C1(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__nand2_2 _17838_ (.A(_07432_),
    .B(_07443_),
    .Y(_07445_));
 sky130_fd_sc_hd__xnor2_1 _17839_ (.A(_07432_),
    .B(_07443_),
    .Y(_07446_));
 sky130_fd_sc_hd__o21bai_1 _17840_ (.A1(_07429_),
    .A2(_07430_),
    .B1_N(_07446_),
    .Y(_07447_));
 sky130_fd_sc_hd__nand3b_1 _17841_ (.A_N(_07429_),
    .B(_07431_),
    .C(_07446_),
    .Y(_07448_));
 sky130_fd_sc_hd__nand4b_2 _17842_ (.A_N(_07429_),
    .B(_07431_),
    .C(_07444_),
    .D(_07445_),
    .Y(_07449_));
 sky130_fd_sc_hd__o21ai_1 _17843_ (.A1(_07429_),
    .A2(_07430_),
    .B1(_07446_),
    .Y(_07451_));
 sky130_fd_sc_hd__nand4_4 _17844_ (.A(_07046_),
    .B(_07048_),
    .C(_07449_),
    .D(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__nand3_2 _17845_ (.A(_07413_),
    .B(_07447_),
    .C(_07448_),
    .Y(_07453_));
 sky130_fd_sc_hd__a21oi_1 _17846_ (.A1(_07136_),
    .A2(_07151_),
    .B1(_07137_),
    .Y(_07454_));
 sky130_fd_sc_hd__a221oi_2 _17847_ (.A1(_07136_),
    .A2(_07151_),
    .B1(_07452_),
    .B2(_07453_),
    .C1(_07137_),
    .Y(_07455_));
 sky130_fd_sc_hd__and3b_1 _17848_ (.A_N(_07454_),
    .B(_07453_),
    .C(_07452_),
    .X(_07456_));
 sky130_fd_sc_hd__and3_1 _17849_ (.A(_07452_),
    .B(_07453_),
    .C(_07454_),
    .X(_07457_));
 sky130_fd_sc_hd__a21oi_2 _17850_ (.A1(_07452_),
    .A2(_07453_),
    .B1(_07454_),
    .Y(_07458_));
 sky130_fd_sc_hd__a21oi_2 _17851_ (.A1(_07037_),
    .A2(_07038_),
    .B1(_07033_),
    .Y(_07459_));
 sky130_fd_sc_hd__o21ai_2 _17852_ (.A1(_07052_),
    .A2(_07060_),
    .B1(_07059_),
    .Y(_07460_));
 sky130_fd_sc_hd__nand3_4 _17853_ (.A(net181),
    .B(net180),
    .C(net292),
    .Y(_07462_));
 sky130_fd_sc_hd__or3b_4 _17854_ (.A(net62),
    .B(_04135_),
    .C_N(net61),
    .X(_07463_));
 sky130_fd_sc_hd__o211ai_4 _17855_ (.A1(net185),
    .A2(_05551_),
    .B1(_05688_),
    .C1(_05549_),
    .Y(_07464_));
 sky130_fd_sc_hd__or3b_2 _17856_ (.A(net61),
    .B(_04146_),
    .C_N(net60),
    .X(_07465_));
 sky130_fd_sc_hd__a22oi_4 _17857_ (.A1(_07462_),
    .A2(_07463_),
    .B1(_07464_),
    .B2(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__a22o_4 _17858_ (.A1(_07462_),
    .A2(_07463_),
    .B1(_07464_),
    .B2(_07465_),
    .X(_07467_));
 sky130_fd_sc_hd__o2111a_2 _17859_ (.A1(_04146_),
    .A2(_05720_),
    .B1(_07462_),
    .C1(_07463_),
    .D1(_07464_),
    .X(_07468_));
 sky130_fd_sc_hd__o2111ai_4 _17860_ (.A1(_04146_),
    .A2(_05720_),
    .B1(_07462_),
    .C1(_07463_),
    .D1(_07464_),
    .Y(_07469_));
 sky130_fd_sc_hd__a32o_2 _17861_ (.A1(net212),
    .A2(net183),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net13),
    .X(_07470_));
 sky130_fd_sc_hd__o21bai_4 _17862_ (.A1(_07466_),
    .A2(_07468_),
    .B1_N(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nand2_2 _17863_ (.A(_07467_),
    .B(_07470_),
    .Y(_07473_));
 sky130_fd_sc_hd__nand3_4 _17864_ (.A(_07467_),
    .B(_07469_),
    .C(_07470_),
    .Y(_07474_));
 sky130_fd_sc_hd__a21oi_2 _17865_ (.A1(_07471_),
    .A2(_07474_),
    .B1(_07460_),
    .Y(_07475_));
 sky130_fd_sc_hd__a21o_1 _17866_ (.A1(_07471_),
    .A2(_07474_),
    .B1(_07460_),
    .X(_07476_));
 sky130_fd_sc_hd__o211a_1 _17867_ (.A1(_07468_),
    .A2(_07473_),
    .B1(_07471_),
    .C1(_07460_),
    .X(_07477_));
 sky130_fd_sc_hd__o221ai_4 _17868_ (.A1(_07468_),
    .A2(_07473_),
    .B1(_07058_),
    .B2(_07065_),
    .C1(_07471_),
    .Y(_07478_));
 sky130_fd_sc_hd__o21ai_4 _17869_ (.A1(_07475_),
    .A2(_07477_),
    .B1(_07459_),
    .Y(_07479_));
 sky130_fd_sc_hd__nand3b_4 _17870_ (.A_N(_07459_),
    .B(_07476_),
    .C(_07478_),
    .Y(_07480_));
 sky130_fd_sc_hd__nand2_2 _17871_ (.A(_07479_),
    .B(_07480_),
    .Y(_07481_));
 sky130_fd_sc_hd__o22ai_4 _17872_ (.A1(_04157_),
    .A2(_05260_),
    .B1(net155),
    .B2(_05238_),
    .Y(_07482_));
 sky130_fd_sc_hd__a32oi_4 _17873_ (.A1(_06219_),
    .A2(_06221_),
    .A3(_04889_),
    .B1(_04911_),
    .B2(net17),
    .Y(_07484_));
 sky130_fd_sc_hd__nor2_1 _17874_ (.A(_04179_),
    .B(net316),
    .Y(_07485_));
 sky130_fd_sc_hd__a31oi_4 _17875_ (.A1(net199),
    .A2(net172),
    .A3(_04627_),
    .B1(_07485_),
    .Y(_07486_));
 sky130_fd_sc_hd__nor2_2 _17876_ (.A(_07484_),
    .B(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__o221a_2 _17877_ (.A1(_04179_),
    .A2(net316),
    .B1(_06454_),
    .B2(_04638_),
    .C1(_07484_),
    .X(_07488_));
 sky130_fd_sc_hd__nand2_1 _17878_ (.A(_07484_),
    .B(_07486_),
    .Y(_07489_));
 sky130_fd_sc_hd__o21ba_2 _17879_ (.A1(_07487_),
    .A2(_07488_),
    .B1_N(_07482_),
    .X(_07490_));
 sky130_fd_sc_hd__o21bai_2 _17880_ (.A1(_07487_),
    .A2(_07488_),
    .B1_N(_07482_),
    .Y(_07491_));
 sky130_fd_sc_hd__o21ai_4 _17881_ (.A1(_07484_),
    .A2(_07486_),
    .B1(_07482_),
    .Y(_07492_));
 sky130_fd_sc_hd__a21oi_4 _17882_ (.A1(_07484_),
    .A2(_07486_),
    .B1(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__o21ai_2 _17883_ (.A1(_07488_),
    .A2(_07492_),
    .B1(_07491_),
    .Y(_07495_));
 sky130_fd_sc_hd__nand2_1 _17884_ (.A(net171),
    .B(_04342_),
    .Y(_07496_));
 sky130_fd_sc_hd__o22ai_4 _17885_ (.A1(_04201_),
    .A2(_04375_),
    .B1(_06756_),
    .B2(_07496_),
    .Y(_07497_));
 sky130_fd_sc_hd__a41oi_4 _17886_ (.A1(_11420_),
    .A2(net284),
    .A3(_05926_),
    .A4(net270),
    .B1(_04223_),
    .Y(_07498_));
 sky130_fd_sc_hd__a41o_4 _17887_ (.A1(_06519_),
    .A2(_03955_),
    .A3(_05926_),
    .A4(net271),
    .B1(_04223_),
    .X(_07499_));
 sky130_fd_sc_hd__and3_4 _17888_ (.A(_06758_),
    .B(_04223_),
    .C(_04212_),
    .X(_07500_));
 sky130_fd_sc_hd__nand2_8 _17889_ (.A(net272),
    .B(_04223_),
    .Y(_07501_));
 sky130_fd_sc_hd__nor4_4 _17890_ (.A(net262),
    .B(net244),
    .C(_05927_),
    .D(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__nand4_4 _17891_ (.A(_06519_),
    .B(_03955_),
    .C(_05926_),
    .D(_07500_),
    .Y(_07503_));
 sky130_fd_sc_hd__o31a_1 _17892_ (.A1(net233),
    .A2(_05927_),
    .A3(_07501_),
    .B1(_07499_),
    .X(_07504_));
 sky130_fd_sc_hd__o21ai_4 _17893_ (.A1(_05931_),
    .A2(_07501_),
    .B1(_07499_),
    .Y(_07506_));
 sky130_fd_sc_hd__a41oi_1 _17894_ (.A1(_11420_),
    .A2(net283),
    .A3(_05926_),
    .A4(_07500_),
    .B1(_03286_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand2_1 _17895_ (.A(_07499_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__o211ai_2 _17896_ (.A1(net175),
    .A2(_07074_),
    .B1(_04484_),
    .C1(_07072_),
    .Y(_07509_));
 sky130_fd_sc_hd__nor2_1 _17897_ (.A(_04212_),
    .B(_04331_),
    .Y(_07510_));
 sky130_fd_sc_hd__or3_2 _17898_ (.A(net44),
    .B(_04212_),
    .C(_03286_),
    .X(_07511_));
 sky130_fd_sc_hd__and4_1 _17899_ (.A(_07499_),
    .B(net167),
    .C(_07510_),
    .D(net33),
    .X(_07512_));
 sky130_fd_sc_hd__nand4_2 _17900_ (.A(_07499_),
    .B(net167),
    .C(_07510_),
    .D(net33),
    .Y(_07513_));
 sky130_fd_sc_hd__o311a_2 _17901_ (.A1(_03286_),
    .A2(net44),
    .A3(_04212_),
    .B1(_07508_),
    .C1(_07509_),
    .X(_07514_));
 sky130_fd_sc_hd__o211ai_4 _17902_ (.A1(_04212_),
    .A2(_04331_),
    .B1(_07508_),
    .C1(_07509_),
    .Y(_07515_));
 sky130_fd_sc_hd__a21oi_2 _17903_ (.A1(_07513_),
    .A2(_07515_),
    .B1(_07497_),
    .Y(_07517_));
 sky130_fd_sc_hd__o21bai_4 _17904_ (.A1(_07512_),
    .A2(_07514_),
    .B1_N(_07497_),
    .Y(_07518_));
 sky130_fd_sc_hd__nand2_2 _17905_ (.A(_07497_),
    .B(_07513_),
    .Y(_07519_));
 sky130_fd_sc_hd__o311a_2 _17906_ (.A1(_03286_),
    .A2(_07506_),
    .A3(_07511_),
    .B1(_07515_),
    .C1(_07497_),
    .X(_07520_));
 sky130_fd_sc_hd__nand3_1 _17907_ (.A(_07497_),
    .B(_07513_),
    .C(_07515_),
    .Y(_07521_));
 sky130_fd_sc_hd__a21oi_2 _17908_ (.A1(_07084_),
    .A2(_07087_),
    .B1(_07081_),
    .Y(_07522_));
 sky130_fd_sc_hd__a32o_2 _17909_ (.A1(net33),
    .A2(_07070_),
    .A3(_07077_),
    .B1(_07084_),
    .B2(_07087_),
    .X(_07523_));
 sky130_fd_sc_hd__a21oi_4 _17910_ (.A1(_07518_),
    .A2(_07521_),
    .B1(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__o21ai_2 _17911_ (.A1(_07517_),
    .A2(_07520_),
    .B1(_07522_),
    .Y(_07525_));
 sky130_fd_sc_hd__nor3_2 _17912_ (.A(_07517_),
    .B(_07520_),
    .C(_07522_),
    .Y(_07526_));
 sky130_fd_sc_hd__o211ai_4 _17913_ (.A1(_07519_),
    .A2(_07514_),
    .B1(_07518_),
    .C1(_07523_),
    .Y(_07528_));
 sky130_fd_sc_hd__o2111ai_4 _17914_ (.A1(_07492_),
    .A2(_07488_),
    .B1(_07491_),
    .C1(_07525_),
    .D1(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__o22ai_4 _17915_ (.A1(_07490_),
    .A2(_07493_),
    .B1(_07524_),
    .B2(_07526_),
    .Y(_07530_));
 sky130_fd_sc_hd__o211ai_4 _17916_ (.A1(_07490_),
    .A2(_07493_),
    .B1(_07525_),
    .C1(_07528_),
    .Y(_07531_));
 sky130_fd_sc_hd__o21bai_4 _17917_ (.A1(_07524_),
    .A2(_07526_),
    .B1_N(_07495_),
    .Y(_07532_));
 sky130_fd_sc_hd__a31oi_4 _17918_ (.A1(_07063_),
    .A2(_07066_),
    .A3(_07093_),
    .B1(_07094_),
    .Y(_07533_));
 sky130_fd_sc_hd__nand2_2 _17919_ (.A(_07095_),
    .B(_07098_),
    .Y(_07534_));
 sky130_fd_sc_hd__a21oi_1 _17920_ (.A1(_07529_),
    .A2(_07530_),
    .B1(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__nand3_2 _17921_ (.A(_07531_),
    .B(_07532_),
    .C(_07533_),
    .Y(_07536_));
 sky130_fd_sc_hd__nand3_4 _17922_ (.A(_07529_),
    .B(_07530_),
    .C(_07534_),
    .Y(_07537_));
 sky130_fd_sc_hd__a22o_1 _17923_ (.A1(_07479_),
    .A2(_07480_),
    .B1(_07536_),
    .B2(_07537_),
    .X(_07539_));
 sky130_fd_sc_hd__nand4_4 _17924_ (.A(_07479_),
    .B(_07480_),
    .C(_07536_),
    .D(_07537_),
    .Y(_07540_));
 sky130_fd_sc_hd__nand3_2 _17925_ (.A(_07481_),
    .B(_07536_),
    .C(_07537_),
    .Y(_07541_));
 sky130_fd_sc_hd__a21o_1 _17926_ (.A1(_07536_),
    .A2(_07537_),
    .B1(_07481_),
    .X(_07542_));
 sky130_fd_sc_hd__nand2_2 _17927_ (.A(_07539_),
    .B(_07540_),
    .Y(_07543_));
 sky130_fd_sc_hd__o21ai_2 _17928_ (.A1(_07101_),
    .A2(_07049_),
    .B1(_07104_),
    .Y(_07544_));
 sky130_fd_sc_hd__inv_2 _17929_ (.A(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__a2bb2oi_1 _17930_ (.A1_N(_07103_),
    .A2_N(_07106_),
    .B1(_07541_),
    .B2(_07542_),
    .Y(_07546_));
 sky130_fd_sc_hd__o211ai_4 _17931_ (.A1(_07103_),
    .A2(_07106_),
    .B1(_07539_),
    .C1(_07540_),
    .Y(_07547_));
 sky130_fd_sc_hd__a21oi_1 _17932_ (.A1(_07539_),
    .A2(_07540_),
    .B1(_07544_),
    .Y(_07548_));
 sky130_fd_sc_hd__o2111ai_4 _17933_ (.A1(_07049_),
    .A2(_07101_),
    .B1(_07104_),
    .C1(_07541_),
    .D1(_07542_),
    .Y(_07550_));
 sky130_fd_sc_hd__o21ai_4 _17934_ (.A1(_07457_),
    .A2(_07458_),
    .B1(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__o211ai_1 _17935_ (.A1(_07455_),
    .A2(_07456_),
    .B1(_07547_),
    .C1(_07550_),
    .Y(_07552_));
 sky130_fd_sc_hd__o22ai_1 _17936_ (.A1(_07457_),
    .A2(_07458_),
    .B1(_07546_),
    .B2(_07548_),
    .Y(_07553_));
 sky130_fd_sc_hd__o22ai_2 _17937_ (.A1(_07455_),
    .A2(_07456_),
    .B1(_07546_),
    .B2(_07548_),
    .Y(_07554_));
 sky130_fd_sc_hd__o211ai_2 _17938_ (.A1(_07457_),
    .A2(_07458_),
    .B1(_07547_),
    .C1(_07550_),
    .Y(_07555_));
 sky130_fd_sc_hd__a32oi_4 _17939_ (.A1(_07108_),
    .A2(_07110_),
    .A3(_07109_),
    .B1(_07169_),
    .B2(_07114_),
    .Y(_07556_));
 sky130_fd_sc_hd__a21boi_1 _17940_ (.A1(_07113_),
    .A2(_07168_),
    .B1_N(_07114_),
    .Y(_07557_));
 sky130_fd_sc_hd__nand3_2 _17941_ (.A(_07552_),
    .B(_07553_),
    .C(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__nand3_4 _17942_ (.A(_07554_),
    .B(_07556_),
    .C(_07555_),
    .Y(_07559_));
 sky130_fd_sc_hd__nand3_2 _17943_ (.A(_07412_),
    .B(_07558_),
    .C(_07559_),
    .Y(_07561_));
 sky130_fd_sc_hd__a21o_1 _17944_ (.A1(_07558_),
    .A2(_07559_),
    .B1(_07412_),
    .X(_07562_));
 sky130_fd_sc_hd__nand2_2 _17945_ (.A(_07558_),
    .B(_07411_),
    .Y(_07563_));
 sky130_fd_sc_hd__and3_1 _17946_ (.A(_07558_),
    .B(_07559_),
    .C(_07411_),
    .X(_07564_));
 sky130_fd_sc_hd__a21o_1 _17947_ (.A1(_07558_),
    .A2(_07559_),
    .B1(_07411_),
    .X(_07565_));
 sky130_fd_sc_hd__o21ai_2 _17948_ (.A1(_07174_),
    .A2(_07182_),
    .B1(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__a2bb2oi_4 _17949_ (.A1_N(_07174_),
    .A2_N(_07182_),
    .B1(_07561_),
    .B2(_07562_),
    .Y(_07567_));
 sky130_fd_sc_hd__o211a_1 _17950_ (.A1(_07177_),
    .A2(_07327_),
    .B1(_07561_),
    .C1(_07562_),
    .X(_07568_));
 sky130_fd_sc_hd__o2111ai_4 _17951_ (.A1(_07177_),
    .A2(_07024_),
    .B1(_07175_),
    .C1(_07561_),
    .D1(_07562_),
    .Y(_07569_));
 sky130_fd_sc_hd__o22ai_4 _17952_ (.A1(_07323_),
    .A2(_07325_),
    .B1(_07567_),
    .B2(_07568_),
    .Y(_07570_));
 sky130_fd_sc_hd__nand2_1 _17953_ (.A(_07569_),
    .B(_07326_),
    .Y(_07572_));
 sky130_fd_sc_hd__o211ai_1 _17954_ (.A1(_07564_),
    .A2(_07566_),
    .B1(_07569_),
    .C1(_07326_),
    .Y(_07573_));
 sky130_fd_sc_hd__o221ai_2 _17955_ (.A1(_07323_),
    .A2(_07325_),
    .B1(_07564_),
    .B2(_07566_),
    .C1(_07569_),
    .Y(_07574_));
 sky130_fd_sc_hd__o21ai_1 _17956_ (.A1(_07567_),
    .A2(_07568_),
    .B1(_07326_),
    .Y(_07575_));
 sky130_fd_sc_hd__o31a_1 _17957_ (.A1(_06852_),
    .A2(_06944_),
    .A3(_07184_),
    .B1(_07240_),
    .X(_07576_));
 sky130_fd_sc_hd__nand2_1 _17958_ (.A(_07188_),
    .B(_07240_),
    .Y(_07577_));
 sky130_fd_sc_hd__a21oi_1 _17959_ (.A1(_07570_),
    .A2(_07573_),
    .B1(_07577_),
    .Y(_07578_));
 sky130_fd_sc_hd__nand3_2 _17960_ (.A(_07576_),
    .B(_07575_),
    .C(_07574_),
    .Y(_07579_));
 sky130_fd_sc_hd__o221a_1 _17961_ (.A1(_07567_),
    .A2(_07572_),
    .B1(_07186_),
    .B2(_07239_),
    .C1(_07570_),
    .X(_07580_));
 sky130_fd_sc_hd__o221ai_4 _17962_ (.A1(_07567_),
    .A2(_07572_),
    .B1(_07186_),
    .B2(_07239_),
    .C1(_07570_),
    .Y(_07581_));
 sky130_fd_sc_hd__a21o_1 _17963_ (.A1(_06898_),
    .A2(_07233_),
    .B1(_07232_),
    .X(_07583_));
 sky130_fd_sc_hd__a21oi_1 _17964_ (.A1(_06898_),
    .A2(_07233_),
    .B1(_07232_),
    .Y(_07584_));
 sky130_fd_sc_hd__a21o_1 _17965_ (.A1(_07579_),
    .A2(_07581_),
    .B1(_07583_),
    .X(_07585_));
 sky130_fd_sc_hd__o211ai_1 _17966_ (.A1(_07232_),
    .A2(_07237_),
    .B1(_07579_),
    .C1(_07581_),
    .Y(_07586_));
 sky130_fd_sc_hd__o22ai_2 _17967_ (.A1(_07232_),
    .A2(_07237_),
    .B1(_07578_),
    .B2(_07580_),
    .Y(_07587_));
 sky130_fd_sc_hd__nand3_1 _17968_ (.A(_07579_),
    .B(_07581_),
    .C(_07584_),
    .Y(_07588_));
 sky130_fd_sc_hd__nand2_1 _17969_ (.A(_07585_),
    .B(_07586_),
    .Y(_07589_));
 sky130_fd_sc_hd__o211ai_1 _17970_ (.A1(_07245_),
    .A2(_07260_),
    .B1(_07587_),
    .C1(_07588_),
    .Y(_07590_));
 sky130_fd_sc_hd__a21boi_2 _17971_ (.A1(_07587_),
    .A2(_07588_),
    .B1_N(_07261_),
    .Y(_07591_));
 sky130_fd_sc_hd__nand3_1 _17972_ (.A(_07585_),
    .B(_07586_),
    .C(_07261_),
    .Y(_07592_));
 sky130_fd_sc_hd__o2bb2ai_1 _17973_ (.A1_N(_07590_),
    .A2_N(_07592_),
    .B1(_06939_),
    .B2(_07251_),
    .Y(_07594_));
 sky130_fd_sc_hd__nand2_1 _17974_ (.A(_07590_),
    .B(_07254_),
    .Y(_07595_));
 sky130_fd_sc_hd__o21ai_1 _17975_ (.A1(_07591_),
    .A2(_07595_),
    .B1(_07594_),
    .Y(_07596_));
 sky130_fd_sc_hd__o2bb2ai_1 _17976_ (.A1_N(_07255_),
    .A2_N(_07257_),
    .B1(_06933_),
    .B2(_07256_),
    .Y(_07597_));
 sky130_fd_sc_hd__a31o_1 _17977_ (.A1(_06934_),
    .A2(_06935_),
    .A3(_07258_),
    .B1(_07597_),
    .X(_07598_));
 sky130_fd_sc_hd__and4_2 _17978_ (.A(_06310_),
    .B(_06621_),
    .C(_06934_),
    .D(_07258_),
    .X(_07599_));
 sky130_fd_sc_hd__a21oi_1 _17979_ (.A1(_06320_),
    .A2(_07599_),
    .B1(_07598_),
    .Y(_07600_));
 sky130_fd_sc_hd__xor2_1 _17980_ (.A(_07596_),
    .B(_07600_),
    .X(net85));
 sky130_fd_sc_hd__o22ai_2 _17981_ (.A1(_07591_),
    .A2(_07595_),
    .B1(_07596_),
    .B2(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__a21o_1 _17982_ (.A1(_07324_),
    .A2(_07320_),
    .B1(_07317_),
    .X(_07602_));
 sky130_fd_sc_hd__inv_2 _17983_ (.A(_07602_),
    .Y(_07604_));
 sky130_fd_sc_hd__o31ai_2 _17984_ (.A1(_07004_),
    .A2(_07292_),
    .A3(_07293_),
    .B1(_07302_),
    .Y(_07605_));
 sky130_fd_sc_hd__a31oi_1 _17985_ (.A1(_07368_),
    .A2(_07369_),
    .A3(_07370_),
    .B1(_07391_),
    .Y(_07606_));
 sky130_fd_sc_hd__a31o_1 _17986_ (.A1(_07368_),
    .A2(_07369_),
    .A3(_07370_),
    .B1(_07391_),
    .X(_07607_));
 sky130_fd_sc_hd__a21o_1 _17987_ (.A1(_07265_),
    .A2(_07273_),
    .B1(_07271_),
    .X(_07608_));
 sky130_fd_sc_hd__a21oi_1 _17988_ (.A1(_07378_),
    .A2(_07381_),
    .B1(_07376_),
    .Y(_07609_));
 sky130_fd_sc_hd__a21o_1 _17989_ (.A1(_07376_),
    .A2(_07386_),
    .B1(_07382_),
    .X(_07610_));
 sky130_fd_sc_hd__o32a_1 _17990_ (.A1(_06864_),
    .A2(net306),
    .A3(_04703_),
    .B1(_03506_),
    .B2(_06866_),
    .X(_07611_));
 sky130_fd_sc_hd__a32o_1 _17991_ (.A1(_06863_),
    .A2(_04747_),
    .A3(net313),
    .B1(net26),
    .B2(_06865_),
    .X(_07612_));
 sky130_fd_sc_hd__or3b_2 _17992_ (.A(_03616_),
    .B(net50),
    .C_N(net49),
    .X(_07613_));
 sky130_fd_sc_hd__nand3_2 _17993_ (.A(net266),
    .B(net301),
    .C(_06324_),
    .Y(_07615_));
 sky130_fd_sc_hd__or3b_2 _17994_ (.A(_03725_),
    .B(net49),
    .C_N(net48),
    .X(_07616_));
 sky130_fd_sc_hd__o211ai_4 _17995_ (.A1(_04747_),
    .A2(_05436_),
    .B1(_06026_),
    .C1(_05414_),
    .Y(_07617_));
 sky130_fd_sc_hd__a22oi_4 _17996_ (.A1(_07613_),
    .A2(_07615_),
    .B1(_07616_),
    .B2(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__a22o_1 _17997_ (.A1(_07613_),
    .A2(_07615_),
    .B1(_07616_),
    .B2(_07617_),
    .X(_07619_));
 sky130_fd_sc_hd__nand4_2 _17998_ (.A(_07613_),
    .B(_07615_),
    .C(_07616_),
    .D(_07617_),
    .Y(_07620_));
 sky130_fd_sc_hd__a21oi_1 _17999_ (.A1(_07619_),
    .A2(_07620_),
    .B1(_07612_),
    .Y(_07621_));
 sky130_fd_sc_hd__a21o_1 _18000_ (.A1(_07619_),
    .A2(_07620_),
    .B1(_07612_),
    .X(_07622_));
 sky130_fd_sc_hd__nor3b_2 _18001_ (.A(_07611_),
    .B(_07618_),
    .C_N(_07620_),
    .Y(_07623_));
 sky130_fd_sc_hd__nand3_1 _18002_ (.A(_07612_),
    .B(_07619_),
    .C(_07620_),
    .Y(_07624_));
 sky130_fd_sc_hd__nand3_2 _18003_ (.A(_07610_),
    .B(_07622_),
    .C(_07624_),
    .Y(_07626_));
 sky130_fd_sc_hd__o22ai_4 _18004_ (.A1(_07385_),
    .A2(_07609_),
    .B1(_07621_),
    .B2(_07623_),
    .Y(_07627_));
 sky130_fd_sc_hd__a21oi_1 _18005_ (.A1(_07626_),
    .A2(_07627_),
    .B1(_07608_),
    .Y(_07628_));
 sky130_fd_sc_hd__a21o_1 _18006_ (.A1(_07626_),
    .A2(_07627_),
    .B1(_07608_),
    .X(_07629_));
 sky130_fd_sc_hd__o211a_1 _18007_ (.A1(_07271_),
    .A2(_07279_),
    .B1(_07626_),
    .C1(_07627_),
    .X(_07630_));
 sky130_fd_sc_hd__o211ai_2 _18008_ (.A1(_07271_),
    .A2(_07279_),
    .B1(_07626_),
    .C1(_07627_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand4_4 _18009_ (.A(_07372_),
    .B(_07607_),
    .C(_07629_),
    .D(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__o22ai_2 _18010_ (.A1(_07371_),
    .A2(_07606_),
    .B1(_07628_),
    .B2(_07630_),
    .Y(_07633_));
 sky130_fd_sc_hd__o21ai_1 _18011_ (.A1(_07204_),
    .A2(_07283_),
    .B1(_07286_),
    .Y(_07634_));
 sky130_fd_sc_hd__nand3_2 _18012_ (.A(_07632_),
    .B(_07633_),
    .C(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__a21o_1 _18013_ (.A1(_07632_),
    .A2(_07633_),
    .B1(_07634_),
    .X(_07637_));
 sky130_fd_sc_hd__a21oi_1 _18014_ (.A1(_07635_),
    .A2(_07637_),
    .B1(_07605_),
    .Y(_07638_));
 sky130_fd_sc_hd__a21o_1 _18015_ (.A1(_07635_),
    .A2(_07637_),
    .B1(_07605_),
    .X(_07639_));
 sky130_fd_sc_hd__and3_1 _18016_ (.A(_07605_),
    .B(_07635_),
    .C(_07637_),
    .X(_07640_));
 sky130_fd_sc_hd__nand3_1 _18017_ (.A(_07605_),
    .B(_07635_),
    .C(_07637_),
    .Y(_07641_));
 sky130_fd_sc_hd__and2_4 _18018_ (.A(_04234_),
    .B(net54),
    .X(_07642_));
 sky130_fd_sc_hd__nor2_8 _18019_ (.A(net54),
    .B(_04234_),
    .Y(_07643_));
 sky130_fd_sc_hd__o21ai_1 _18020_ (.A1(_07642_),
    .A2(_07643_),
    .B1(net1),
    .Y(_07644_));
 sky130_fd_sc_hd__a22o_1 _18021_ (.A1(_04539_),
    .A2(_07305_),
    .B1(_07308_),
    .B2(net12),
    .X(_07645_));
 sky130_fd_sc_hd__a32o_1 _18022_ (.A1(net318),
    .A2(_04452_),
    .A3(_07223_),
    .B1(_07225_),
    .B2(net23),
    .X(_07646_));
 sky130_fd_sc_hd__nand2_1 _18023_ (.A(_07645_),
    .B(_07646_),
    .Y(_07648_));
 sky130_fd_sc_hd__nor2_1 _18024_ (.A(_07645_),
    .B(_07646_),
    .Y(_07649_));
 sky130_fd_sc_hd__a221o_1 _18025_ (.A1(_04539_),
    .A2(_07305_),
    .B1(_07308_),
    .B2(net12),
    .C1(_07646_),
    .X(_07650_));
 sky130_fd_sc_hd__a21boi_1 _18026_ (.A1(_07648_),
    .A2(_07650_),
    .B1_N(_07644_),
    .Y(_07651_));
 sky130_fd_sc_hd__o2111a_1 _18027_ (.A1(_07642_),
    .A2(_07643_),
    .B1(net1),
    .C1(_07648_),
    .D1(_07650_),
    .X(_07652_));
 sky130_fd_sc_hd__nor2_2 _18028_ (.A(_07651_),
    .B(_07652_),
    .Y(_07653_));
 sky130_fd_sc_hd__nand2_2 _18029_ (.A(_07311_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__a21o_1 _18030_ (.A1(_07309_),
    .A2(_07310_),
    .B1(_07653_),
    .X(_07655_));
 sky130_fd_sc_hd__nand2_1 _18031_ (.A(_07654_),
    .B(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__o21ai_2 _18032_ (.A1(_07638_),
    .A2(_07640_),
    .B1(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__nor2_1 _18033_ (.A(_07656_),
    .B(_07638_),
    .Y(_07659_));
 sky130_fd_sc_hd__nand3b_2 _18034_ (.A_N(_07656_),
    .B(_07641_),
    .C(_07639_),
    .Y(_07660_));
 sky130_fd_sc_hd__nand2_1 _18035_ (.A(_07657_),
    .B(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__a31o_1 _18036_ (.A1(_07400_),
    .A2(_07402_),
    .A3(_07403_),
    .B1(_07409_),
    .X(_07662_));
 sky130_fd_sc_hd__nand3_2 _18037_ (.A(_07407_),
    .B(_07410_),
    .C(_07661_),
    .Y(_07663_));
 sky130_fd_sc_hd__inv_2 _18038_ (.A(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__and3_1 _18039_ (.A(_07657_),
    .B(_07660_),
    .C(_07662_),
    .X(_07665_));
 sky130_fd_sc_hd__a21o_2 _18040_ (.A1(_07407_),
    .A2(_07410_),
    .B1(_07661_),
    .X(_07666_));
 sky130_fd_sc_hd__nand2_1 _18041_ (.A(_07304_),
    .B(_07315_),
    .Y(_07667_));
 sky130_fd_sc_hd__inv_2 _18042_ (.A(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__a21oi_1 _18043_ (.A1(_07663_),
    .A2(_07666_),
    .B1(_07667_),
    .Y(_07670_));
 sky130_fd_sc_hd__a21o_2 _18044_ (.A1(_07663_),
    .A2(_07666_),
    .B1(_07667_),
    .X(_07671_));
 sky130_fd_sc_hd__a31o_2 _18045_ (.A1(_07407_),
    .A2(_07410_),
    .A3(_07661_),
    .B1(_07668_),
    .X(_07672_));
 sky130_fd_sc_hd__and3_1 _18046_ (.A(_07663_),
    .B(_07666_),
    .C(_07667_),
    .X(_07673_));
 sky130_fd_sc_hd__a31o_1 _18047_ (.A1(_07657_),
    .A2(_07660_),
    .A3(_07662_),
    .B1(_07672_),
    .X(_07674_));
 sky130_fd_sc_hd__a21oi_1 _18048_ (.A1(_07663_),
    .A2(_07666_),
    .B1(_07668_),
    .Y(_07675_));
 sky130_fd_sc_hd__and3_1 _18049_ (.A(_07663_),
    .B(_07666_),
    .C(_07668_),
    .X(_07676_));
 sky130_fd_sc_hd__o21ai_1 _18050_ (.A1(_07665_),
    .A2(_07672_),
    .B1(_07671_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand2_2 _18051_ (.A(_07559_),
    .B(_07563_),
    .Y(_07678_));
 sky130_fd_sc_hd__nand2_1 _18052_ (.A(_07453_),
    .B(_07454_),
    .Y(_07679_));
 sky130_fd_sc_hd__a21o_1 _18053_ (.A1(_07358_),
    .A2(_07365_),
    .B1(_07366_),
    .X(_07681_));
 sky130_fd_sc_hd__a32o_1 _18054_ (.A1(net256),
    .A2(_08700_),
    .A3(_04985_),
    .B1(_04988_),
    .B2(net32),
    .X(_07682_));
 sky130_fd_sc_hd__o211ai_4 _18055_ (.A1(net260),
    .A2(_09665_),
    .B1(net243),
    .C1(_09698_),
    .Y(_07683_));
 sky130_fd_sc_hd__or3b_1 _18056_ (.A(_03960_),
    .B(net43),
    .C_N(net42),
    .X(_07684_));
 sky130_fd_sc_hd__nor2_1 _18057_ (.A(_03982_),
    .B(_04483_),
    .Y(_07685_));
 sky130_fd_sc_hd__or3b_2 _18058_ (.A(_03982_),
    .B(net42),
    .C_N(net41),
    .X(_07686_));
 sky130_fd_sc_hd__o311a_1 _18059_ (.A1(_04747_),
    .A2(net264),
    .A3(_11387_),
    .B1(net279),
    .C1(_11354_),
    .X(_07687_));
 sky130_fd_sc_hd__nand2_1 _18060_ (.A(_11442_),
    .B(net279),
    .Y(_07688_));
 sky130_fd_sc_hd__a22oi_1 _18061_ (.A1(_07683_),
    .A2(_07684_),
    .B1(_07686_),
    .B2(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__o2bb2ai_2 _18062_ (.A1_N(_07683_),
    .A2_N(_07684_),
    .B1(_07685_),
    .B2(_07687_),
    .Y(_07690_));
 sky130_fd_sc_hd__o2111ai_4 _18063_ (.A1(_03960_),
    .A2(_04898_),
    .B1(_07683_),
    .C1(_07686_),
    .D1(_07688_),
    .Y(_07692_));
 sky130_fd_sc_hd__a21oi_1 _18064_ (.A1(_07690_),
    .A2(_07692_),
    .B1(_07682_),
    .Y(_07693_));
 sky130_fd_sc_hd__a21o_1 _18065_ (.A1(_07690_),
    .A2(_07692_),
    .B1(_07682_),
    .X(_07694_));
 sky130_fd_sc_hd__and3_1 _18066_ (.A(_07682_),
    .B(_07690_),
    .C(_07692_),
    .X(_07695_));
 sky130_fd_sc_hd__nand3_1 _18067_ (.A(_07682_),
    .B(_07690_),
    .C(_07692_),
    .Y(_07696_));
 sky130_fd_sc_hd__a21oi_1 _18068_ (.A1(_07694_),
    .A2(_07696_),
    .B1(_07681_),
    .Y(_07697_));
 sky130_fd_sc_hd__o21bai_1 _18069_ (.A1(_07693_),
    .A2(_07695_),
    .B1_N(_07681_),
    .Y(_07698_));
 sky130_fd_sc_hd__nand3_2 _18070_ (.A(_07681_),
    .B(_07694_),
    .C(_07696_),
    .Y(_07699_));
 sky130_fd_sc_hd__o2bb2a_1 _18071_ (.A1_N(_05874_),
    .A2_N(net275),
    .B1(_05766_),
    .B2(_03835_),
    .X(_07700_));
 sky130_fd_sc_hd__a32oi_4 _18072_ (.A1(_06486_),
    .A2(net260),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net30),
    .Y(_07701_));
 sky130_fd_sc_hd__or3_1 _18073_ (.A(net46),
    .B(_04124_),
    .C(_03938_),
    .X(_07703_));
 sky130_fd_sc_hd__nand3_1 _18074_ (.A(_07242_),
    .B(net257),
    .C(net276),
    .Y(_07704_));
 sky130_fd_sc_hd__a21o_1 _18075_ (.A1(_07703_),
    .A2(_07704_),
    .B1(_07701_),
    .X(_07705_));
 sky130_fd_sc_hd__o221ai_4 _18076_ (.A1(_07263_),
    .A2(_05226_),
    .B1(_05229_),
    .B2(_03938_),
    .C1(_07701_),
    .Y(_07706_));
 sky130_fd_sc_hd__a21o_1 _18077_ (.A1(_07705_),
    .A2(_07706_),
    .B1(_07700_),
    .X(_07707_));
 sky130_fd_sc_hd__nand3_1 _18078_ (.A(_07705_),
    .B(_07706_),
    .C(_07700_),
    .Y(_07708_));
 sky130_fd_sc_hd__nand2_1 _18079_ (.A(_07707_),
    .B(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__a21oi_1 _18080_ (.A1(_07698_),
    .A2(_07699_),
    .B1(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__a21oi_1 _18081_ (.A1(_07707_),
    .A2(_07708_),
    .B1(_07697_),
    .Y(_07711_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(_07698_),
    .B(_07709_),
    .Y(_07712_));
 sky130_fd_sc_hd__a21oi_2 _18083_ (.A1(_07711_),
    .A2(_07699_),
    .B1(_07710_),
    .Y(_07714_));
 sky130_fd_sc_hd__o22a_1 _18084_ (.A1(_07349_),
    .A2(_07344_),
    .B1(_07330_),
    .B2(_07347_),
    .X(_07715_));
 sky130_fd_sc_hd__o22ai_1 _18085_ (.A1(_07349_),
    .A2(_07344_),
    .B1(_07330_),
    .B2(_07347_),
    .Y(_07716_));
 sky130_fd_sc_hd__o21ai_2 _18086_ (.A1(_07334_),
    .A2(_07337_),
    .B1(_07345_),
    .Y(_07717_));
 sky130_fd_sc_hd__o21a_1 _18087_ (.A1(_07435_),
    .A2(_07438_),
    .B1(_07432_),
    .X(_07718_));
 sky130_fd_sc_hd__a21oi_1 _18088_ (.A1(_07432_),
    .A2(_07442_),
    .B1(_07440_),
    .Y(_07719_));
 sky130_fd_sc_hd__o22a_1 _18089_ (.A1(_13021_),
    .A2(_04268_),
    .B1(_04270_),
    .B2(_04004_),
    .X(_07720_));
 sky130_fd_sc_hd__a32o_1 _18090_ (.A1(net234),
    .A2(net251),
    .A3(net280),
    .B1(_04269_),
    .B2(net4),
    .X(_07721_));
 sky130_fd_sc_hd__o211ai_4 _18091_ (.A1(net254),
    .A2(_02442_),
    .B1(net285),
    .C1(_02421_),
    .Y(_07722_));
 sky130_fd_sc_hd__or3_2 _18092_ (.A(net39),
    .B(_04037_),
    .C(_04026_),
    .X(_07723_));
 sky130_fd_sc_hd__or3b_4 _18093_ (.A(_04015_),
    .B(net40),
    .C_N(net39),
    .X(_07725_));
 sky130_fd_sc_hd__o211ai_4 _18094_ (.A1(net254),
    .A2(_00646_),
    .B1(net281),
    .C1(_00625_),
    .Y(_07726_));
 sky130_fd_sc_hd__a22oi_4 _18095_ (.A1(_07722_),
    .A2(_07723_),
    .B1(_07725_),
    .B2(_07726_),
    .Y(_07727_));
 sky130_fd_sc_hd__a22o_1 _18096_ (.A1(_07722_),
    .A2(_07723_),
    .B1(_07725_),
    .B2(_07726_),
    .X(_07728_));
 sky130_fd_sc_hd__o2111a_1 _18097_ (.A1(_04026_),
    .A2(_03737_),
    .B1(_07722_),
    .C1(_07725_),
    .D1(_07726_),
    .X(_07729_));
 sky130_fd_sc_hd__o2111ai_4 _18098_ (.A1(_04026_),
    .A2(_03737_),
    .B1(_07722_),
    .C1(_07725_),
    .D1(_07726_),
    .Y(_07730_));
 sky130_fd_sc_hd__o21ai_1 _18099_ (.A1(_07727_),
    .A2(_07729_),
    .B1(_07721_),
    .Y(_07731_));
 sky130_fd_sc_hd__nand3_1 _18100_ (.A(_07720_),
    .B(_07728_),
    .C(_07730_),
    .Y(_07732_));
 sky130_fd_sc_hd__nor2_1 _18101_ (.A(_07720_),
    .B(_07729_),
    .Y(_07733_));
 sky130_fd_sc_hd__a21oi_1 _18102_ (.A1(_07721_),
    .A2(_07730_),
    .B1(_07727_),
    .Y(_07734_));
 sky130_fd_sc_hd__o21ai_1 _18103_ (.A1(_07727_),
    .A2(_07729_),
    .B1(_07720_),
    .Y(_07736_));
 sky130_fd_sc_hd__and3_1 _18104_ (.A(_07721_),
    .B(_07728_),
    .C(_07730_),
    .X(_07737_));
 sky130_fd_sc_hd__nand3_1 _18105_ (.A(_07721_),
    .B(_07728_),
    .C(_07730_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand3_2 _18106_ (.A(_07719_),
    .B(_07731_),
    .C(_07732_),
    .Y(_07739_));
 sky130_fd_sc_hd__o21ai_1 _18107_ (.A1(_07440_),
    .A2(_07718_),
    .B1(_07736_),
    .Y(_07740_));
 sky130_fd_sc_hd__o211a_1 _18108_ (.A1(_07440_),
    .A2(_07718_),
    .B1(_07736_),
    .C1(_07738_),
    .X(_07741_));
 sky130_fd_sc_hd__o211ai_2 _18109_ (.A1(_07440_),
    .A2(_07718_),
    .B1(_07736_),
    .C1(_07738_),
    .Y(_07742_));
 sky130_fd_sc_hd__a21o_1 _18110_ (.A1(_07739_),
    .A2(_07742_),
    .B1(_07717_),
    .X(_07743_));
 sky130_fd_sc_hd__nand2_1 _18111_ (.A(_07717_),
    .B(_07739_),
    .Y(_07744_));
 sky130_fd_sc_hd__o2111ai_1 _18112_ (.A1(_07334_),
    .A2(_07337_),
    .B1(_07345_),
    .C1(_07739_),
    .D1(_07742_),
    .Y(_07745_));
 sky130_fd_sc_hd__a22o_1 _18113_ (.A1(_07339_),
    .A2(_07345_),
    .B1(_07739_),
    .B2(_07742_),
    .X(_07747_));
 sky130_fd_sc_hd__nand3_2 _18114_ (.A(_07715_),
    .B(_07745_),
    .C(_07747_),
    .Y(_07748_));
 sky130_fd_sc_hd__o211ai_2 _18115_ (.A1(_07744_),
    .A2(_07741_),
    .B1(_07716_),
    .C1(_07743_),
    .Y(_07749_));
 sky130_fd_sc_hd__a21oi_1 _18116_ (.A1(_07748_),
    .A2(_07749_),
    .B1(_07714_),
    .Y(_07750_));
 sky130_fd_sc_hd__a21o_1 _18117_ (.A1(_07748_),
    .A2(_07749_),
    .B1(_07714_),
    .X(_07751_));
 sky130_fd_sc_hd__and3_1 _18118_ (.A(_07748_),
    .B(_07749_),
    .C(_07714_),
    .X(_07752_));
 sky130_fd_sc_hd__nand3_1 _18119_ (.A(_07748_),
    .B(_07749_),
    .C(_07714_),
    .Y(_07753_));
 sky130_fd_sc_hd__o2bb2ai_1 _18120_ (.A1_N(_07452_),
    .A2_N(_07679_),
    .B1(_07750_),
    .B2(_07752_),
    .Y(_07754_));
 sky130_fd_sc_hd__nand3_1 _18121_ (.A(_07452_),
    .B(_07679_),
    .C(_07751_),
    .Y(_07755_));
 sky130_fd_sc_hd__nand4_1 _18122_ (.A(_07452_),
    .B(_07679_),
    .C(_07751_),
    .D(_07753_),
    .Y(_07756_));
 sky130_fd_sc_hd__a21bo_1 _18123_ (.A1(_07397_),
    .A2(_07355_),
    .B1_N(_07356_),
    .X(_07758_));
 sky130_fd_sc_hd__a21oi_2 _18124_ (.A1(_07754_),
    .A2(_07756_),
    .B1(_07758_),
    .Y(_07759_));
 sky130_fd_sc_hd__o221a_2 _18125_ (.A1(_07357_),
    .A2(_07401_),
    .B1(_07752_),
    .B2(_07755_),
    .C1(_07754_),
    .X(_07760_));
 sky130_fd_sc_hd__nor2_2 _18126_ (.A(_07759_),
    .B(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__a21oi_2 _18127_ (.A1(_07497_),
    .A2(_07515_),
    .B1(_07512_),
    .Y(_07762_));
 sky130_fd_sc_hd__o32ai_4 _18128_ (.A1(_03286_),
    .A2(_07506_),
    .A3(_07511_),
    .B1(_07519_),
    .B2(_07514_),
    .Y(_07763_));
 sky130_fd_sc_hd__nor2_4 _18129_ (.A(net21),
    .B(net22),
    .Y(_07764_));
 sky130_fd_sc_hd__or2_4 _18130_ (.A(net21),
    .B(net22),
    .X(_07765_));
 sky130_fd_sc_hd__and3_4 _18131_ (.A(_06758_),
    .B(_07764_),
    .C(_04212_),
    .X(_07766_));
 sky130_fd_sc_hd__nand2_8 _18132_ (.A(net270),
    .B(_07764_),
    .Y(_07767_));
 sky130_fd_sc_hd__nand4_4 _18133_ (.A(_03957_),
    .B(_05926_),
    .C(net270),
    .D(_07764_),
    .Y(_07769_));
 sky130_fd_sc_hd__a41oi_2 _18134_ (.A1(_11420_),
    .A2(net284),
    .A3(_05926_),
    .A4(_07500_),
    .B1(_04245_),
    .Y(_07770_));
 sky130_fd_sc_hd__nand2_8 _18135_ (.A(_07503_),
    .B(net22),
    .Y(_07771_));
 sky130_fd_sc_hd__a31o_1 _18136_ (.A1(net204),
    .A2(net270),
    .A3(_07764_),
    .B1(_07770_),
    .X(_07772_));
 sky130_fd_sc_hd__o211ai_2 _18137_ (.A1(_07076_),
    .A2(_07765_),
    .B1(net33),
    .C1(_07771_),
    .Y(_07773_));
 sky130_fd_sc_hd__o211ai_2 _18138_ (.A1(net175),
    .A2(_07501_),
    .B1(_04484_),
    .C1(_07499_),
    .Y(_07774_));
 sky130_fd_sc_hd__o211ai_4 _18139_ (.A1(_04223_),
    .A2(_04331_),
    .B1(_07773_),
    .C1(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__inv_2 _18140_ (.A(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__and3_2 _18141_ (.A(net21),
    .B(_04320_),
    .C(_04245_),
    .X(_07777_));
 sky130_fd_sc_hd__or4_4 _18142_ (.A(net44),
    .B(net22),
    .C(_04223_),
    .D(_03286_),
    .X(_07778_));
 sky130_fd_sc_hd__nor2_1 _18143_ (.A(_04212_),
    .B(_04375_),
    .Y(_07780_));
 sky130_fd_sc_hd__o311a_1 _18144_ (.A1(net245),
    .A2(net241),
    .A3(_07074_),
    .B1(_04342_),
    .C1(_07072_),
    .X(_07781_));
 sky130_fd_sc_hd__a31o_1 _18145_ (.A1(_07072_),
    .A2(net168),
    .A3(_04342_),
    .B1(_07780_),
    .X(_07782_));
 sky130_fd_sc_hd__a21o_1 _18146_ (.A1(_07775_),
    .A2(_07778_),
    .B1(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__o21a_1 _18147_ (.A1(_07780_),
    .A2(_07781_),
    .B1(_07775_),
    .X(_07784_));
 sky130_fd_sc_hd__o21ai_2 _18148_ (.A1(_07780_),
    .A2(_07781_),
    .B1(_07775_),
    .Y(_07785_));
 sky130_fd_sc_hd__nand3b_2 _18149_ (.A_N(_07782_),
    .B(_07778_),
    .C(_07775_),
    .Y(_07786_));
 sky130_fd_sc_hd__o2bb2ai_2 _18150_ (.A1_N(_07775_),
    .A2_N(_07778_),
    .B1(_07780_),
    .B2(_07781_),
    .Y(_07787_));
 sky130_fd_sc_hd__nand2_1 _18151_ (.A(_07786_),
    .B(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__and3_1 _18152_ (.A(_07787_),
    .B(_07762_),
    .C(_07786_),
    .X(_07789_));
 sky130_fd_sc_hd__nand3_4 _18153_ (.A(_07787_),
    .B(_07762_),
    .C(_07786_),
    .Y(_07791_));
 sky130_fd_sc_hd__o211ai_4 _18154_ (.A1(_07785_),
    .A2(_07777_),
    .B1(_07763_),
    .C1(_07783_),
    .Y(_07792_));
 sky130_fd_sc_hd__a32o_1 _18155_ (.A1(_06219_),
    .A2(_06221_),
    .A3(_05227_),
    .B1(_05249_),
    .B2(net17),
    .X(_07793_));
 sky130_fd_sc_hd__or3b_2 _18156_ (.A(net58),
    .B(_04201_),
    .C_N(net55),
    .X(_07794_));
 sky130_fd_sc_hd__o211ai_4 _18157_ (.A1(net175),
    .A2(_06759_),
    .B1(_04627_),
    .C1(net196),
    .Y(_07795_));
 sky130_fd_sc_hd__o211ai_2 _18158_ (.A1(net175),
    .A2(_06451_),
    .B1(_04889_),
    .C1(net200),
    .Y(_07796_));
 sky130_fd_sc_hd__and3b_1 _18159_ (.A_N(net59),
    .B(net18),
    .C(net58),
    .X(_07797_));
 sky130_fd_sc_hd__or3b_1 _18160_ (.A(net59),
    .B(_04179_),
    .C_N(net58),
    .X(_07798_));
 sky130_fd_sc_hd__a31oi_2 _18161_ (.A1(net200),
    .A2(net172),
    .A3(_04889_),
    .B1(_07797_),
    .Y(_07799_));
 sky130_fd_sc_hd__o211a_2 _18162_ (.A1(_04201_),
    .A2(net316),
    .B1(_07795_),
    .C1(_07799_),
    .X(_07800_));
 sky130_fd_sc_hd__nand4_2 _18163_ (.A(_07794_),
    .B(_07795_),
    .C(_07796_),
    .D(_07798_),
    .Y(_07802_));
 sky130_fd_sc_hd__a21oi_2 _18164_ (.A1(_07794_),
    .A2(_07795_),
    .B1(_07799_),
    .Y(_07803_));
 sky130_fd_sc_hd__a22o_1 _18165_ (.A1(_07794_),
    .A2(_07795_),
    .B1(_07796_),
    .B2(_07798_),
    .X(_07804_));
 sky130_fd_sc_hd__nor2_1 _18166_ (.A(_07793_),
    .B(_07803_),
    .Y(_07805_));
 sky130_fd_sc_hd__a21o_1 _18167_ (.A1(_07793_),
    .A2(_07802_),
    .B1(_07803_),
    .X(_07806_));
 sky130_fd_sc_hd__a21oi_1 _18168_ (.A1(_07802_),
    .A2(_07804_),
    .B1(_07793_),
    .Y(_07807_));
 sky130_fd_sc_hd__o21bai_4 _18169_ (.A1(_07800_),
    .A2(_07803_),
    .B1_N(_07793_),
    .Y(_07808_));
 sky130_fd_sc_hd__and3_1 _18170_ (.A(_07793_),
    .B(_07802_),
    .C(_07804_),
    .X(_07809_));
 sky130_fd_sc_hd__nand3_2 _18171_ (.A(_07793_),
    .B(_07802_),
    .C(_07804_),
    .Y(_07810_));
 sky130_fd_sc_hd__o2bb2ai_4 _18172_ (.A1_N(_07791_),
    .A2_N(_07792_),
    .B1(_07807_),
    .B2(_07809_),
    .Y(_07811_));
 sky130_fd_sc_hd__nand3_2 _18173_ (.A(_07791_),
    .B(_07808_),
    .C(_07810_),
    .Y(_07813_));
 sky130_fd_sc_hd__nand4_4 _18174_ (.A(_07791_),
    .B(_07792_),
    .C(_07808_),
    .D(_07810_),
    .Y(_07814_));
 sky130_fd_sc_hd__o32a_1 _18175_ (.A1(_07517_),
    .A2(_07520_),
    .A3(_07522_),
    .B1(_07493_),
    .B2(_07490_),
    .X(_07815_));
 sky130_fd_sc_hd__o21ai_4 _18176_ (.A1(_07495_),
    .A2(_07524_),
    .B1(_07528_),
    .Y(_07816_));
 sky130_fd_sc_hd__a21oi_2 _18177_ (.A1(_07811_),
    .A2(_07814_),
    .B1(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__o2bb2ai_4 _18178_ (.A1_N(_07811_),
    .A2_N(_07814_),
    .B1(_07815_),
    .B2(_07524_),
    .Y(_07818_));
 sky130_fd_sc_hd__and3_1 _18179_ (.A(_07816_),
    .B(_07814_),
    .C(_07811_),
    .X(_07819_));
 sky130_fd_sc_hd__nand3_4 _18180_ (.A(_07816_),
    .B(_07814_),
    .C(_07811_),
    .Y(_07820_));
 sky130_fd_sc_hd__a21o_1 _18181_ (.A1(_07469_),
    .A2(_07470_),
    .B1(_07466_),
    .X(_07821_));
 sky130_fd_sc_hd__a21oi_4 _18182_ (.A1(_07482_),
    .A2(_07489_),
    .B1(_07487_),
    .Y(_07822_));
 sky130_fd_sc_hd__o22a_2 _18183_ (.A1(_04135_),
    .A2(_07691_),
    .B1(_05294_),
    .B2(_07669_),
    .X(_07824_));
 sky130_fd_sc_hd__a32o_1 _18184_ (.A1(net181),
    .A2(net180),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net14),
    .X(_07825_));
 sky130_fd_sc_hd__a221oi_2 _18185_ (.A1(_03957_),
    .A2(_05926_),
    .B1(net177),
    .B2(net16),
    .C1(_05699_),
    .Y(_07826_));
 sky130_fd_sc_hd__nor2_1 _18186_ (.A(_04157_),
    .B(_05720_),
    .Y(_07827_));
 sky130_fd_sc_hd__and3_1 _18187_ (.A(_03927_),
    .B(net15),
    .C(net61),
    .X(_07828_));
 sky130_fd_sc_hd__a31oi_4 _18188_ (.A1(_05549_),
    .A2(net177),
    .A3(net292),
    .B1(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__a31o_1 _18189_ (.A1(_05549_),
    .A2(net177),
    .A3(net292),
    .B1(_07828_),
    .X(_07830_));
 sky130_fd_sc_hd__o21ai_4 _18190_ (.A1(_07826_),
    .A2(_07827_),
    .B1(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__o221a_4 _18191_ (.A1(_04157_),
    .A2(_05720_),
    .B1(net155),
    .B2(_05699_),
    .C1(_07829_),
    .X(_07832_));
 sky130_fd_sc_hd__o221ai_4 _18192_ (.A1(_04157_),
    .A2(_05720_),
    .B1(net155),
    .B2(_05699_),
    .C1(_07829_),
    .Y(_07833_));
 sky130_fd_sc_hd__nand2_1 _18193_ (.A(_07831_),
    .B(_07833_),
    .Y(_07835_));
 sky130_fd_sc_hd__a21o_1 _18194_ (.A1(_07831_),
    .A2(_07833_),
    .B1(_07825_),
    .X(_07836_));
 sky130_fd_sc_hd__nand2_1 _18195_ (.A(_07825_),
    .B(_07831_),
    .Y(_07837_));
 sky130_fd_sc_hd__nand3_2 _18196_ (.A(_07825_),
    .B(_07831_),
    .C(_07833_),
    .Y(_07838_));
 sky130_fd_sc_hd__nand3_2 _18197_ (.A(_07831_),
    .B(_07833_),
    .C(_07824_),
    .Y(_07839_));
 sky130_fd_sc_hd__a21o_1 _18198_ (.A1(_07831_),
    .A2(_07833_),
    .B1(_07824_),
    .X(_07840_));
 sky130_fd_sc_hd__nand3_4 _18199_ (.A(_07840_),
    .B(_07822_),
    .C(_07839_),
    .Y(_07841_));
 sky130_fd_sc_hd__a21oi_2 _18200_ (.A1(_07835_),
    .A2(_07824_),
    .B1(_07822_),
    .Y(_07842_));
 sky130_fd_sc_hd__o221a_2 _18201_ (.A1(_07832_),
    .A2(_07837_),
    .B1(_07487_),
    .B2(_07493_),
    .C1(_07836_),
    .X(_07843_));
 sky130_fd_sc_hd__o221ai_4 _18202_ (.A1(_07832_),
    .A2(_07837_),
    .B1(_07487_),
    .B2(_07493_),
    .C1(_07836_),
    .Y(_07844_));
 sky130_fd_sc_hd__a22oi_1 _18203_ (.A1(_07467_),
    .A2(_07474_),
    .B1(_07841_),
    .B2(_07844_),
    .Y(_07846_));
 sky130_fd_sc_hd__a22o_1 _18204_ (.A1(_07467_),
    .A2(_07474_),
    .B1(_07841_),
    .B2(_07844_),
    .X(_07847_));
 sky130_fd_sc_hd__and4_1 _18205_ (.A(_07467_),
    .B(_07474_),
    .C(_07841_),
    .D(_07844_),
    .X(_07848_));
 sky130_fd_sc_hd__o2111ai_4 _18206_ (.A1(_07468_),
    .A2(_07473_),
    .B1(_07841_),
    .C1(_07844_),
    .D1(_07467_),
    .Y(_07849_));
 sky130_fd_sc_hd__a21oi_1 _18207_ (.A1(_07841_),
    .A2(_07844_),
    .B1(_07821_),
    .Y(_07850_));
 sky130_fd_sc_hd__a21o_1 _18208_ (.A1(_07841_),
    .A2(_07844_),
    .B1(_07821_),
    .X(_07851_));
 sky130_fd_sc_hd__a32oi_4 _18209_ (.A1(_07840_),
    .A2(_07822_),
    .A3(_07839_),
    .B1(_07474_),
    .B2(_07467_),
    .Y(_07852_));
 sky130_fd_sc_hd__and3_1 _18210_ (.A(_07821_),
    .B(_07841_),
    .C(_07844_),
    .X(_07853_));
 sky130_fd_sc_hd__nand2_1 _18211_ (.A(_07852_),
    .B(_07844_),
    .Y(_07854_));
 sky130_fd_sc_hd__o2bb2ai_1 _18212_ (.A1_N(_07818_),
    .A2_N(_07820_),
    .B1(_07850_),
    .B2(_07853_),
    .Y(_07855_));
 sky130_fd_sc_hd__nand3_2 _18213_ (.A(_07818_),
    .B(_07851_),
    .C(_07854_),
    .Y(_07857_));
 sky130_fd_sc_hd__o2bb2ai_1 _18214_ (.A1_N(_07818_),
    .A2_N(_07820_),
    .B1(_07846_),
    .B2(_07848_),
    .Y(_07858_));
 sky130_fd_sc_hd__nand4_2 _18215_ (.A(_07818_),
    .B(_07820_),
    .C(_07847_),
    .D(_07849_),
    .Y(_07859_));
 sky130_fd_sc_hd__a32oi_4 _18216_ (.A1(_07529_),
    .A2(_07530_),
    .A3(_07534_),
    .B1(_07480_),
    .B2(_07479_),
    .Y(_07860_));
 sky130_fd_sc_hd__a32oi_4 _18217_ (.A1(_07531_),
    .A2(_07533_),
    .A3(_07532_),
    .B1(_07481_),
    .B2(_07537_),
    .Y(_07861_));
 sky130_fd_sc_hd__o211ai_4 _18218_ (.A1(_07535_),
    .A2(_07860_),
    .B1(_07859_),
    .C1(_07858_),
    .Y(_07862_));
 sky130_fd_sc_hd__inv_2 _18219_ (.A(_07862_),
    .Y(_07863_));
 sky130_fd_sc_hd__o211ai_4 _18220_ (.A1(_07819_),
    .A2(_07857_),
    .B1(_07855_),
    .C1(_07861_),
    .Y(_07864_));
 sky130_fd_sc_hd__o21ai_2 _18221_ (.A1(_07459_),
    .A2(_07475_),
    .B1(_07478_),
    .Y(_07865_));
 sky130_fd_sc_hd__a21oi_2 _18222_ (.A1(_07414_),
    .A2(_07423_),
    .B1(_07420_),
    .Y(_07866_));
 sky130_fd_sc_hd__a21o_1 _18223_ (.A1(_07414_),
    .A2(_07423_),
    .B1(_07420_),
    .X(_07868_));
 sky130_fd_sc_hd__a32oi_4 _18224_ (.A1(net219),
    .A2(_04559_),
    .A3(net252),
    .B1(_11793_),
    .B2(net10),
    .Y(_07869_));
 sky130_fd_sc_hd__and3_1 _18225_ (.A(_03971_),
    .B(net11),
    .C(net64),
    .X(_07870_));
 sky130_fd_sc_hd__a31oi_4 _18226_ (.A1(net215),
    .A2(net289),
    .A3(net185),
    .B1(_07870_),
    .Y(_07871_));
 sky130_fd_sc_hd__o211ai_2 _18227_ (.A1(_04787_),
    .A2(net208),
    .B1(net291),
    .C1(net211),
    .Y(_07872_));
 sky130_fd_sc_hd__or3b_1 _18228_ (.A(net64),
    .B(_04113_),
    .C_N(net63),
    .X(_07873_));
 sky130_fd_sc_hd__o22a_1 _18229_ (.A1(_04113_),
    .A2(_08283_),
    .B1(_05077_),
    .B2(_08261_),
    .X(_07874_));
 sky130_fd_sc_hd__a21oi_2 _18230_ (.A1(_07872_),
    .A2(_07873_),
    .B1(_07871_),
    .Y(_07875_));
 sky130_fd_sc_hd__o221a_1 _18231_ (.A1(_04113_),
    .A2(_08283_),
    .B1(_05077_),
    .B2(_08261_),
    .C1(_07871_),
    .X(_07876_));
 sky130_fd_sc_hd__nand2_2 _18232_ (.A(_07871_),
    .B(_07874_),
    .Y(_07877_));
 sky130_fd_sc_hd__o21ai_1 _18233_ (.A1(_07875_),
    .A2(_07876_),
    .B1(_07869_),
    .Y(_07879_));
 sky130_fd_sc_hd__a31o_1 _18234_ (.A1(_07871_),
    .A2(_07872_),
    .A3(_07873_),
    .B1(_07869_),
    .X(_07880_));
 sky130_fd_sc_hd__nand3b_2 _18235_ (.A_N(_07875_),
    .B(_07877_),
    .C(_07869_),
    .Y(_07881_));
 sky130_fd_sc_hd__o21bai_2 _18236_ (.A1(_07875_),
    .A2(_07876_),
    .B1_N(_07869_),
    .Y(_07882_));
 sky130_fd_sc_hd__nand3_2 _18237_ (.A(_07881_),
    .B(_07882_),
    .C(_07866_),
    .Y(_07883_));
 sky130_fd_sc_hd__o211ai_4 _18238_ (.A1(_07875_),
    .A2(_07880_),
    .B1(_07879_),
    .C1(_07868_),
    .Y(_07884_));
 sky130_fd_sc_hd__o32a_1 _18239_ (.A1(_02869_),
    .A2(net247),
    .A3(_03957_),
    .B1(_02891_),
    .B2(_04048_),
    .X(_07885_));
 sky130_fd_sc_hd__a32o_1 _18240_ (.A1(_03952_),
    .A2(net232),
    .A3(_02858_),
    .B1(_02880_),
    .B2(net7),
    .X(_07886_));
 sky130_fd_sc_hd__a32o_1 _18241_ (.A1(net228),
    .A2(_01293_),
    .A3(net230),
    .B1(_01315_),
    .B2(net8),
    .X(_07887_));
 sky130_fd_sc_hd__nor2_1 _18242_ (.A(_04069_),
    .B(_12363_),
    .Y(_07888_));
 sky130_fd_sc_hd__a31oi_1 _18243_ (.A1(net223),
    .A2(_12330_),
    .A3(net188),
    .B1(_07888_),
    .Y(_07890_));
 sky130_fd_sc_hd__a31o_1 _18244_ (.A1(net223),
    .A2(_12330_),
    .A3(net188),
    .B1(_07888_),
    .X(_07891_));
 sky130_fd_sc_hd__nand2_2 _18245_ (.A(_07887_),
    .B(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__nor2_1 _18246_ (.A(_07887_),
    .B(_07891_),
    .Y(_07893_));
 sky130_fd_sc_hd__o221ai_2 _18247_ (.A1(_04059_),
    .A2(_01326_),
    .B1(_04133_),
    .B2(_01304_),
    .C1(_07890_),
    .Y(_07894_));
 sky130_fd_sc_hd__a21o_1 _18248_ (.A1(_07892_),
    .A2(_07894_),
    .B1(_07886_),
    .X(_07895_));
 sky130_fd_sc_hd__nand3_1 _18249_ (.A(_07886_),
    .B(_07892_),
    .C(_07894_),
    .Y(_07896_));
 sky130_fd_sc_hd__nand2_2 _18250_ (.A(_07895_),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__a21bo_1 _18251_ (.A1(_07883_),
    .A2(_07884_),
    .B1_N(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__nand4_2 _18252_ (.A(_07883_),
    .B(_07884_),
    .C(_07895_),
    .D(_07896_),
    .Y(_07899_));
 sky130_fd_sc_hd__nand3_1 _18253_ (.A(_07883_),
    .B(_07884_),
    .C(_07897_),
    .Y(_07901_));
 sky130_fd_sc_hd__a21o_1 _18254_ (.A1(_07883_),
    .A2(_07884_),
    .B1(_07897_),
    .X(_07902_));
 sky130_fd_sc_hd__nand4_4 _18255_ (.A(_07478_),
    .B(_07480_),
    .C(_07901_),
    .D(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand3_4 _18256_ (.A(_07865_),
    .B(_07898_),
    .C(_07899_),
    .Y(_07904_));
 sky130_fd_sc_hd__and3_1 _18257_ (.A(_07431_),
    .B(_07444_),
    .C(_07445_),
    .X(_07905_));
 sky130_fd_sc_hd__a31oi_4 _18258_ (.A1(_07431_),
    .A2(_07444_),
    .A3(_07445_),
    .B1(_07429_),
    .Y(_07906_));
 sky130_fd_sc_hd__a21oi_2 _18259_ (.A1(_07903_),
    .A2(_07904_),
    .B1(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__a21o_1 _18260_ (.A1(_07903_),
    .A2(_07904_),
    .B1(_07906_),
    .X(_07908_));
 sky130_fd_sc_hd__and3_1 _18261_ (.A(_07903_),
    .B(_07904_),
    .C(_07906_),
    .X(_07909_));
 sky130_fd_sc_hd__nand3_1 _18262_ (.A(_07903_),
    .B(_07904_),
    .C(_07906_),
    .Y(_07910_));
 sky130_fd_sc_hd__a211oi_2 _18263_ (.A1(_07903_),
    .A2(_07904_),
    .B1(_07905_),
    .C1(_07429_),
    .Y(_07912_));
 sky130_fd_sc_hd__o211a_1 _18264_ (.A1(_07429_),
    .A2(_07905_),
    .B1(_07904_),
    .C1(_07903_),
    .X(_07913_));
 sky130_fd_sc_hd__o211ai_4 _18265_ (.A1(_07907_),
    .A2(_07909_),
    .B1(_07862_),
    .C1(_07864_),
    .Y(_07914_));
 sky130_fd_sc_hd__o2bb2ai_4 _18266_ (.A1_N(_07862_),
    .A2_N(_07864_),
    .B1(_07912_),
    .B2(_07913_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand3_1 _18267_ (.A(_07862_),
    .B(_07908_),
    .C(_07910_),
    .Y(_07916_));
 sky130_fd_sc_hd__o2111a_2 _18268_ (.A1(_07543_),
    .A2(_07545_),
    .B1(_07551_),
    .C1(_07914_),
    .D1(_07915_),
    .X(_07917_));
 sky130_fd_sc_hd__o2111ai_4 _18269_ (.A1(_07543_),
    .A2(_07545_),
    .B1(_07551_),
    .C1(_07914_),
    .D1(_07915_),
    .Y(_07918_));
 sky130_fd_sc_hd__a22oi_4 _18270_ (.A1(_07547_),
    .A2(_07551_),
    .B1(_07914_),
    .B2(_07915_),
    .Y(_07919_));
 sky130_fd_sc_hd__a22o_2 _18271_ (.A1(_07547_),
    .A2(_07551_),
    .B1(_07914_),
    .B2(_07915_),
    .X(_07920_));
 sky130_fd_sc_hd__o21ai_1 _18272_ (.A1(_07917_),
    .A2(_07919_),
    .B1(_07761_),
    .Y(_07921_));
 sky130_fd_sc_hd__o211ai_2 _18273_ (.A1(_07759_),
    .A2(_07760_),
    .B1(_07918_),
    .C1(_07920_),
    .Y(_07923_));
 sky130_fd_sc_hd__o22ai_4 _18274_ (.A1(_07759_),
    .A2(_07760_),
    .B1(_07917_),
    .B2(_07919_),
    .Y(_07924_));
 sky130_fd_sc_hd__nand2_1 _18275_ (.A(_07761_),
    .B(_07918_),
    .Y(_07925_));
 sky130_fd_sc_hd__nand3_4 _18276_ (.A(_07920_),
    .B(_07761_),
    .C(_07918_),
    .Y(_07926_));
 sky130_fd_sc_hd__a22oi_2 _18277_ (.A1(_07559_),
    .A2(_07563_),
    .B1(_07921_),
    .B2(_07923_),
    .Y(_07927_));
 sky130_fd_sc_hd__nand3_2 _18278_ (.A(_07678_),
    .B(_07924_),
    .C(_07926_),
    .Y(_07928_));
 sky130_fd_sc_hd__a21oi_4 _18279_ (.A1(_07924_),
    .A2(_07926_),
    .B1(_07678_),
    .Y(_07929_));
 sky130_fd_sc_hd__nand4_2 _18280_ (.A(_07559_),
    .B(_07563_),
    .C(_07921_),
    .D(_07923_),
    .Y(_07930_));
 sky130_fd_sc_hd__a32oi_4 _18281_ (.A1(_07678_),
    .A2(_07924_),
    .A3(_07926_),
    .B1(_07674_),
    .B2(_07671_),
    .Y(_07931_));
 sky130_fd_sc_hd__o21ai_1 _18282_ (.A1(_07677_),
    .A2(_07929_),
    .B1(_07928_),
    .Y(_07932_));
 sky130_fd_sc_hd__o211ai_2 _18283_ (.A1(_07670_),
    .A2(_07673_),
    .B1(_07928_),
    .C1(_07930_),
    .Y(_07934_));
 sky130_fd_sc_hd__o22ai_2 _18284_ (.A1(_07675_),
    .A2(_07676_),
    .B1(_07927_),
    .B2(_07929_),
    .Y(_07935_));
 sky130_fd_sc_hd__o22ai_2 _18285_ (.A1(_07670_),
    .A2(_07673_),
    .B1(_07927_),
    .B2(_07929_),
    .Y(_07936_));
 sky130_fd_sc_hd__o2111ai_4 _18286_ (.A1(_07672_),
    .A2(_07665_),
    .B1(_07671_),
    .C1(_07928_),
    .D1(_07930_),
    .Y(_07937_));
 sky130_fd_sc_hd__o2bb2ai_1 _18287_ (.A1_N(_07326_),
    .A2_N(_07569_),
    .B1(_07566_),
    .B2(_07564_),
    .Y(_07938_));
 sky130_fd_sc_hd__a21oi_2 _18288_ (.A1(_07569_),
    .A2(_07326_),
    .B1(_07567_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand3_2 _18289_ (.A(_07934_),
    .B(_07935_),
    .C(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__and3_1 _18290_ (.A(_07936_),
    .B(_07938_),
    .C(_07937_),
    .X(_07941_));
 sky130_fd_sc_hd__nand3_2 _18291_ (.A(_07936_),
    .B(_07938_),
    .C(_07937_),
    .Y(_07942_));
 sky130_fd_sc_hd__a21o_1 _18292_ (.A1(_07940_),
    .A2(_07942_),
    .B1(_07602_),
    .X(_07943_));
 sky130_fd_sc_hd__a31oi_2 _18293_ (.A1(_07934_),
    .A2(_07935_),
    .A3(_07939_),
    .B1(_07604_),
    .Y(_07945_));
 sky130_fd_sc_hd__o211ai_1 _18294_ (.A1(_07317_),
    .A2(_07325_),
    .B1(_07940_),
    .C1(_07942_),
    .Y(_07946_));
 sky130_fd_sc_hd__a21o_1 _18295_ (.A1(_07940_),
    .A2(_07942_),
    .B1(_07604_),
    .X(_07947_));
 sky130_fd_sc_hd__nand3_1 _18296_ (.A(_07940_),
    .B(_07942_),
    .C(_07604_),
    .Y(_07948_));
 sky130_fd_sc_hd__nand2_1 _18297_ (.A(_07581_),
    .B(_07584_),
    .Y(_07949_));
 sky130_fd_sc_hd__a21oi_1 _18298_ (.A1(_07579_),
    .A2(_07583_),
    .B1(_07580_),
    .Y(_07950_));
 sky130_fd_sc_hd__nand3_2 _18299_ (.A(_07947_),
    .B(_07948_),
    .C(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__a21oi_1 _18300_ (.A1(_07947_),
    .A2(_07948_),
    .B1(_07950_),
    .Y(_07952_));
 sky130_fd_sc_hd__nand4_2 _18301_ (.A(_07579_),
    .B(_07943_),
    .C(_07946_),
    .D(_07949_),
    .Y(_07953_));
 sky130_fd_sc_hd__nand2_1 _18302_ (.A(_07951_),
    .B(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__nand3_1 _18303_ (.A(_07591_),
    .B(_07951_),
    .C(_07953_),
    .Y(_07956_));
 sky130_fd_sc_hd__o2bb2ai_2 _18304_ (.A1_N(_07951_),
    .A2_N(_07953_),
    .B1(_07262_),
    .B2(_07589_),
    .Y(_07957_));
 sky130_fd_sc_hd__a21o_1 _18305_ (.A1(_07956_),
    .A2(_07957_),
    .B1(_07601_),
    .X(_07958_));
 sky130_fd_sc_hd__o2111a_1 _18306_ (.A1(_07591_),
    .A2(_07595_),
    .B1(_07956_),
    .C1(_07957_),
    .D1(_07594_),
    .X(_07959_));
 sky130_fd_sc_hd__nand3_1 _18307_ (.A(_07601_),
    .B(_07956_),
    .C(_07957_),
    .Y(_07960_));
 sky130_fd_sc_hd__and2_1 _18308_ (.A(_07958_),
    .B(_07960_),
    .X(net86));
 sky130_fd_sc_hd__a21oi_2 _18309_ (.A1(_07602_),
    .A2(_07940_),
    .B1(_07941_),
    .Y(_07961_));
 sky130_fd_sc_hd__o21ai_1 _18310_ (.A1(_07656_),
    .A2(_07638_),
    .B1(_07641_),
    .Y(_07962_));
 sky130_fd_sc_hd__inv_2 _18311_ (.A(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__o2bb2a_1 _18312_ (.A1_N(_07758_),
    .A2_N(_07754_),
    .B1(_07752_),
    .B2(_07755_),
    .X(_07964_));
 sky130_fd_sc_hd__a2bb2o_1 _18313_ (.A1_N(_07752_),
    .A2_N(_07755_),
    .B1(_07758_),
    .B2(_07754_),
    .X(_07966_));
 sky130_fd_sc_hd__nand2_1 _18314_ (.A(_07632_),
    .B(_07635_),
    .Y(_07967_));
 sky130_fd_sc_hd__a21bo_1 _18315_ (.A1(_07608_),
    .A2(_07627_),
    .B1_N(_07626_),
    .X(_07968_));
 sky130_fd_sc_hd__a21oi_1 _18316_ (.A1(_07612_),
    .A2(_07620_),
    .B1(_07618_),
    .Y(_07969_));
 sky130_fd_sc_hd__a21o_1 _18317_ (.A1(_07612_),
    .A2(_07620_),
    .B1(_07618_),
    .X(_07970_));
 sky130_fd_sc_hd__nand2_1 _18318_ (.A(_07705_),
    .B(_07700_),
    .Y(_07971_));
 sky130_fd_sc_hd__a32oi_2 _18319_ (.A1(_06863_),
    .A2(net301),
    .A3(net266),
    .B1(net27),
    .B2(_06865_),
    .Y(_07972_));
 sky130_fd_sc_hd__a32o_1 _18320_ (.A1(net266),
    .A2(net301),
    .A3(_06863_),
    .B1(_06865_),
    .B2(net27),
    .X(_07973_));
 sky130_fd_sc_hd__o211ai_2 _18321_ (.A1(_04747_),
    .A2(_05436_),
    .B1(net273),
    .C1(_05414_),
    .Y(_07974_));
 sky130_fd_sc_hd__or3b_2 _18322_ (.A(_03725_),
    .B(net50),
    .C_N(net49),
    .X(_07975_));
 sky130_fd_sc_hd__nand3_1 _18323_ (.A(_05841_),
    .B(net265),
    .C(_06026_),
    .Y(_07977_));
 sky130_fd_sc_hd__or3b_2 _18324_ (.A(_03835_),
    .B(net49),
    .C_N(net48),
    .X(_07978_));
 sky130_fd_sc_hd__a22oi_1 _18325_ (.A1(_07974_),
    .A2(_07975_),
    .B1(_07977_),
    .B2(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__a22o_1 _18326_ (.A1(_07974_),
    .A2(_07975_),
    .B1(_07977_),
    .B2(_07978_),
    .X(_07980_));
 sky130_fd_sc_hd__and4_1 _18327_ (.A(_07974_),
    .B(_07975_),
    .C(_07977_),
    .D(_07978_),
    .X(_07981_));
 sky130_fd_sc_hd__nand4_2 _18328_ (.A(_07974_),
    .B(_07975_),
    .C(_07977_),
    .D(_07978_),
    .Y(_07982_));
 sky130_fd_sc_hd__nor3b_1 _18329_ (.A(_07972_),
    .B(_07979_),
    .C_N(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__nand3_1 _18330_ (.A(_07973_),
    .B(_07980_),
    .C(_07982_),
    .Y(_07984_));
 sky130_fd_sc_hd__a21oi_1 _18331_ (.A1(_07980_),
    .A2(_07982_),
    .B1(_07973_),
    .Y(_07985_));
 sky130_fd_sc_hd__o21ai_1 _18332_ (.A1(_07979_),
    .A2(_07981_),
    .B1(_07972_),
    .Y(_07986_));
 sky130_fd_sc_hd__nand4_2 _18333_ (.A(_07706_),
    .B(_07971_),
    .C(_07984_),
    .D(_07986_),
    .Y(_07988_));
 sky130_fd_sc_hd__o2bb2ai_2 _18334_ (.A1_N(_07706_),
    .A2_N(_07971_),
    .B1(_07983_),
    .B2(_07985_),
    .Y(_07989_));
 sky130_fd_sc_hd__a21oi_1 _18335_ (.A1(_07988_),
    .A2(_07989_),
    .B1(_07970_),
    .Y(_07990_));
 sky130_fd_sc_hd__o211a_1 _18336_ (.A1(_07618_),
    .A2(_07623_),
    .B1(_07988_),
    .C1(_07989_),
    .X(_07991_));
 sky130_fd_sc_hd__and3_1 _18337_ (.A(_07988_),
    .B(_07989_),
    .C(_07969_),
    .X(_07992_));
 sky130_fd_sc_hd__a21oi_1 _18338_ (.A1(_07988_),
    .A2(_07989_),
    .B1(_07969_),
    .Y(_07993_));
 sky130_fd_sc_hd__o211ai_2 _18339_ (.A1(_07990_),
    .A2(_07991_),
    .B1(_07699_),
    .C1(_07712_),
    .Y(_07994_));
 sky130_fd_sc_hd__o2bb2a_1 _18340_ (.A1_N(_07699_),
    .A2_N(_07712_),
    .B1(_07992_),
    .B2(_07993_),
    .X(_07995_));
 sky130_fd_sc_hd__o2bb2ai_1 _18341_ (.A1_N(_07699_),
    .A2_N(_07712_),
    .B1(_07992_),
    .B2(_07993_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_1 _18342_ (.A(_07994_),
    .B(_07968_),
    .Y(_07997_));
 sky130_fd_sc_hd__and3_1 _18343_ (.A(_07994_),
    .B(_07996_),
    .C(_07968_),
    .X(_07999_));
 sky130_fd_sc_hd__a21oi_1 _18344_ (.A1(_07994_),
    .A2(_07996_),
    .B1(_07968_),
    .Y(_08000_));
 sky130_fd_sc_hd__a21o_1 _18345_ (.A1(_07994_),
    .A2(_07996_),
    .B1(_07968_),
    .X(_08001_));
 sky130_fd_sc_hd__o211a_2 _18346_ (.A1(_07999_),
    .A2(_08000_),
    .B1(_07632_),
    .C1(_07635_),
    .X(_08002_));
 sky130_fd_sc_hd__o211ai_2 _18347_ (.A1(_07999_),
    .A2(_08000_),
    .B1(_07632_),
    .C1(_07635_),
    .Y(_08003_));
 sky130_fd_sc_hd__o211ai_4 _18348_ (.A1(_07997_),
    .A2(_07995_),
    .B1(_07967_),
    .C1(_08001_),
    .Y(_08004_));
 sky130_fd_sc_hd__nor2_8 _18349_ (.A(net54),
    .B(_04266_),
    .Y(_08005_));
 sky130_fd_sc_hd__and2_4 _18350_ (.A(_04266_),
    .B(net54),
    .X(_08006_));
 sky130_fd_sc_hd__nand2_8 _18351_ (.A(_04266_),
    .B(net54),
    .Y(_08007_));
 sky130_fd_sc_hd__o21a_1 _18352_ (.A1(_08005_),
    .A2(_08006_),
    .B1(net1),
    .X(_08008_));
 sky130_fd_sc_hd__o21ai_1 _18353_ (.A1(_07644_),
    .A2(_07649_),
    .B1(_07648_),
    .Y(_08010_));
 sky130_fd_sc_hd__a22oi_1 _18354_ (.A1(net12),
    .A2(_07643_),
    .B1(_04539_),
    .B2(_07642_),
    .Y(_08011_));
 sky130_fd_sc_hd__a22o_1 _18355_ (.A1(net12),
    .A2(_07643_),
    .B1(_04539_),
    .B2(_07642_),
    .X(_08012_));
 sky130_fd_sc_hd__or3b_1 _18356_ (.A(_03396_),
    .B(net53),
    .C_N(net52),
    .X(_08013_));
 sky130_fd_sc_hd__a211o_4 _18357_ (.A1(_03176_),
    .A2(_04430_),
    .B1(_07306_),
    .C1(_04408_),
    .X(_08014_));
 sky130_fd_sc_hd__nand3_1 _18358_ (.A(net313),
    .B(_04747_),
    .C(_07223_),
    .Y(_08015_));
 sky130_fd_sc_hd__nand2_1 _18359_ (.A(net26),
    .B(_07225_),
    .Y(_08016_));
 sky130_fd_sc_hd__a22oi_2 _18360_ (.A1(_08013_),
    .A2(_08014_),
    .B1(_08015_),
    .B2(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__and4_1 _18361_ (.A(_08013_),
    .B(_08014_),
    .C(_08015_),
    .D(_08016_),
    .X(_08018_));
 sky130_fd_sc_hd__nand4_1 _18362_ (.A(_08013_),
    .B(_08014_),
    .C(_08015_),
    .D(_08016_),
    .Y(_08019_));
 sky130_fd_sc_hd__o21ai_1 _18363_ (.A1(_08017_),
    .A2(_08018_),
    .B1(_08011_),
    .Y(_08021_));
 sky130_fd_sc_hd__or3_1 _18364_ (.A(_08011_),
    .B(_08017_),
    .C(_08018_),
    .X(_08022_));
 sky130_fd_sc_hd__nand3_2 _18365_ (.A(_08010_),
    .B(_08021_),
    .C(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__a21o_1 _18366_ (.A1(_08021_),
    .A2(_08022_),
    .B1(_08010_),
    .X(_08024_));
 sky130_fd_sc_hd__a21oi_1 _18367_ (.A1(_08023_),
    .A2(_08024_),
    .B1(_08008_),
    .Y(_08025_));
 sky130_fd_sc_hd__o211a_1 _18368_ (.A1(_08005_),
    .A2(_08006_),
    .B1(net1),
    .C1(_08024_),
    .X(_08026_));
 sky130_fd_sc_hd__nand2_1 _18369_ (.A(_08024_),
    .B(_08008_),
    .Y(_08027_));
 sky130_fd_sc_hd__a21o_2 _18370_ (.A1(_08026_),
    .A2(_08023_),
    .B1(_08025_),
    .X(_08028_));
 sky130_fd_sc_hd__or2_1 _18371_ (.A(_07654_),
    .B(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__a31o_1 _18372_ (.A1(_07309_),
    .A2(_07310_),
    .A3(_07653_),
    .B1(_08028_),
    .X(_08030_));
 sky130_fd_sc_hd__nand4_2 _18373_ (.A(_07310_),
    .B(_08028_),
    .C(_07653_),
    .D(_07309_),
    .Y(_08032_));
 sky130_fd_sc_hd__nand2_1 _18374_ (.A(_08030_),
    .B(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__a21o_1 _18375_ (.A1(_08003_),
    .A2(_08004_),
    .B1(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__nand3_1 _18376_ (.A(_08003_),
    .B(_08033_),
    .C(_08004_),
    .Y(_08035_));
 sky130_fd_sc_hd__a22o_1 _18377_ (.A1(_08003_),
    .A2(_08004_),
    .B1(_08030_),
    .B2(_08032_),
    .X(_08036_));
 sky130_fd_sc_hd__nand4_1 _18378_ (.A(_08003_),
    .B(_08004_),
    .C(_08030_),
    .D(_08032_),
    .Y(_08037_));
 sky130_fd_sc_hd__and3_2 _18379_ (.A(_07966_),
    .B(_08034_),
    .C(_08035_),
    .X(_08038_));
 sky130_fd_sc_hd__and3_1 _18380_ (.A(_07964_),
    .B(_08036_),
    .C(_08037_),
    .X(_08039_));
 sky130_fd_sc_hd__o21ai_4 _18381_ (.A1(_08038_),
    .A2(_08039_),
    .B1(_07963_),
    .Y(_08040_));
 sky130_fd_sc_hd__a31o_1 _18382_ (.A1(_07964_),
    .A2(_08036_),
    .A3(_08037_),
    .B1(_07963_),
    .X(_08041_));
 sky130_fd_sc_hd__a31o_1 _18383_ (.A1(_07966_),
    .A2(_08034_),
    .A3(_08035_),
    .B1(_08041_),
    .X(_08043_));
 sky130_fd_sc_hd__o22a_1 _18384_ (.A1(_07640_),
    .A2(_07659_),
    .B1(_08038_),
    .B2(_08039_),
    .X(_08044_));
 sky130_fd_sc_hd__nor4_1 _18385_ (.A(_07640_),
    .B(_07659_),
    .C(_08038_),
    .D(_08039_),
    .Y(_08045_));
 sky130_fd_sc_hd__o21ai_1 _18386_ (.A1(_08038_),
    .A2(_08041_),
    .B1(_08040_),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_1 _18387_ (.A(_07761_),
    .B(_07919_),
    .Y(_08047_));
 sky130_fd_sc_hd__a21o_1 _18388_ (.A1(_07761_),
    .A2(_07918_),
    .B1(_07919_),
    .X(_08048_));
 sky130_fd_sc_hd__a31o_2 _18389_ (.A1(_07865_),
    .A2(_07898_),
    .A3(_07899_),
    .B1(_07906_),
    .X(_08049_));
 sky130_fd_sc_hd__o2bb2ai_2 _18390_ (.A1_N(_07717_),
    .A2_N(_07739_),
    .B1(_07740_),
    .B2(_07737_),
    .Y(_08050_));
 sky130_fd_sc_hd__a21oi_1 _18391_ (.A1(_07887_),
    .A2(_07891_),
    .B1(_07886_),
    .Y(_08051_));
 sky130_fd_sc_hd__o21ai_1 _18392_ (.A1(_07887_),
    .A2(_07891_),
    .B1(_07886_),
    .Y(_08052_));
 sky130_fd_sc_hd__o21ai_1 _18393_ (.A1(_07885_),
    .A2(_07893_),
    .B1(_07892_),
    .Y(_08054_));
 sky130_fd_sc_hd__a32o_1 _18394_ (.A1(_00625_),
    .A2(net250),
    .A3(net280),
    .B1(_04269_),
    .B2(net5),
    .X(_08055_));
 sky130_fd_sc_hd__or3b_1 _18395_ (.A(_04026_),
    .B(net40),
    .C_N(net39),
    .X(_08056_));
 sky130_fd_sc_hd__o211ai_2 _18396_ (.A1(net254),
    .A2(_02442_),
    .B1(net281),
    .C1(_02421_),
    .Y(_08057_));
 sky130_fd_sc_hd__a32oi_4 _18397_ (.A1(_02421_),
    .A2(net249),
    .A3(net281),
    .B1(_04217_),
    .B2(net6),
    .Y(_08058_));
 sky130_fd_sc_hd__nor2_1 _18398_ (.A(_04048_),
    .B(_03737_),
    .Y(_08059_));
 sky130_fd_sc_hd__o311a_1 _18399_ (.A1(net260),
    .A2(_11387_),
    .A3(_03954_),
    .B1(net285),
    .C1(_03952_),
    .X(_08060_));
 sky130_fd_sc_hd__o211ai_1 _18400_ (.A1(net254),
    .A2(_03954_),
    .B1(net285),
    .C1(_03952_),
    .Y(_08061_));
 sky130_fd_sc_hd__a31oi_2 _18401_ (.A1(_03952_),
    .A2(net232),
    .A3(net285),
    .B1(_08059_),
    .Y(_08062_));
 sky130_fd_sc_hd__o211ai_1 _18402_ (.A1(_04026_),
    .A2(_04218_),
    .B1(_08057_),
    .C1(_08061_),
    .Y(_08063_));
 sky130_fd_sc_hd__nand2_2 _18403_ (.A(_08058_),
    .B(_08062_),
    .Y(_08065_));
 sky130_fd_sc_hd__o2bb2ai_2 _18404_ (.A1_N(_08056_),
    .A2_N(_08057_),
    .B1(_08059_),
    .B2(_08060_),
    .Y(_08066_));
 sky130_fd_sc_hd__o21a_1 _18405_ (.A1(_08058_),
    .A2(_08062_),
    .B1(_08055_),
    .X(_08067_));
 sky130_fd_sc_hd__o211a_1 _18406_ (.A1(_08059_),
    .A2(_08063_),
    .B1(_08066_),
    .C1(_08055_),
    .X(_08068_));
 sky130_fd_sc_hd__o21ai_1 _18407_ (.A1(_08059_),
    .A2(_08063_),
    .B1(_08067_),
    .Y(_08069_));
 sky130_fd_sc_hd__a21oi_4 _18408_ (.A1(_08065_),
    .A2(_08066_),
    .B1(_08055_),
    .Y(_08070_));
 sky130_fd_sc_hd__a221oi_4 _18409_ (.A1(_08067_),
    .A2(_08065_),
    .B1(_08052_),
    .B2(_07892_),
    .C1(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__nand3b_2 _18410_ (.A_N(_08070_),
    .B(_08054_),
    .C(_08069_),
    .Y(_08072_));
 sky130_fd_sc_hd__o22a_1 _18411_ (.A1(_07893_),
    .A2(_08051_),
    .B1(_08068_),
    .B2(_08070_),
    .X(_08073_));
 sky130_fd_sc_hd__o221ai_4 _18412_ (.A1(_07885_),
    .A2(_07893_),
    .B1(_08068_),
    .B2(_08070_),
    .C1(_07892_),
    .Y(_08074_));
 sky130_fd_sc_hd__o22ai_2 _18413_ (.A1(_07727_),
    .A2(_07733_),
    .B1(_08071_),
    .B2(_08073_),
    .Y(_08076_));
 sky130_fd_sc_hd__o2111ai_4 _18414_ (.A1(_07720_),
    .A2(_07729_),
    .B1(_08072_),
    .C1(_08074_),
    .D1(_07728_),
    .Y(_08077_));
 sky130_fd_sc_hd__o21ai_1 _18415_ (.A1(_07727_),
    .A2(_07733_),
    .B1(_08074_),
    .Y(_08078_));
 sky130_fd_sc_hd__o21ai_1 _18416_ (.A1(_08071_),
    .A2(_08073_),
    .B1(_07734_),
    .Y(_08079_));
 sky130_fd_sc_hd__o211ai_4 _18417_ (.A1(_08071_),
    .A2(_08078_),
    .B1(_08050_),
    .C1(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__nand3b_4 _18418_ (.A_N(_08050_),
    .B(_08076_),
    .C(_08077_),
    .Y(_08081_));
 sky130_fd_sc_hd__a21oi_1 _18419_ (.A1(_07682_),
    .A2(_07692_),
    .B1(_07689_),
    .Y(_08082_));
 sky130_fd_sc_hd__o211ai_1 _18420_ (.A1(_11387_),
    .A2(_12988_),
    .B1(net279),
    .C1(net234),
    .Y(_08083_));
 sky130_fd_sc_hd__or3b_1 _18421_ (.A(_04004_),
    .B(net42),
    .C_N(net41),
    .X(_08084_));
 sky130_fd_sc_hd__a32oi_4 _18422_ (.A1(net234),
    .A2(net251),
    .A3(net279),
    .B1(_04482_),
    .B2(net4),
    .Y(_08085_));
 sky130_fd_sc_hd__or3b_1 _18423_ (.A(_03982_),
    .B(net43),
    .C_N(net42),
    .X(_08087_));
 sky130_fd_sc_hd__o211ai_1 _18424_ (.A1(net260),
    .A2(_11387_),
    .B1(net243),
    .C1(_11354_),
    .Y(_08088_));
 sky130_fd_sc_hd__o221ai_4 _18425_ (.A1(_11453_),
    .A2(_04896_),
    .B1(_04898_),
    .B2(_03982_),
    .C1(_08085_),
    .Y(_08089_));
 sky130_fd_sc_hd__a21oi_1 _18426_ (.A1(_08087_),
    .A2(_08088_),
    .B1(_08085_),
    .Y(_08090_));
 sky130_fd_sc_hd__a22o_1 _18427_ (.A1(_08083_),
    .A2(_08084_),
    .B1(_08087_),
    .B2(_08088_),
    .X(_08091_));
 sky130_fd_sc_hd__and3_1 _18428_ (.A(_04124_),
    .B(net43),
    .C(net2),
    .X(_08092_));
 sky130_fd_sc_hd__o311a_1 _18429_ (.A1(_04747_),
    .A2(net264),
    .A3(_09665_),
    .B1(_04985_),
    .C1(_09698_),
    .X(_08093_));
 sky130_fd_sc_hd__a31o_1 _18430_ (.A1(net255),
    .A2(_09698_),
    .A3(_04985_),
    .B1(_08092_),
    .X(_08094_));
 sky130_fd_sc_hd__a21o_1 _18431_ (.A1(_08089_),
    .A2(_08091_),
    .B1(_08094_),
    .X(_08095_));
 sky130_fd_sc_hd__o211ai_1 _18432_ (.A1(_08092_),
    .A2(_08093_),
    .B1(_08089_),
    .C1(_08091_),
    .Y(_08096_));
 sky130_fd_sc_hd__o2bb2ai_1 _18433_ (.A1_N(_08089_),
    .A2_N(_08091_),
    .B1(_08092_),
    .B2(_08093_),
    .Y(_08098_));
 sky130_fd_sc_hd__nand3b_1 _18434_ (.A_N(_08094_),
    .B(_08091_),
    .C(_08089_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand4_1 _18435_ (.A(_07690_),
    .B(_07696_),
    .C(_08098_),
    .D(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__a21oi_2 _18436_ (.A1(_08098_),
    .A2(_08099_),
    .B1(_08082_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand3b_1 _18437_ (.A_N(_08082_),
    .B(_08095_),
    .C(_08096_),
    .Y(_08102_));
 sky130_fd_sc_hd__o22a_1 _18438_ (.A1(_06552_),
    .A2(_05763_),
    .B1(_05766_),
    .B2(_03916_),
    .X(_08103_));
 sky130_fd_sc_hd__nand3_1 _18439_ (.A(_07242_),
    .B(net257),
    .C(_05462_),
    .Y(_08104_));
 sky130_fd_sc_hd__a32oi_2 _18440_ (.A1(_07242_),
    .A2(net257),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net31),
    .Y(_08105_));
 sky130_fd_sc_hd__or3_1 _18441_ (.A(net46),
    .B(_04124_),
    .C(_03949_),
    .X(_08106_));
 sky130_fd_sc_hd__o211ai_2 _18442_ (.A1(net260),
    .A2(_08656_),
    .B1(net276),
    .C1(_08700_),
    .Y(_08107_));
 sky130_fd_sc_hd__a21oi_1 _18443_ (.A1(_08106_),
    .A2(_08107_),
    .B1(_08105_),
    .Y(_08109_));
 sky130_fd_sc_hd__a21o_1 _18444_ (.A1(_08106_),
    .A2(_08107_),
    .B1(_08105_),
    .X(_08110_));
 sky130_fd_sc_hd__o2111a_1 _18445_ (.A1(_03938_),
    .A2(_05465_),
    .B1(_08104_),
    .C1(_08106_),
    .D1(_08107_),
    .X(_08111_));
 sky130_fd_sc_hd__o21bai_1 _18446_ (.A1(_08109_),
    .A2(_08111_),
    .B1_N(_08103_),
    .Y(_08112_));
 sky130_fd_sc_hd__nand3b_1 _18447_ (.A_N(_08111_),
    .B(_08103_),
    .C(_08110_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand2_1 _18448_ (.A(_08112_),
    .B(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__a21o_1 _18449_ (.A1(_08100_),
    .A2(_08102_),
    .B1(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__inv_2 _18450_ (.A(_08115_),
    .Y(_08116_));
 sky130_fd_sc_hd__a32o_1 _18451_ (.A1(_08098_),
    .A2(_08099_),
    .A3(_08082_),
    .B1(_08112_),
    .B2(_08113_),
    .X(_08117_));
 sky130_fd_sc_hd__and3_1 _18452_ (.A(_08100_),
    .B(_08102_),
    .C(_08114_),
    .X(_08118_));
 sky130_fd_sc_hd__o21ai_1 _18453_ (.A1(_08101_),
    .A2(_08117_),
    .B1(_08115_),
    .Y(_08120_));
 sky130_fd_sc_hd__a21boi_1 _18454_ (.A1(_08080_),
    .A2(_08081_),
    .B1_N(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__o2bb2ai_1 _18455_ (.A1_N(_08080_),
    .A2_N(_08081_),
    .B1(_08116_),
    .B2(_08118_),
    .Y(_08122_));
 sky130_fd_sc_hd__o2111a_1 _18456_ (.A1(_08101_),
    .A2(_08117_),
    .B1(_08115_),
    .C1(_08080_),
    .D1(_08081_),
    .X(_08123_));
 sky130_fd_sc_hd__o2111ai_4 _18457_ (.A1(_08101_),
    .A2(_08117_),
    .B1(_08115_),
    .C1(_08080_),
    .D1(_08081_),
    .Y(_08124_));
 sky130_fd_sc_hd__o2bb2ai_4 _18458_ (.A1_N(_07903_),
    .A2_N(_08049_),
    .B1(_08121_),
    .B2(_08123_),
    .Y(_08125_));
 sky130_fd_sc_hd__nand4_4 _18459_ (.A(_07903_),
    .B(_08049_),
    .C(_08122_),
    .D(_08124_),
    .Y(_08126_));
 sky130_fd_sc_hd__inv_2 _18460_ (.A(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__a21bo_2 _18461_ (.A1(_07714_),
    .A2(_07748_),
    .B1_N(_07749_),
    .X(_08128_));
 sky130_fd_sc_hd__a21oi_1 _18462_ (.A1(_08125_),
    .A2(_08126_),
    .B1(_08128_),
    .Y(_08129_));
 sky130_fd_sc_hd__a21o_1 _18463_ (.A1(_08125_),
    .A2(_08126_),
    .B1(_08128_),
    .X(_08131_));
 sky130_fd_sc_hd__nand2_2 _18464_ (.A(_08125_),
    .B(_08128_),
    .Y(_08132_));
 sky130_fd_sc_hd__and3_1 _18465_ (.A(_08125_),
    .B(_08126_),
    .C(_08128_),
    .X(_08133_));
 sky130_fd_sc_hd__o21ai_4 _18466_ (.A1(_08127_),
    .A2(_08132_),
    .B1(_08131_),
    .Y(_08134_));
 sky130_fd_sc_hd__o21a_1 _18467_ (.A1(_07907_),
    .A2(_07909_),
    .B1(_07864_),
    .X(_08135_));
 sky130_fd_sc_hd__o21ai_1 _18468_ (.A1(_07907_),
    .A2(_07909_),
    .B1(_07864_),
    .Y(_08136_));
 sky130_fd_sc_hd__nand2_1 _18469_ (.A(_07864_),
    .B(_07916_),
    .Y(_08137_));
 sky130_fd_sc_hd__nand2_1 _18470_ (.A(_07862_),
    .B(_08136_),
    .Y(_08138_));
 sky130_fd_sc_hd__a32o_1 _18471_ (.A1(_07811_),
    .A2(_07814_),
    .A3(_07816_),
    .B1(_07851_),
    .B2(_07854_),
    .X(_08139_));
 sky130_fd_sc_hd__a31oi_4 _18472_ (.A1(_07820_),
    .A2(_07847_),
    .A3(_07849_),
    .B1(_07817_),
    .Y(_08140_));
 sky130_fd_sc_hd__a31o_1 _18473_ (.A1(_07820_),
    .A2(_07847_),
    .A3(_07849_),
    .B1(_07817_),
    .X(_08142_));
 sky130_fd_sc_hd__o311a_1 _18474_ (.A1(net231),
    .A2(_04787_),
    .A3(_05551_),
    .B1(_05549_),
    .C1(_07658_),
    .X(_08143_));
 sky130_fd_sc_hd__nor2_1 _18475_ (.A(_04146_),
    .B(_07691_),
    .Y(_08144_));
 sky130_fd_sc_hd__o32a_1 _18476_ (.A1(_07669_),
    .A2(_05548_),
    .A3(net206),
    .B1(_07691_),
    .B2(_04146_),
    .X(_08145_));
 sky130_fd_sc_hd__o311a_1 _18477_ (.A1(_05551_),
    .A2(_05925_),
    .A3(_06220_),
    .B1(_06219_),
    .C1(_05688_),
    .X(_08146_));
 sky130_fd_sc_hd__o211ai_4 _18478_ (.A1(_05927_),
    .A2(_06220_),
    .B1(_05688_),
    .C1(net201),
    .Y(_08147_));
 sky130_fd_sc_hd__nor2_1 _18479_ (.A(_04168_),
    .B(_05720_),
    .Y(_08148_));
 sky130_fd_sc_hd__or3b_4 _18480_ (.A(net61),
    .B(_04168_),
    .C_N(net60),
    .X(_08149_));
 sky130_fd_sc_hd__o221ai_4 _18481_ (.A1(net232),
    .A2(_05927_),
    .B1(_04157_),
    .B2(net206),
    .C1(net292),
    .Y(_08150_));
 sky130_fd_sc_hd__or3b_2 _18482_ (.A(net62),
    .B(_04157_),
    .C_N(net61),
    .X(_08151_));
 sky130_fd_sc_hd__o31ai_2 _18483_ (.A1(_06837_),
    .A2(net205),
    .A3(_05932_),
    .B1(_08151_),
    .Y(_08153_));
 sky130_fd_sc_hd__a22oi_4 _18484_ (.A1(_08147_),
    .A2(_08149_),
    .B1(_08150_),
    .B2(_08151_),
    .Y(_08154_));
 sky130_fd_sc_hd__o21ai_4 _18485_ (.A1(_08146_),
    .A2(_08148_),
    .B1(_08153_),
    .Y(_08155_));
 sky130_fd_sc_hd__o2111a_4 _18486_ (.A1(_04157_),
    .A2(_06859_),
    .B1(_08147_),
    .C1(_08149_),
    .D1(_08150_),
    .X(_08156_));
 sky130_fd_sc_hd__o2111ai_4 _18487_ (.A1(_04157_),
    .A2(_06859_),
    .B1(_08147_),
    .C1(_08149_),
    .D1(_08150_),
    .Y(_08157_));
 sky130_fd_sc_hd__a21boi_4 _18488_ (.A1(_08155_),
    .A2(_08157_),
    .B1_N(_08145_),
    .Y(_08158_));
 sky130_fd_sc_hd__o21ai_1 _18489_ (.A1(_08154_),
    .A2(_08156_),
    .B1(_08145_),
    .Y(_08159_));
 sky130_fd_sc_hd__o21ai_4 _18490_ (.A1(_08143_),
    .A2(_08144_),
    .B1(_08155_),
    .Y(_08160_));
 sky130_fd_sc_hd__o211a_2 _18491_ (.A1(_08143_),
    .A2(_08144_),
    .B1(_08155_),
    .C1(_08157_),
    .X(_08161_));
 sky130_fd_sc_hd__o21ai_4 _18492_ (.A1(_08156_),
    .A2(_08160_),
    .B1(_07806_),
    .Y(_08162_));
 sky130_fd_sc_hd__o211ai_4 _18493_ (.A1(_08156_),
    .A2(_08160_),
    .B1(_08159_),
    .C1(_07806_),
    .Y(_08164_));
 sky130_fd_sc_hd__o22ai_4 _18494_ (.A1(_07800_),
    .A2(_07805_),
    .B1(_08158_),
    .B2(_08161_),
    .Y(_08165_));
 sky130_fd_sc_hd__o221a_1 _18495_ (.A1(_04135_),
    .A2(_07691_),
    .B1(_05294_),
    .B2(_07669_),
    .C1(_07831_),
    .X(_08166_));
 sky130_fd_sc_hd__o21ai_4 _18496_ (.A1(_07824_),
    .A2(_07832_),
    .B1(_07831_),
    .Y(_08167_));
 sky130_fd_sc_hd__a21oi_2 _18497_ (.A1(_08164_),
    .A2(_08165_),
    .B1(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__o2bb2ai_4 _18498_ (.A1_N(_08164_),
    .A2_N(_08165_),
    .B1(_08166_),
    .B2(_07832_),
    .Y(_08169_));
 sky130_fd_sc_hd__o211a_1 _18499_ (.A1(_08158_),
    .A2(_08162_),
    .B1(_08167_),
    .C1(_08165_),
    .X(_08170_));
 sky130_fd_sc_hd__o211ai_4 _18500_ (.A1(_08158_),
    .A2(_08162_),
    .B1(_08167_),
    .C1(_08165_),
    .Y(_08171_));
 sky130_fd_sc_hd__nor2_1 _18501_ (.A(_08168_),
    .B(_08170_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_2 _18502_ (.A(_08169_),
    .B(_08171_),
    .Y(_08173_));
 sky130_fd_sc_hd__a22oi_2 _18503_ (.A1(_07808_),
    .A2(_07810_),
    .B1(_07788_),
    .B2(_07763_),
    .Y(_08175_));
 sky130_fd_sc_hd__nand2_1 _18504_ (.A(_07792_),
    .B(_07813_),
    .Y(_08176_));
 sky130_fd_sc_hd__o311a_1 _18505_ (.A1(net245),
    .A2(net241),
    .A3(_06451_),
    .B1(_05227_),
    .C1(net200),
    .X(_08177_));
 sky130_fd_sc_hd__nor2_1 _18506_ (.A(_04179_),
    .B(_05260_),
    .Y(_08178_));
 sky130_fd_sc_hd__a31o_1 _18507_ (.A1(net200),
    .A2(net172),
    .A3(_05227_),
    .B1(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__o211ai_1 _18508_ (.A1(_05931_),
    .A2(_06759_),
    .B1(_04889_),
    .C1(_06757_),
    .Y(_08180_));
 sky130_fd_sc_hd__and3b_1 _18509_ (.A_N(net59),
    .B(net19),
    .C(net58),
    .X(_08181_));
 sky130_fd_sc_hd__or3b_1 _18510_ (.A(net59),
    .B(_04201_),
    .C_N(net58),
    .X(_08182_));
 sky130_fd_sc_hd__a31oi_2 _18511_ (.A1(_06757_),
    .A2(_06762_),
    .A3(_04889_),
    .B1(_08181_),
    .Y(_08183_));
 sky130_fd_sc_hd__o221ai_4 _18512_ (.A1(_05931_),
    .A2(_07074_),
    .B1(_04212_),
    .B2(_06761_),
    .C1(_04627_),
    .Y(_08184_));
 sky130_fd_sc_hd__or3b_1 _18513_ (.A(net58),
    .B(_04212_),
    .C_N(net55),
    .X(_08186_));
 sky130_fd_sc_hd__a21oi_2 _18514_ (.A1(_08184_),
    .A2(_08186_),
    .B1(_08183_),
    .Y(_08187_));
 sky130_fd_sc_hd__a22o_1 _18515_ (.A1(_08180_),
    .A2(_08182_),
    .B1(_08184_),
    .B2(_08186_),
    .X(_08188_));
 sky130_fd_sc_hd__o221a_2 _18516_ (.A1(_04212_),
    .A2(net316),
    .B1(_07079_),
    .B2(_04638_),
    .C1(_08183_),
    .X(_08189_));
 sky130_fd_sc_hd__o211ai_2 _18517_ (.A1(_04212_),
    .A2(net316),
    .B1(_08184_),
    .C1(_08183_),
    .Y(_08190_));
 sky130_fd_sc_hd__a21o_1 _18518_ (.A1(_08188_),
    .A2(_08190_),
    .B1(_08179_),
    .X(_08191_));
 sky130_fd_sc_hd__o21ai_1 _18519_ (.A1(_08177_),
    .A2(_08178_),
    .B1(_08188_),
    .Y(_08192_));
 sky130_fd_sc_hd__o22a_2 _18520_ (.A1(_08177_),
    .A2(_08178_),
    .B1(_08187_),
    .B2(_08189_),
    .X(_08193_));
 sky130_fd_sc_hd__o21ai_1 _18521_ (.A1(_08187_),
    .A2(_08189_),
    .B1(_08179_),
    .Y(_08194_));
 sky130_fd_sc_hd__nor4_2 _18522_ (.A(_08177_),
    .B(_08178_),
    .C(_08187_),
    .D(_08189_),
    .Y(_08195_));
 sky130_fd_sc_hd__nand3b_1 _18523_ (.A_N(_08179_),
    .B(_08188_),
    .C(_08190_),
    .Y(_08197_));
 sky130_fd_sc_hd__nand2_2 _18524_ (.A(_08194_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__o21ai_4 _18525_ (.A1(_08189_),
    .A2(_08192_),
    .B1(_08191_),
    .Y(_08199_));
 sky130_fd_sc_hd__o221a_1 _18526_ (.A1(_04212_),
    .A2(_04375_),
    .B1(_07079_),
    .B2(_04353_),
    .C1(_07778_),
    .X(_08200_));
 sky130_fd_sc_hd__a32oi_1 _18527_ (.A1(_07499_),
    .A2(net167),
    .A3(_04342_),
    .B1(_04364_),
    .B2(net21),
    .Y(_08201_));
 sky130_fd_sc_hd__a32o_2 _18528_ (.A1(_07499_),
    .A2(net167),
    .A3(_04342_),
    .B1(_04364_),
    .B2(net21),
    .X(_08202_));
 sky130_fd_sc_hd__a31oi_4 _18529_ (.A1(_03957_),
    .A2(_05926_),
    .A3(_07766_),
    .B1(_04256_),
    .Y(_08203_));
 sky130_fd_sc_hd__a31o_4 _18530_ (.A1(_03957_),
    .A2(_05926_),
    .A3(_07766_),
    .B1(_04256_),
    .X(_08204_));
 sky130_fd_sc_hd__and3_1 _18531_ (.A(_04223_),
    .B(_04245_),
    .C(_04256_),
    .X(_08205_));
 sky130_fd_sc_hd__or3_4 _18532_ (.A(net21),
    .B(net22),
    .C(net24),
    .X(_08206_));
 sky130_fd_sc_hd__nor3_4 _18533_ (.A(_07767_),
    .B(net24),
    .C(_05931_),
    .Y(_08207_));
 sky130_fd_sc_hd__nand3_4 _18534_ (.A(_05930_),
    .B(_07766_),
    .C(_04256_),
    .Y(_08208_));
 sky130_fd_sc_hd__o21ai_4 _18535_ (.A1(_07076_),
    .A2(net268),
    .B1(_08204_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand3_1 _18536_ (.A(_08204_),
    .B(net163),
    .C(net33),
    .Y(_08210_));
 sky130_fd_sc_hd__or3_2 _18537_ (.A(net44),
    .B(_04245_),
    .C(_03286_),
    .X(_08211_));
 sky130_fd_sc_hd__o211ai_2 _18538_ (.A1(_07076_),
    .A2(_07765_),
    .B1(_04484_),
    .C1(_07771_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand3_4 _18539_ (.A(_08210_),
    .B(_08211_),
    .C(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__and4b_1 _18540_ (.A_N(net44),
    .B(_04256_),
    .C(net22),
    .D(net33),
    .X(_08214_));
 sky130_fd_sc_hd__or4_2 _18541_ (.A(net44),
    .B(net24),
    .C(_04245_),
    .D(_03286_),
    .X(_08215_));
 sky130_fd_sc_hd__nor2_1 _18542_ (.A(_08201_),
    .B(_08214_),
    .Y(_08216_));
 sky130_fd_sc_hd__o311a_4 _18543_ (.A1(_03286_),
    .A2(_08209_),
    .A3(_08211_),
    .B1(_08213_),
    .C1(_08202_),
    .X(_08218_));
 sky130_fd_sc_hd__nand2_1 _18544_ (.A(_08216_),
    .B(_08213_),
    .Y(_08219_));
 sky130_fd_sc_hd__a21oi_2 _18545_ (.A1(_08213_),
    .A2(_08215_),
    .B1(_08202_),
    .Y(_08220_));
 sky130_fd_sc_hd__a21o_1 _18546_ (.A1(_08213_),
    .A2(_08215_),
    .B1(_08202_),
    .X(_08221_));
 sky130_fd_sc_hd__o21ai_4 _18547_ (.A1(_07777_),
    .A2(_07784_),
    .B1(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__a221oi_4 _18548_ (.A1(_08216_),
    .A2(_08213_),
    .B1(_07785_),
    .B2(_07778_),
    .C1(_08220_),
    .Y(_08223_));
 sky130_fd_sc_hd__a31o_1 _18549_ (.A1(_08202_),
    .A2(_08213_),
    .A3(_08215_),
    .B1(_08222_),
    .X(_08224_));
 sky130_fd_sc_hd__a2bb2oi_2 _18550_ (.A1_N(_07776_),
    .A2_N(_08200_),
    .B1(_08219_),
    .B2(_08221_),
    .Y(_08225_));
 sky130_fd_sc_hd__o22ai_4 _18551_ (.A1(_07776_),
    .A2(_08200_),
    .B1(_08218_),
    .B2(_08220_),
    .Y(_08226_));
 sky130_fd_sc_hd__o21ai_1 _18552_ (.A1(_08218_),
    .A2(_08222_),
    .B1(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__o21ai_2 _18553_ (.A1(_08193_),
    .A2(_08195_),
    .B1(_08226_),
    .Y(_08229_));
 sky130_fd_sc_hd__o211ai_4 _18554_ (.A1(_08218_),
    .A2(_08222_),
    .B1(_08198_),
    .C1(_08226_),
    .Y(_08230_));
 sky130_fd_sc_hd__o21ai_2 _18555_ (.A1(_08223_),
    .A2(_08225_),
    .B1(_08199_),
    .Y(_08231_));
 sky130_fd_sc_hd__o211ai_4 _18556_ (.A1(_08218_),
    .A2(_08222_),
    .B1(_08226_),
    .C1(_08199_),
    .Y(_08232_));
 sky130_fd_sc_hd__o22ai_4 _18557_ (.A1(_08193_),
    .A2(_08195_),
    .B1(_08223_),
    .B2(_08225_),
    .Y(_08233_));
 sky130_fd_sc_hd__a22oi_2 _18558_ (.A1(_07792_),
    .A2(_07813_),
    .B1(_08199_),
    .B2(_08227_),
    .Y(_08234_));
 sky130_fd_sc_hd__and3_2 _18559_ (.A(_08231_),
    .B(_08176_),
    .C(_08230_),
    .X(_08235_));
 sky130_fd_sc_hd__nand3_4 _18560_ (.A(_08231_),
    .B(_08176_),
    .C(_08230_),
    .Y(_08236_));
 sky130_fd_sc_hd__o211ai_4 _18561_ (.A1(_07789_),
    .A2(_08175_),
    .B1(_08232_),
    .C1(_08233_),
    .Y(_08237_));
 sky130_fd_sc_hd__a21o_1 _18562_ (.A1(_08236_),
    .A2(_08237_),
    .B1(_08173_),
    .X(_08238_));
 sky130_fd_sc_hd__o211ai_4 _18563_ (.A1(_08168_),
    .A2(_08170_),
    .B1(_08236_),
    .C1(_08237_),
    .Y(_08240_));
 sky130_fd_sc_hd__a41oi_4 _18564_ (.A1(_07792_),
    .A2(_07813_),
    .A3(_08232_),
    .A4(_08233_),
    .B1(_08173_),
    .Y(_08241_));
 sky130_fd_sc_hd__nand4_4 _18565_ (.A(_08169_),
    .B(_08171_),
    .C(_08236_),
    .D(_08237_),
    .Y(_08242_));
 sky130_fd_sc_hd__a22o_2 _18566_ (.A1(_08169_),
    .A2(_08171_),
    .B1(_08236_),
    .B2(_08237_),
    .X(_08243_));
 sky130_fd_sc_hd__a22oi_4 _18567_ (.A1(_07820_),
    .A2(_07857_),
    .B1(_08238_),
    .B2(_08240_),
    .Y(_08244_));
 sky130_fd_sc_hd__nand3_4 _18568_ (.A(_08243_),
    .B(_08140_),
    .C(_08242_),
    .Y(_08245_));
 sky130_fd_sc_hd__a22oi_4 _18569_ (.A1(_07818_),
    .A2(_08139_),
    .B1(_08242_),
    .B2(_08243_),
    .Y(_08246_));
 sky130_fd_sc_hd__nand3_4 _18570_ (.A(_08142_),
    .B(_08238_),
    .C(_08240_),
    .Y(_08247_));
 sky130_fd_sc_hd__a32oi_4 _18571_ (.A1(_07866_),
    .A2(_07881_),
    .A3(_07882_),
    .B1(_07884_),
    .B2(_07897_),
    .Y(_08248_));
 sky130_fd_sc_hd__a32o_1 _18572_ (.A1(_07866_),
    .A2(_07881_),
    .A3(_07882_),
    .B1(_07884_),
    .B2(_07897_),
    .X(_08249_));
 sky130_fd_sc_hd__a22oi_4 _18573_ (.A1(_07842_),
    .A2(_07838_),
    .B1(_07821_),
    .B2(_07841_),
    .Y(_08251_));
 sky130_fd_sc_hd__a22o_1 _18574_ (.A1(_07842_),
    .A2(_07838_),
    .B1(_07821_),
    .B2(_07841_),
    .X(_08252_));
 sky130_fd_sc_hd__a32oi_4 _18575_ (.A1(net228),
    .A2(_02858_),
    .A3(net230),
    .B1(_02880_),
    .B2(net8),
    .Y(_08253_));
 sky130_fd_sc_hd__a32oi_4 _18576_ (.A1(net223),
    .A2(_01293_),
    .A3(net188),
    .B1(_01315_),
    .B2(net9),
    .Y(_08254_));
 sky130_fd_sc_hd__o2111ai_4 _18577_ (.A1(net231),
    .A2(_04557_),
    .B1(net36),
    .C1(net218),
    .D1(_03993_),
    .Y(_08255_));
 sky130_fd_sc_hd__or3_2 _18578_ (.A(net36),
    .B(_04080_),
    .C(_03993_),
    .X(_08256_));
 sky130_fd_sc_hd__o31a_1 _18579_ (.A1(net216),
    .A2(_12341_),
    .A3(_04554_),
    .B1(_08256_),
    .X(_08257_));
 sky130_fd_sc_hd__a21oi_1 _18580_ (.A1(_08255_),
    .A2(_08256_),
    .B1(_08254_),
    .Y(_08258_));
 sky130_fd_sc_hd__a21o_1 _18581_ (.A1(_08255_),
    .A2(_08256_),
    .B1(_08254_),
    .X(_08259_));
 sky130_fd_sc_hd__nand2_4 _18582_ (.A(_08254_),
    .B(_08257_),
    .Y(_08260_));
 sky130_fd_sc_hd__and3_2 _18583_ (.A(_08259_),
    .B(_08260_),
    .C(_08253_),
    .X(_08262_));
 sky130_fd_sc_hd__nand3_2 _18584_ (.A(_08259_),
    .B(_08260_),
    .C(_08253_),
    .Y(_08263_));
 sky130_fd_sc_hd__a21oi_4 _18585_ (.A1(_08259_),
    .A2(_08260_),
    .B1(_08253_),
    .Y(_08264_));
 sky130_fd_sc_hd__a21o_1 _18586_ (.A1(_08259_),
    .A2(_08260_),
    .B1(_08253_),
    .X(_08265_));
 sky130_fd_sc_hd__nand2_1 _18587_ (.A(_08263_),
    .B(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__o21ai_2 _18588_ (.A1(_07871_),
    .A2(_07874_),
    .B1(_07869_),
    .Y(_08267_));
 sky130_fd_sc_hd__o21ai_1 _18589_ (.A1(_07871_),
    .A2(_07874_),
    .B1(_07880_),
    .Y(_08268_));
 sky130_fd_sc_hd__o311a_1 _18590_ (.A1(net7),
    .A2(net249),
    .A3(_04787_),
    .B1(net252),
    .C1(net215),
    .X(_08269_));
 sky130_fd_sc_hd__and3_1 _18591_ (.A(_03993_),
    .B(net11),
    .C(net34),
    .X(_08270_));
 sky130_fd_sc_hd__a31o_1 _18592_ (.A1(net215),
    .A2(net252),
    .A3(net185),
    .B1(_08270_),
    .X(_08271_));
 sky130_fd_sc_hd__nand3_4 _18593_ (.A(net181),
    .B(net179),
    .C(net291),
    .Y(_08273_));
 sky130_fd_sc_hd__or3b_2 _18594_ (.A(net64),
    .B(_04135_),
    .C_N(net63),
    .X(_08274_));
 sky130_fd_sc_hd__and3_1 _18595_ (.A(_03971_),
    .B(net13),
    .C(net64),
    .X(_08275_));
 sky130_fd_sc_hd__o311a_1 _18596_ (.A1(net11),
    .A2(_04557_),
    .A3(net208),
    .B1(net289),
    .C1(net211),
    .X(_08276_));
 sky130_fd_sc_hd__a31oi_4 _18597_ (.A1(net211),
    .A2(net183),
    .A3(net289),
    .B1(_08275_),
    .Y(_08277_));
 sky130_fd_sc_hd__o211a_1 _18598_ (.A1(_04135_),
    .A2(_08283_),
    .B1(_08273_),
    .C1(_08277_),
    .X(_08278_));
 sky130_fd_sc_hd__o211ai_4 _18599_ (.A1(_04135_),
    .A2(_08283_),
    .B1(_08273_),
    .C1(_08277_),
    .Y(_08279_));
 sky130_fd_sc_hd__a21oi_4 _18600_ (.A1(_08273_),
    .A2(_08274_),
    .B1(_08277_),
    .Y(_08280_));
 sky130_fd_sc_hd__o2bb2ai_1 _18601_ (.A1_N(_08273_),
    .A2_N(_08274_),
    .B1(_08275_),
    .B2(_08276_),
    .Y(_08281_));
 sky130_fd_sc_hd__o21ai_2 _18602_ (.A1(_08269_),
    .A2(_08270_),
    .B1(_08279_),
    .Y(_08282_));
 sky130_fd_sc_hd__o211a_1 _18603_ (.A1(_08269_),
    .A2(_08270_),
    .B1(_08279_),
    .C1(_08281_),
    .X(_08284_));
 sky130_fd_sc_hd__o211ai_1 _18604_ (.A1(_08269_),
    .A2(_08270_),
    .B1(_08279_),
    .C1(_08281_),
    .Y(_08285_));
 sky130_fd_sc_hd__a21oi_1 _18605_ (.A1(_08279_),
    .A2(_08281_),
    .B1(_08271_),
    .Y(_08286_));
 sky130_fd_sc_hd__o21bai_2 _18606_ (.A1(_08278_),
    .A2(_08280_),
    .B1_N(_08271_),
    .Y(_08287_));
 sky130_fd_sc_hd__o211a_2 _18607_ (.A1(_08280_),
    .A2(_08282_),
    .B1(_08268_),
    .C1(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__o2111ai_4 _18608_ (.A1(_08282_),
    .A2(_08280_),
    .B1(_08267_),
    .C1(_07877_),
    .D1(_08287_),
    .Y(_08289_));
 sky130_fd_sc_hd__a21oi_2 _18609_ (.A1(_08285_),
    .A2(_08287_),
    .B1(_08268_),
    .Y(_08290_));
 sky130_fd_sc_hd__o2bb2ai_4 _18610_ (.A1_N(_07877_),
    .A2_N(_08267_),
    .B1(_08284_),
    .B2(_08286_),
    .Y(_08291_));
 sky130_fd_sc_hd__o21ai_4 _18611_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__o211ai_2 _18612_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08289_),
    .C1(_08291_),
    .Y(_08293_));
 sky130_fd_sc_hd__a21o_2 _18613_ (.A1(_08289_),
    .A2(_08291_),
    .B1(_08266_),
    .X(_08295_));
 sky130_fd_sc_hd__nand4_4 _18614_ (.A(_08263_),
    .B(_08265_),
    .C(_08289_),
    .D(_08291_),
    .Y(_08296_));
 sky130_fd_sc_hd__o22ai_4 _18615_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08288_),
    .B2(_08290_),
    .Y(_08297_));
 sky130_fd_sc_hd__o221a_1 _18616_ (.A1(_07843_),
    .A2(_07852_),
    .B1(_08288_),
    .B2(_08292_),
    .C1(_08295_),
    .X(_08298_));
 sky130_fd_sc_hd__o221ai_4 _18617_ (.A1(_07843_),
    .A2(_07852_),
    .B1(_08288_),
    .B2(_08292_),
    .C1(_08295_),
    .Y(_08299_));
 sky130_fd_sc_hd__nand3_4 _18618_ (.A(_08297_),
    .B(_08251_),
    .C(_08296_),
    .Y(_08300_));
 sky130_fd_sc_hd__a31oi_4 _18619_ (.A1(_08297_),
    .A2(_08251_),
    .A3(_08296_),
    .B1(_08249_),
    .Y(_08301_));
 sky130_fd_sc_hd__nand3_4 _18620_ (.A(_08299_),
    .B(_08300_),
    .C(_08248_),
    .Y(_08302_));
 sky130_fd_sc_hd__inv_2 _18621_ (.A(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__a21oi_2 _18622_ (.A1(_08299_),
    .A2(_08300_),
    .B1(_08248_),
    .Y(_08304_));
 sky130_fd_sc_hd__a21o_2 _18623_ (.A1(_08299_),
    .A2(_08300_),
    .B1(_08248_),
    .X(_08306_));
 sky130_fd_sc_hd__nand2_1 _18624_ (.A(_08302_),
    .B(_08306_),
    .Y(_08307_));
 sky130_fd_sc_hd__o211ai_4 _18625_ (.A1(_08303_),
    .A2(_08304_),
    .B1(_08245_),
    .C1(_08247_),
    .Y(_08308_));
 sky130_fd_sc_hd__o21bai_4 _18626_ (.A1(_08244_),
    .A2(_08246_),
    .B1_N(_08307_),
    .Y(_08309_));
 sky130_fd_sc_hd__o2bb2ai_2 _18627_ (.A1_N(_08245_),
    .A2_N(_08247_),
    .B1(_08303_),
    .B2(_08304_),
    .Y(_08310_));
 sky130_fd_sc_hd__nand3_1 _18628_ (.A(_08247_),
    .B(_08302_),
    .C(_08306_),
    .Y(_08311_));
 sky130_fd_sc_hd__nand4_2 _18629_ (.A(_08245_),
    .B(_08247_),
    .C(_08302_),
    .D(_08306_),
    .Y(_08312_));
 sky130_fd_sc_hd__and3_2 _18630_ (.A(_08137_),
    .B(_08310_),
    .C(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__nand3_4 _18631_ (.A(_08137_),
    .B(_08310_),
    .C(_08312_),
    .Y(_08314_));
 sky130_fd_sc_hd__and3_1 _18632_ (.A(_08138_),
    .B(_08308_),
    .C(_08309_),
    .X(_08315_));
 sky130_fd_sc_hd__o211ai_4 _18633_ (.A1(_07863_),
    .A2(_08135_),
    .B1(_08308_),
    .C1(_08309_),
    .Y(_08317_));
 sky130_fd_sc_hd__a31oi_4 _18634_ (.A1(_08138_),
    .A2(_08308_),
    .A3(_08309_),
    .B1(_08134_),
    .Y(_08318_));
 sky130_fd_sc_hd__o2111a_1 _18635_ (.A1(_08132_),
    .A2(_08127_),
    .B1(_08131_),
    .C1(_08314_),
    .D1(_08317_),
    .X(_08319_));
 sky130_fd_sc_hd__o2111ai_4 _18636_ (.A1(_08132_),
    .A2(_08127_),
    .B1(_08131_),
    .C1(_08314_),
    .D1(_08317_),
    .Y(_08320_));
 sky130_fd_sc_hd__a2bb2oi_1 _18637_ (.A1_N(_08129_),
    .A2_N(_08133_),
    .B1(_08314_),
    .B2(_08317_),
    .Y(_08321_));
 sky130_fd_sc_hd__a2bb2o_2 _18638_ (.A1_N(_08129_),
    .A2_N(_08133_),
    .B1(_08314_),
    .B2(_08317_),
    .X(_08322_));
 sky130_fd_sc_hd__a221oi_2 _18639_ (.A1(_07920_),
    .A2(_07925_),
    .B1(_08318_),
    .B2(_08314_),
    .C1(_08321_),
    .Y(_08323_));
 sky130_fd_sc_hd__nand3_2 _18640_ (.A(_08322_),
    .B(_08048_),
    .C(_08320_),
    .Y(_08324_));
 sky130_fd_sc_hd__a2bb2oi_4 _18641_ (.A1_N(_07917_),
    .A2_N(_08047_),
    .B1(_08320_),
    .B2(_08322_),
    .Y(_08325_));
 sky130_fd_sc_hd__o22ai_2 _18642_ (.A1(_07917_),
    .A2(_08047_),
    .B1(_08319_),
    .B2(_08321_),
    .Y(_08326_));
 sky130_fd_sc_hd__nand3_1 _18643_ (.A(_08046_),
    .B(_08324_),
    .C(_08326_),
    .Y(_08328_));
 sky130_fd_sc_hd__o22ai_2 _18644_ (.A1(_08044_),
    .A2(_08045_),
    .B1(_08323_),
    .B2(_08325_),
    .Y(_08329_));
 sky130_fd_sc_hd__o211a_1 _18645_ (.A1(_08044_),
    .A2(_08045_),
    .B1(_08324_),
    .C1(_08326_),
    .X(_08330_));
 sky130_fd_sc_hd__o2111ai_2 _18646_ (.A1(_08041_),
    .A2(_08038_),
    .B1(_08040_),
    .C1(_08324_),
    .D1(_08326_),
    .Y(_08331_));
 sky130_fd_sc_hd__o2bb2ai_1 _18647_ (.A1_N(_08040_),
    .A2_N(_08043_),
    .B1(_08323_),
    .B2(_08325_),
    .Y(_08332_));
 sky130_fd_sc_hd__nand2_1 _18648_ (.A(_07932_),
    .B(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__and3_1 _18649_ (.A(_07932_),
    .B(_08331_),
    .C(_08332_),
    .X(_08334_));
 sky130_fd_sc_hd__nand3_1 _18650_ (.A(_07932_),
    .B(_08331_),
    .C(_08332_),
    .Y(_08335_));
 sky130_fd_sc_hd__o211ai_4 _18651_ (.A1(_07929_),
    .A2(_07931_),
    .B1(_08328_),
    .C1(_08329_),
    .Y(_08336_));
 sky130_fd_sc_hd__and3_1 _18652_ (.A(_07304_),
    .B(_07315_),
    .C(_07666_),
    .X(_08337_));
 sky130_fd_sc_hd__a32o_1 _18653_ (.A1(_07657_),
    .A2(_07660_),
    .A3(_07662_),
    .B1(_07663_),
    .B2(_07667_),
    .X(_08339_));
 sky130_fd_sc_hd__o2111ai_2 _18654_ (.A1(_08330_),
    .A2(_08333_),
    .B1(_08336_),
    .C1(_07672_),
    .D1(_07666_),
    .Y(_08340_));
 sky130_fd_sc_hd__a22o_1 _18655_ (.A1(_07666_),
    .A2(_07672_),
    .B1(_08335_),
    .B2(_08336_),
    .X(_08341_));
 sky130_fd_sc_hd__o2bb2ai_2 _18656_ (.A1_N(_08335_),
    .A2_N(_08336_),
    .B1(_08337_),
    .B2(_07664_),
    .Y(_08342_));
 sky130_fd_sc_hd__nand2_2 _18657_ (.A(_08336_),
    .B(_08339_),
    .Y(_08343_));
 sky130_fd_sc_hd__o21ai_2 _18658_ (.A1(_08343_),
    .A2(_08334_),
    .B1(_08342_),
    .Y(_08344_));
 sky130_fd_sc_hd__nand3_1 _18659_ (.A(_07961_),
    .B(_08340_),
    .C(_08341_),
    .Y(_08345_));
 sky130_fd_sc_hd__o221a_1 _18660_ (.A1(_07941_),
    .A2(_07945_),
    .B1(_08334_),
    .B2(_08343_),
    .C1(_08342_),
    .X(_08346_));
 sky130_fd_sc_hd__o221ai_2 _18661_ (.A1(_07941_),
    .A2(_07945_),
    .B1(_08343_),
    .B2(_08334_),
    .C1(_08342_),
    .Y(_08347_));
 sky130_fd_sc_hd__a21oi_1 _18662_ (.A1(_08345_),
    .A2(_08347_),
    .B1(_07952_),
    .Y(_08348_));
 sky130_fd_sc_hd__a21oi_1 _18663_ (.A1(_08344_),
    .A2(_07961_),
    .B1(_07953_),
    .Y(_08350_));
 sky130_fd_sc_hd__and3_1 _18664_ (.A(_07952_),
    .B(_08345_),
    .C(_08347_),
    .X(_08351_));
 sky130_fd_sc_hd__o21ai_1 _18665_ (.A1(_07961_),
    .A2(_08344_),
    .B1(_08350_),
    .Y(_08352_));
 sky130_fd_sc_hd__a21oi_1 _18666_ (.A1(_08350_),
    .A2(_08347_),
    .B1(_08348_),
    .Y(_08353_));
 sky130_fd_sc_hd__a21oi_1 _18667_ (.A1(_07592_),
    .A2(_07595_),
    .B1(_07954_),
    .Y(_08354_));
 sky130_fd_sc_hd__a21boi_1 _18668_ (.A1(_07601_),
    .A2(_07957_),
    .B1_N(_07956_),
    .Y(_08355_));
 sky130_fd_sc_hd__or3_1 _18669_ (.A(_08348_),
    .B(_08351_),
    .C(_08355_),
    .X(_08356_));
 sky130_fd_sc_hd__xnor2_1 _18670_ (.A(_08353_),
    .B(_08355_),
    .Y(net88));
 sky130_fd_sc_hd__o21ai_2 _18671_ (.A1(_08330_),
    .A2(_08333_),
    .B1(_08343_),
    .Y(_08357_));
 sky130_fd_sc_hd__o2bb2a_1 _18672_ (.A1_N(_08336_),
    .A2_N(_08339_),
    .B1(_08330_),
    .B2(_08333_),
    .X(_08358_));
 sky130_fd_sc_hd__o21ba_1 _18673_ (.A1(_07963_),
    .A2(_08039_),
    .B1_N(_08038_),
    .X(_08360_));
 sky130_fd_sc_hd__inv_2 _18674_ (.A(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__a32oi_4 _18675_ (.A1(_08320_),
    .A2(_08322_),
    .A3(_08048_),
    .B1(_08043_),
    .B2(_08040_),
    .Y(_08362_));
 sky130_fd_sc_hd__a21oi_1 _18676_ (.A1(_08046_),
    .A2(_08324_),
    .B1(_08325_),
    .Y(_08363_));
 sky130_fd_sc_hd__a21boi_4 _18677_ (.A1(_08125_),
    .A2(_08128_),
    .B1_N(_08126_),
    .Y(_08364_));
 sky130_fd_sc_hd__nand2_1 _18678_ (.A(_08126_),
    .B(_08132_),
    .Y(_08365_));
 sky130_fd_sc_hd__o211ai_2 _18679_ (.A1(_04747_),
    .A2(net264),
    .B1(_06026_),
    .C1(_06486_),
    .Y(_08366_));
 sky130_fd_sc_hd__or3b_1 _18680_ (.A(_03916_),
    .B(net49),
    .C_N(net48),
    .X(_08367_));
 sky130_fd_sc_hd__or3b_2 _18681_ (.A(_03938_),
    .B(net48),
    .C_N(net47),
    .X(_08368_));
 sky130_fd_sc_hd__nand3_1 _18682_ (.A(_07242_),
    .B(net257),
    .C(net275),
    .Y(_08369_));
 sky130_fd_sc_hd__o2111a_1 _18683_ (.A1(_03916_),
    .A2(_06030_),
    .B1(_08366_),
    .C1(_08368_),
    .D1(_08369_),
    .X(_08371_));
 sky130_fd_sc_hd__o2111ai_1 _18684_ (.A1(_03916_),
    .A2(_06030_),
    .B1(_08366_),
    .C1(_08368_),
    .D1(_08369_),
    .Y(_08372_));
 sky130_fd_sc_hd__a22oi_2 _18685_ (.A1(_08366_),
    .A2(_08367_),
    .B1(_08368_),
    .B2(_08369_),
    .Y(_08373_));
 sky130_fd_sc_hd__a22o_1 _18686_ (.A1(_08366_),
    .A2(_08367_),
    .B1(_08368_),
    .B2(_08369_),
    .X(_08374_));
 sky130_fd_sc_hd__a32o_1 _18687_ (.A1(_05841_),
    .A2(net265),
    .A3(net273),
    .B1(_06326_),
    .B2(net29),
    .X(_08375_));
 sky130_fd_sc_hd__o21bai_2 _18688_ (.A1(_08371_),
    .A2(_08373_),
    .B1_N(_08375_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand3_1 _18689_ (.A(_08372_),
    .B(_08374_),
    .C(_08375_),
    .Y(_08377_));
 sky130_fd_sc_hd__o21ai_2 _18690_ (.A1(_08103_),
    .A2(_08111_),
    .B1(_08110_),
    .Y(_08378_));
 sky130_fd_sc_hd__a21o_1 _18691_ (.A1(_08376_),
    .A2(_08377_),
    .B1(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__nand3_4 _18692_ (.A(_08378_),
    .B(_08377_),
    .C(_08376_),
    .Y(_08380_));
 sky130_fd_sc_hd__o221a_1 _18693_ (.A1(_05020_),
    .A2(_06864_),
    .B1(_06866_),
    .B2(_03616_),
    .C1(_07980_),
    .X(_08382_));
 sky130_fd_sc_hd__nand2_1 _18694_ (.A(_07980_),
    .B(_07972_),
    .Y(_08383_));
 sky130_fd_sc_hd__o2bb2ai_1 _18695_ (.A1_N(_08379_),
    .A2_N(_08380_),
    .B1(_08382_),
    .B2(_07981_),
    .Y(_08384_));
 sky130_fd_sc_hd__nand4_4 _18696_ (.A(_07982_),
    .B(_08379_),
    .C(_08380_),
    .D(_08383_),
    .Y(_08385_));
 sky130_fd_sc_hd__a21o_1 _18697_ (.A1(_08100_),
    .A2(_08114_),
    .B1(_08101_),
    .X(_08386_));
 sky130_fd_sc_hd__a21o_1 _18698_ (.A1(_08384_),
    .A2(_08385_),
    .B1(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__nand3_1 _18699_ (.A(_08386_),
    .B(_08385_),
    .C(_08384_),
    .Y(_08388_));
 sky130_fd_sc_hd__a21bo_1 _18700_ (.A1(_07970_),
    .A2(_07989_),
    .B1_N(_07988_),
    .X(_08389_));
 sky130_fd_sc_hd__a21o_1 _18701_ (.A1(_08387_),
    .A2(_08388_),
    .B1(_08389_),
    .X(_08390_));
 sky130_fd_sc_hd__nand3_1 _18702_ (.A(_08387_),
    .B(_08388_),
    .C(_08389_),
    .Y(_08391_));
 sky130_fd_sc_hd__nand2_1 _18703_ (.A(_07996_),
    .B(_07997_),
    .Y(_08393_));
 sky130_fd_sc_hd__a21oi_1 _18704_ (.A1(_08390_),
    .A2(_08391_),
    .B1(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__a21o_1 _18705_ (.A1(_08390_),
    .A2(_08391_),
    .B1(_08393_),
    .X(_08395_));
 sky130_fd_sc_hd__and3_1 _18706_ (.A(_08390_),
    .B(_08391_),
    .C(_08393_),
    .X(_08396_));
 sky130_fd_sc_hd__nand3_1 _18707_ (.A(_08390_),
    .B(_08391_),
    .C(_08393_),
    .Y(_08397_));
 sky130_fd_sc_hd__a22oi_1 _18708_ (.A1(_04539_),
    .A2(_08005_),
    .B1(_08006_),
    .B2(net12),
    .Y(_08398_));
 sky130_fd_sc_hd__a22o_1 _18709_ (.A1(_04539_),
    .A2(_08005_),
    .B1(_08006_),
    .B2(net12),
    .X(_08399_));
 sky130_fd_sc_hd__and3_1 _18710_ (.A(_07642_),
    .B(_04452_),
    .C(net318),
    .X(_08400_));
 sky130_fd_sc_hd__a21oi_1 _18711_ (.A1(net23),
    .A2(_07643_),
    .B1(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__a21oi_1 _18712_ (.A1(_08012_),
    .A2(_08019_),
    .B1(_08017_),
    .Y(_08402_));
 sky130_fd_sc_hd__a32o_1 _18713_ (.A1(net313),
    .A2(_04747_),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net26),
    .X(_08404_));
 sky130_fd_sc_hd__or3b_1 _18714_ (.A(_03616_),
    .B(net52),
    .C_N(net51),
    .X(_08405_));
 sky130_fd_sc_hd__nand3_2 _18715_ (.A(net266),
    .B(net301),
    .C(_07223_),
    .Y(_08406_));
 sky130_fd_sc_hd__or3_2 _18716_ (.A(net51),
    .B(_04190_),
    .C(_03725_),
    .X(_08407_));
 sky130_fd_sc_hd__nand3_2 _18717_ (.A(_05414_),
    .B(_05446_),
    .C(_06863_),
    .Y(_08408_));
 sky130_fd_sc_hd__a22oi_1 _18718_ (.A1(_08405_),
    .A2(_08406_),
    .B1(_08407_),
    .B2(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__a22o_1 _18719_ (.A1(_08405_),
    .A2(_08406_),
    .B1(_08407_),
    .B2(_08408_),
    .X(_08410_));
 sky130_fd_sc_hd__o2111ai_4 _18720_ (.A1(_03616_),
    .A2(_07226_),
    .B1(_08406_),
    .C1(_08407_),
    .D1(_08408_),
    .Y(_08411_));
 sky130_fd_sc_hd__nand3_1 _18721_ (.A(_08404_),
    .B(_08410_),
    .C(_08411_),
    .Y(_08412_));
 sky130_fd_sc_hd__a21o_1 _18722_ (.A1(_08410_),
    .A2(_08411_),
    .B1(_08404_),
    .X(_08413_));
 sky130_fd_sc_hd__a21bo_1 _18723_ (.A1(_08410_),
    .A2(_08411_),
    .B1_N(_08404_),
    .X(_08415_));
 sky130_fd_sc_hd__nand3b_1 _18724_ (.A_N(_08404_),
    .B(_08410_),
    .C(_08411_),
    .Y(_08416_));
 sky130_fd_sc_hd__nand3_2 _18725_ (.A(_08415_),
    .B(_08416_),
    .C(_08402_),
    .Y(_08417_));
 sky130_fd_sc_hd__nand3b_1 _18726_ (.A_N(_08402_),
    .B(_08412_),
    .C(_08413_),
    .Y(_08418_));
 sky130_fd_sc_hd__and3b_1 _18727_ (.A_N(_08401_),
    .B(_08417_),
    .C(_08418_),
    .X(_08419_));
 sky130_fd_sc_hd__a221oi_2 _18728_ (.A1(net23),
    .A2(_07643_),
    .B1(_08417_),
    .B2(_08418_),
    .C1(_08400_),
    .Y(_08420_));
 sky130_fd_sc_hd__a211oi_2 _18729_ (.A1(_08023_),
    .A2(_08027_),
    .B1(_08419_),
    .C1(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__o211ai_2 _18730_ (.A1(_08419_),
    .A2(_08420_),
    .B1(_08023_),
    .C1(_08027_),
    .Y(_08422_));
 sky130_fd_sc_hd__inv_2 _18731_ (.A(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__o21ai_1 _18732_ (.A1(_08421_),
    .A2(_08423_),
    .B1(_08399_),
    .Y(_08424_));
 sky130_fd_sc_hd__nand3b_1 _18733_ (.A_N(_08421_),
    .B(_08422_),
    .C(_08398_),
    .Y(_08426_));
 sky130_fd_sc_hd__nand2_1 _18734_ (.A(_08424_),
    .B(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__o211a_1 _18735_ (.A1(_08394_),
    .A2(_08396_),
    .B1(_08424_),
    .C1(_08426_),
    .X(_08428_));
 sky130_fd_sc_hd__o21bai_2 _18736_ (.A1(_08394_),
    .A2(_08396_),
    .B1_N(_08427_),
    .Y(_08429_));
 sky130_fd_sc_hd__nand3_2 _18737_ (.A(_08395_),
    .B(_08397_),
    .C(_08427_),
    .Y(_08430_));
 sky130_fd_sc_hd__nand2_2 _18738_ (.A(_08429_),
    .B(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__a21oi_2 _18739_ (.A1(_08429_),
    .A2(_08430_),
    .B1(_08365_),
    .Y(_08432_));
 sky130_fd_sc_hd__a221o_1 _18740_ (.A1(_08125_),
    .A2(_08128_),
    .B1(_08429_),
    .B2(_08430_),
    .C1(_08127_),
    .X(_08433_));
 sky130_fd_sc_hd__a31o_1 _18741_ (.A1(_08395_),
    .A2(_08397_),
    .A3(_08427_),
    .B1(_08364_),
    .X(_08434_));
 sky130_fd_sc_hd__and3_2 _18742_ (.A(_08365_),
    .B(_08429_),
    .C(_08430_),
    .X(_08435_));
 sky130_fd_sc_hd__and3_2 _18743_ (.A(_08004_),
    .B(_08030_),
    .C(_08032_),
    .X(_08437_));
 sky130_fd_sc_hd__or2_1 _18744_ (.A(_08002_),
    .B(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__o22a_1 _18745_ (.A1(_08432_),
    .A2(_08435_),
    .B1(_08437_),
    .B2(_08002_),
    .X(_08439_));
 sky130_fd_sc_hd__o21ai_1 _18746_ (.A1(_08432_),
    .A2(_08435_),
    .B1(_08438_),
    .Y(_08440_));
 sky130_fd_sc_hd__a21oi_2 _18747_ (.A1(_08431_),
    .A2(_08364_),
    .B1(_08438_),
    .Y(_08441_));
 sky130_fd_sc_hd__a31o_1 _18748_ (.A1(_08126_),
    .A2(_08132_),
    .A3(_08431_),
    .B1(_08438_),
    .X(_08442_));
 sky130_fd_sc_hd__o21a_1 _18749_ (.A1(_08364_),
    .A2(_08431_),
    .B1(_08441_),
    .X(_08443_));
 sky130_fd_sc_hd__o221a_1 _18750_ (.A1(_08428_),
    .A2(_08434_),
    .B1(_08437_),
    .B2(_08002_),
    .C1(_08433_),
    .X(_08444_));
 sky130_fd_sc_hd__o221ai_4 _18751_ (.A1(_08428_),
    .A2(_08434_),
    .B1(_08437_),
    .B2(_08002_),
    .C1(_08433_),
    .Y(_08445_));
 sky130_fd_sc_hd__o21ba_1 _18752_ (.A1(_08432_),
    .A2(_08435_),
    .B1_N(_08438_),
    .X(_08446_));
 sky130_fd_sc_hd__o21bai_1 _18753_ (.A1(_08432_),
    .A2(_08435_),
    .B1_N(_08438_),
    .Y(_08448_));
 sky130_fd_sc_hd__o21ai_1 _18754_ (.A1(_08435_),
    .A2(_08442_),
    .B1(_08440_),
    .Y(_08449_));
 sky130_fd_sc_hd__o21a_1 _18755_ (.A1(_08129_),
    .A2(_08133_),
    .B1(_08314_),
    .X(_08450_));
 sky130_fd_sc_hd__a32o_1 _18756_ (.A1(_08138_),
    .A2(_08308_),
    .A3(_08309_),
    .B1(_08314_),
    .B2(_08134_),
    .X(_08451_));
 sky130_fd_sc_hd__o21ai_2 _18757_ (.A1(_08116_),
    .A2(_08118_),
    .B1(_08080_),
    .Y(_08452_));
 sky130_fd_sc_hd__nand2_1 _18758_ (.A(_08080_),
    .B(_08124_),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_1 _18759_ (.A(_08081_),
    .B(_08452_),
    .Y(_08454_));
 sky130_fd_sc_hd__a32oi_4 _18760_ (.A1(_08252_),
    .A2(_08293_),
    .A3(_08295_),
    .B1(_08300_),
    .B2(_08248_),
    .Y(_08455_));
 sky130_fd_sc_hd__o21a_2 _18761_ (.A1(_08058_),
    .A2(_08062_),
    .B1(_08069_),
    .X(_08456_));
 sky130_fd_sc_hd__o21ai_2 _18762_ (.A1(_08254_),
    .A2(_08257_),
    .B1(_08253_),
    .Y(_08457_));
 sky130_fd_sc_hd__a31oi_2 _18763_ (.A1(_08254_),
    .A2(_08255_),
    .A3(_08256_),
    .B1(_08253_),
    .Y(_08459_));
 sky130_fd_sc_hd__a32o_1 _18764_ (.A1(_03952_),
    .A2(net231),
    .A3(net281),
    .B1(_04217_),
    .B2(net7),
    .X(_08460_));
 sky130_fd_sc_hd__nand3_2 _18765_ (.A(net223),
    .B(_02858_),
    .C(net188),
    .Y(_08461_));
 sky130_fd_sc_hd__or3b_2 _18766_ (.A(net38),
    .B(_04069_),
    .C_N(net37),
    .X(_08462_));
 sky130_fd_sc_hd__nor2_1 _18767_ (.A(_04059_),
    .B(_03737_),
    .Y(_08463_));
 sky130_fd_sc_hd__a31oi_4 _18768_ (.A1(net228),
    .A2(net285),
    .A3(net230),
    .B1(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__a21oi_4 _18769_ (.A1(_08461_),
    .A2(_08462_),
    .B1(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__a21o_1 _18770_ (.A1(_08461_),
    .A2(_08462_),
    .B1(_08464_),
    .X(_08466_));
 sky130_fd_sc_hd__o211a_1 _18771_ (.A1(_04069_),
    .A2(_02891_),
    .B1(_08461_),
    .C1(_08464_),
    .X(_08467_));
 sky130_fd_sc_hd__o221ai_4 _18772_ (.A1(_04069_),
    .A2(_02891_),
    .B1(net187),
    .B2(_02869_),
    .C1(_08464_),
    .Y(_08468_));
 sky130_fd_sc_hd__o21bai_4 _18773_ (.A1(_08465_),
    .A2(_08467_),
    .B1_N(_08460_),
    .Y(_08470_));
 sky130_fd_sc_hd__and3_1 _18774_ (.A(_08460_),
    .B(_08466_),
    .C(_08468_),
    .X(_08471_));
 sky130_fd_sc_hd__nand3_2 _18775_ (.A(_08460_),
    .B(_08466_),
    .C(_08468_),
    .Y(_08472_));
 sky130_fd_sc_hd__o211a_1 _18776_ (.A1(_08258_),
    .A2(_08459_),
    .B1(_08470_),
    .C1(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__o211ai_2 _18777_ (.A1(_08258_),
    .A2(_08459_),
    .B1(_08470_),
    .C1(_08472_),
    .Y(_08474_));
 sky130_fd_sc_hd__a22oi_4 _18778_ (.A1(_08260_),
    .A2(_08457_),
    .B1(_08470_),
    .B2(_08472_),
    .Y(_08475_));
 sky130_fd_sc_hd__a22o_1 _18779_ (.A1(_08260_),
    .A2(_08457_),
    .B1(_08470_),
    .B2(_08472_),
    .X(_08476_));
 sky130_fd_sc_hd__o21ai_4 _18780_ (.A1(_08473_),
    .A2(_08475_),
    .B1(_08456_),
    .Y(_08477_));
 sky130_fd_sc_hd__nand3b_2 _18781_ (.A_N(_08456_),
    .B(_08474_),
    .C(_08476_),
    .Y(_08478_));
 sky130_fd_sc_hd__o21ai_2 _18782_ (.A1(_07734_),
    .A2(_08073_),
    .B1(_08072_),
    .Y(_08479_));
 sky130_fd_sc_hd__a21oi_2 _18783_ (.A1(_08477_),
    .A2(_08478_),
    .B1(_08479_),
    .Y(_08481_));
 sky130_fd_sc_hd__a21o_1 _18784_ (.A1(_08477_),
    .A2(_08478_),
    .B1(_08479_),
    .X(_08482_));
 sky130_fd_sc_hd__o311a_1 _18785_ (.A1(_07727_),
    .A2(_07733_),
    .A3(_08071_),
    .B1(_08074_),
    .C1(_08477_),
    .X(_08483_));
 sky130_fd_sc_hd__nand2_1 _18786_ (.A(_08477_),
    .B(_08479_),
    .Y(_08484_));
 sky130_fd_sc_hd__o21ai_2 _18787_ (.A1(_08094_),
    .A2(_08090_),
    .B1(_08089_),
    .Y(_08485_));
 sky130_fd_sc_hd__o22a_1 _18788_ (.A1(_13021_),
    .A2(_04896_),
    .B1(_04898_),
    .B2(_04004_),
    .X(_08486_));
 sky130_fd_sc_hd__a32o_1 _18789_ (.A1(net234),
    .A2(net251),
    .A3(net243),
    .B1(_04897_),
    .B2(net4),
    .X(_08487_));
 sky130_fd_sc_hd__o211ai_4 _18790_ (.A1(net253),
    .A2(_02442_),
    .B1(net280),
    .C1(_02421_),
    .Y(_08488_));
 sky130_fd_sc_hd__or3b_1 _18791_ (.A(_04026_),
    .B(net41),
    .C_N(net40),
    .X(_08489_));
 sky130_fd_sc_hd__or3b_2 _18792_ (.A(_04015_),
    .B(net42),
    .C_N(net41),
    .X(_08490_));
 sky130_fd_sc_hd__o211ai_4 _18793_ (.A1(net253),
    .A2(_00646_),
    .B1(net279),
    .C1(_00625_),
    .Y(_08492_));
 sky130_fd_sc_hd__a22oi_1 _18794_ (.A1(_08488_),
    .A2(_08489_),
    .B1(_08490_),
    .B2(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__a22o_2 _18795_ (.A1(_08488_),
    .A2(_08489_),
    .B1(_08490_),
    .B2(_08492_),
    .X(_08494_));
 sky130_fd_sc_hd__o2111a_1 _18796_ (.A1(_04026_),
    .A2(_04270_),
    .B1(_08488_),
    .C1(_08490_),
    .D1(_08492_),
    .X(_08495_));
 sky130_fd_sc_hd__o2111ai_4 _18797_ (.A1(_04026_),
    .A2(_04270_),
    .B1(_08488_),
    .C1(_08490_),
    .D1(_08492_),
    .Y(_08496_));
 sky130_fd_sc_hd__a21oi_2 _18798_ (.A1(_08494_),
    .A2(_08496_),
    .B1(_08487_),
    .Y(_08497_));
 sky130_fd_sc_hd__nand3_1 _18799_ (.A(_08494_),
    .B(_08496_),
    .C(_08486_),
    .Y(_08498_));
 sky130_fd_sc_hd__o21ai_1 _18800_ (.A1(_08493_),
    .A2(_08495_),
    .B1(_08487_),
    .Y(_08499_));
 sky130_fd_sc_hd__nand3_2 _18801_ (.A(_08499_),
    .B(_08485_),
    .C(_08498_),
    .Y(_08500_));
 sky130_fd_sc_hd__a31o_1 _18802_ (.A1(_08487_),
    .A2(_08494_),
    .A3(_08496_),
    .B1(_08485_),
    .X(_08501_));
 sky130_fd_sc_hd__a21o_1 _18803_ (.A1(_08498_),
    .A2(_08499_),
    .B1(_08485_),
    .X(_08503_));
 sky130_fd_sc_hd__a32o_1 _18804_ (.A1(net256),
    .A2(_08700_),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net32),
    .X(_08504_));
 sky130_fd_sc_hd__a31o_1 _18805_ (.A1(net309),
    .A2(net295),
    .A3(net290),
    .B1(_05226_),
    .X(_08505_));
 sky130_fd_sc_hd__o32a_4 _18806_ (.A1(_03960_),
    .A2(_04124_),
    .A3(net46),
    .B1(_09687_),
    .B2(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__or3_1 _18807_ (.A(net45),
    .B(_04102_),
    .C(_03982_),
    .X(_08507_));
 sky130_fd_sc_hd__o2111ai_4 _18808_ (.A1(net260),
    .A2(_11387_),
    .B1(net45),
    .C1(_11354_),
    .D1(_04102_),
    .Y(_08508_));
 sky130_fd_sc_hd__a21oi_1 _18809_ (.A1(_08507_),
    .A2(_08508_),
    .B1(_08506_),
    .Y(_08509_));
 sky130_fd_sc_hd__a21o_1 _18810_ (.A1(_08507_),
    .A2(_08508_),
    .B1(_08506_),
    .X(_08510_));
 sky130_fd_sc_hd__o311a_1 _18811_ (.A1(_03982_),
    .A2(_04102_),
    .A3(net45),
    .B1(_08508_),
    .C1(_08506_),
    .X(_08511_));
 sky130_fd_sc_hd__o221ai_2 _18812_ (.A1(_11453_),
    .A2(_04986_),
    .B1(_04989_),
    .B2(_03982_),
    .C1(_08506_),
    .Y(_08512_));
 sky130_fd_sc_hd__o21ai_1 _18813_ (.A1(_08509_),
    .A2(_08511_),
    .B1(_08504_),
    .Y(_08514_));
 sky130_fd_sc_hd__nand3b_1 _18814_ (.A_N(_08504_),
    .B(_08510_),
    .C(_08512_),
    .Y(_08515_));
 sky130_fd_sc_hd__nand2_1 _18815_ (.A(_08514_),
    .B(_08515_),
    .Y(_08516_));
 sky130_fd_sc_hd__o211ai_2 _18816_ (.A1(_08497_),
    .A2(_08501_),
    .B1(_08516_),
    .C1(_08500_),
    .Y(_08517_));
 sky130_fd_sc_hd__a21o_1 _18817_ (.A1(_08500_),
    .A2(_08503_),
    .B1(_08516_),
    .X(_08518_));
 sky130_fd_sc_hd__nand2_1 _18818_ (.A(_08517_),
    .B(_08518_),
    .Y(_08519_));
 sky130_fd_sc_hd__nand3_2 _18819_ (.A(_08482_),
    .B(_08484_),
    .C(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__o21bai_2 _18820_ (.A1(_08481_),
    .A2(_08483_),
    .B1_N(_08519_),
    .Y(_08521_));
 sky130_fd_sc_hd__o21ai_2 _18821_ (.A1(_08481_),
    .A2(_08483_),
    .B1(_08519_),
    .Y(_08522_));
 sky130_fd_sc_hd__nand4_2 _18822_ (.A(_08482_),
    .B(_08484_),
    .C(_08517_),
    .D(_08518_),
    .Y(_08523_));
 sky130_fd_sc_hd__o211ai_4 _18823_ (.A1(_08298_),
    .A2(_08301_),
    .B1(_08522_),
    .C1(_08523_),
    .Y(_08525_));
 sky130_fd_sc_hd__nand3_4 _18824_ (.A(_08521_),
    .B(_08455_),
    .C(_08520_),
    .Y(_08526_));
 sky130_fd_sc_hd__a31oi_1 _18825_ (.A1(_08521_),
    .A2(_08455_),
    .A3(_08520_),
    .B1(_08454_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand2_1 _18826_ (.A(_08527_),
    .B(_08525_),
    .Y(_08528_));
 sky130_fd_sc_hd__a22oi_1 _18827_ (.A1(_08081_),
    .A2(_08452_),
    .B1(_08525_),
    .B2(_08526_),
    .Y(_08529_));
 sky130_fd_sc_hd__a22o_1 _18828_ (.A1(_08081_),
    .A2(_08452_),
    .B1(_08525_),
    .B2(_08526_),
    .X(_08530_));
 sky130_fd_sc_hd__and4b_1 _18829_ (.A_N(_08455_),
    .B(_08522_),
    .C(_08523_),
    .D(_08453_),
    .X(_08531_));
 sky130_fd_sc_hd__a21oi_1 _18830_ (.A1(_08081_),
    .A2(_08452_),
    .B1(_08526_),
    .Y(_08532_));
 sky130_fd_sc_hd__nand2_2 _18831_ (.A(_08454_),
    .B(_08525_),
    .Y(_08533_));
 sky130_fd_sc_hd__a21oi_1 _18832_ (.A1(_08526_),
    .A2(_08533_),
    .B1(_08532_),
    .Y(_08534_));
 sky130_fd_sc_hd__a21oi_1 _18833_ (.A1(_08525_),
    .A2(_08527_),
    .B1(_08529_),
    .Y(_08536_));
 sky130_fd_sc_hd__a31o_1 _18834_ (.A1(_08453_),
    .A2(_08525_),
    .A3(_08526_),
    .B1(_08529_),
    .X(_08537_));
 sky130_fd_sc_hd__a32oi_4 _18835_ (.A1(_08243_),
    .A2(_08140_),
    .A3(_08242_),
    .B1(_08302_),
    .B2(_08306_),
    .Y(_08538_));
 sky130_fd_sc_hd__a31o_1 _18836_ (.A1(_08247_),
    .A2(_08302_),
    .A3(_08306_),
    .B1(_08244_),
    .X(_08539_));
 sky130_fd_sc_hd__a2bb2oi_2 _18837_ (.A1_N(_08158_),
    .A2_N(_08162_),
    .B1(_08167_),
    .B2(_08165_),
    .Y(_08540_));
 sky130_fd_sc_hd__o2bb2ai_2 _18838_ (.A1_N(_08167_),
    .A2_N(_08165_),
    .B1(_08162_),
    .B2(_08158_),
    .Y(_08541_));
 sky130_fd_sc_hd__a21oi_2 _18839_ (.A1(_08271_),
    .A2(_08279_),
    .B1(_08280_),
    .Y(_08542_));
 sky130_fd_sc_hd__a21o_1 _18840_ (.A1(_08271_),
    .A2(_08279_),
    .B1(_08280_),
    .X(_08543_));
 sky130_fd_sc_hd__and3_1 _18841_ (.A(_03971_),
    .B(net14),
    .C(net64),
    .X(_08544_));
 sky130_fd_sc_hd__a31oi_2 _18842_ (.A1(net181),
    .A2(net179),
    .A3(net289),
    .B1(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__a31o_2 _18843_ (.A1(net181),
    .A2(net179),
    .A3(net289),
    .B1(_08544_),
    .X(_08547_));
 sky130_fd_sc_hd__nor2_1 _18844_ (.A(_04146_),
    .B(_08283_),
    .Y(_08548_));
 sky130_fd_sc_hd__a31oi_4 _18845_ (.A1(_05549_),
    .A2(net177),
    .A3(net291),
    .B1(_08548_),
    .Y(_08549_));
 sky130_fd_sc_hd__a31o_1 _18846_ (.A1(_05549_),
    .A2(net177),
    .A3(net291),
    .B1(_08548_),
    .X(_08550_));
 sky130_fd_sc_hd__a221oi_2 _18847_ (.A1(_03957_),
    .A2(_05926_),
    .B1(net177),
    .B2(net16),
    .C1(_07669_),
    .Y(_08551_));
 sky130_fd_sc_hd__nor2_1 _18848_ (.A(_04157_),
    .B(_07691_),
    .Y(_08552_));
 sky130_fd_sc_hd__o32a_1 _18849_ (.A1(_07669_),
    .A2(net205),
    .A3(_05932_),
    .B1(_07691_),
    .B2(_04157_),
    .X(_08553_));
 sky130_fd_sc_hd__o21ai_4 _18850_ (.A1(_08551_),
    .A2(_08552_),
    .B1(_08550_),
    .Y(_08554_));
 sky130_fd_sc_hd__o221a_2 _18851_ (.A1(_04157_),
    .A2(_07691_),
    .B1(net155),
    .B2(_07669_),
    .C1(_08549_),
    .X(_08555_));
 sky130_fd_sc_hd__o221ai_4 _18852_ (.A1(_04157_),
    .A2(_07691_),
    .B1(net155),
    .B2(_07669_),
    .C1(_08549_),
    .Y(_08556_));
 sky130_fd_sc_hd__a21oi_4 _18853_ (.A1(_08554_),
    .A2(_08556_),
    .B1(_08547_),
    .Y(_08558_));
 sky130_fd_sc_hd__a21o_1 _18854_ (.A1(_08554_),
    .A2(_08556_),
    .B1(_08547_),
    .X(_08559_));
 sky130_fd_sc_hd__o21ai_2 _18855_ (.A1(_08549_),
    .A2(_08553_),
    .B1(_08547_),
    .Y(_08560_));
 sky130_fd_sc_hd__nand3_1 _18856_ (.A(_08554_),
    .B(_08556_),
    .C(_08545_),
    .Y(_08561_));
 sky130_fd_sc_hd__a21o_1 _18857_ (.A1(_08554_),
    .A2(_08556_),
    .B1(_08545_),
    .X(_08562_));
 sky130_fd_sc_hd__o21ai_4 _18858_ (.A1(_08555_),
    .A2(_08560_),
    .B1(_08543_),
    .Y(_08563_));
 sky130_fd_sc_hd__o211ai_2 _18859_ (.A1(_08560_),
    .A2(_08555_),
    .B1(_08543_),
    .C1(_08559_),
    .Y(_08564_));
 sky130_fd_sc_hd__and3_1 _18860_ (.A(_08562_),
    .B(_08542_),
    .C(_08561_),
    .X(_08565_));
 sky130_fd_sc_hd__nand3_4 _18861_ (.A(_08562_),
    .B(_08542_),
    .C(_08561_),
    .Y(_08566_));
 sky130_fd_sc_hd__o32a_1 _18862_ (.A1(net216),
    .A2(_01304_),
    .A3(_04554_),
    .B1(_01326_),
    .B2(_04080_),
    .X(_08567_));
 sky130_fd_sc_hd__a32o_1 _18863_ (.A1(net218),
    .A2(_04559_),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net10),
    .X(_08569_));
 sky130_fd_sc_hd__o211ai_4 _18864_ (.A1(net231),
    .A2(_04787_),
    .B1(_12330_),
    .C1(net215),
    .Y(_08570_));
 sky130_fd_sc_hd__or3_2 _18865_ (.A(net36),
    .B(_04091_),
    .C(_03993_),
    .X(_08571_));
 sky130_fd_sc_hd__or3_2 _18866_ (.A(net35),
    .B(_04113_),
    .C(_03971_),
    .X(_08572_));
 sky130_fd_sc_hd__o211ai_4 _18867_ (.A1(_04787_),
    .A2(net208),
    .B1(net252),
    .C1(net211),
    .Y(_08573_));
 sky130_fd_sc_hd__a22oi_4 _18868_ (.A1(_08570_),
    .A2(_08571_),
    .B1(_08572_),
    .B2(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__and4_1 _18869_ (.A(_08570_),
    .B(_08571_),
    .C(_08572_),
    .D(_08573_),
    .X(_08575_));
 sky130_fd_sc_hd__nand4_2 _18870_ (.A(_08570_),
    .B(_08571_),
    .C(_08572_),
    .D(_08573_),
    .Y(_08576_));
 sky130_fd_sc_hd__a21oi_4 _18871_ (.A1(_08569_),
    .A2(_08576_),
    .B1(_08574_),
    .Y(_08577_));
 sky130_fd_sc_hd__nor2_1 _18872_ (.A(_08574_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__o21a_1 _18873_ (.A1(_08574_),
    .A2(_08575_),
    .B1(_08569_),
    .X(_08580_));
 sky130_fd_sc_hd__nor3_1 _18874_ (.A(_08569_),
    .B(_08574_),
    .C(_08575_),
    .Y(_08581_));
 sky130_fd_sc_hd__o21a_1 _18875_ (.A1(_08574_),
    .A2(_08575_),
    .B1(_08567_),
    .X(_08582_));
 sky130_fd_sc_hd__o21ai_1 _18876_ (.A1(_08574_),
    .A2(_08575_),
    .B1(_08567_),
    .Y(_08583_));
 sky130_fd_sc_hd__o21a_1 _18877_ (.A1(_08574_),
    .A2(_08577_),
    .B1(_08583_),
    .X(_08584_));
 sky130_fd_sc_hd__o2bb2ai_2 _18878_ (.A1_N(_08564_),
    .A2_N(_08566_),
    .B1(_08580_),
    .B2(_08581_),
    .Y(_08585_));
 sky130_fd_sc_hd__o221ai_4 _18879_ (.A1(_08558_),
    .A2(_08563_),
    .B1(_08578_),
    .B2(_08582_),
    .C1(_08566_),
    .Y(_08586_));
 sky130_fd_sc_hd__o2bb2ai_2 _18880_ (.A1_N(_08564_),
    .A2_N(_08566_),
    .B1(_08578_),
    .B2(_08582_),
    .Y(_08587_));
 sky130_fd_sc_hd__o21ai_2 _18881_ (.A1(_08558_),
    .A2(_08563_),
    .B1(_08584_),
    .Y(_08588_));
 sky130_fd_sc_hd__nand4_2 _18882_ (.A(_08164_),
    .B(_08171_),
    .C(_08585_),
    .D(_08586_),
    .Y(_08589_));
 sky130_fd_sc_hd__o211a_2 _18883_ (.A1(_08588_),
    .A2(_08565_),
    .B1(_08541_),
    .C1(_08587_),
    .X(_08591_));
 sky130_fd_sc_hd__o211ai_4 _18884_ (.A1(_08588_),
    .A2(_08565_),
    .B1(_08541_),
    .C1(_08587_),
    .Y(_08592_));
 sky130_fd_sc_hd__a31o_1 _18885_ (.A1(_08263_),
    .A2(_08265_),
    .A3(_08289_),
    .B1(_08290_),
    .X(_08593_));
 sky130_fd_sc_hd__a31oi_4 _18886_ (.A1(_08585_),
    .A2(_08586_),
    .A3(_08540_),
    .B1(_08593_),
    .Y(_08594_));
 sky130_fd_sc_hd__a31o_2 _18887_ (.A1(_08585_),
    .A2(_08586_),
    .A3(_08540_),
    .B1(_08593_),
    .X(_08595_));
 sky130_fd_sc_hd__nand2_2 _18888_ (.A(_08594_),
    .B(_08592_),
    .Y(_08596_));
 sky130_fd_sc_hd__a21bo_2 _18889_ (.A1(_08589_),
    .A2(_08592_),
    .B1_N(_08593_),
    .X(_08597_));
 sky130_fd_sc_hd__a22o_1 _18890_ (.A1(_08289_),
    .A2(_08292_),
    .B1(_08589_),
    .B2(_08592_),
    .X(_08598_));
 sky130_fd_sc_hd__nand4_4 _18891_ (.A(_08289_),
    .B(_08292_),
    .C(_08589_),
    .D(_08592_),
    .Y(_08599_));
 sky130_fd_sc_hd__o21ai_1 _18892_ (.A1(_08591_),
    .A2(_08595_),
    .B1(_08597_),
    .Y(_08600_));
 sky130_fd_sc_hd__a22oi_4 _18893_ (.A1(_08230_),
    .A2(_08234_),
    .B1(_08172_),
    .B2(_08237_),
    .Y(_08602_));
 sky130_fd_sc_hd__a31o_1 _18894_ (.A1(_08169_),
    .A2(_08171_),
    .A3(_08237_),
    .B1(_08235_),
    .X(_08603_));
 sky130_fd_sc_hd__o21a_2 _18895_ (.A1(_08145_),
    .A2(_08156_),
    .B1(_08155_),
    .X(_08604_));
 sky130_fd_sc_hd__a21o_2 _18896_ (.A1(_08179_),
    .A2(_08190_),
    .B1(_08187_),
    .X(_08605_));
 sky130_fd_sc_hd__or3b_2 _18897_ (.A(net60),
    .B(_04201_),
    .C_N(net59),
    .X(_08606_));
 sky130_fd_sc_hd__o211ai_4 _18898_ (.A1(net175),
    .A2(_06759_),
    .B1(_05227_),
    .C1(net196),
    .Y(_08607_));
 sky130_fd_sc_hd__o211ai_4 _18899_ (.A1(net175),
    .A2(_06451_),
    .B1(_05688_),
    .C1(net199),
    .Y(_08608_));
 sky130_fd_sc_hd__or3b_4 _18900_ (.A(net61),
    .B(_04179_),
    .C_N(net60),
    .X(_08609_));
 sky130_fd_sc_hd__o2111a_1 _18901_ (.A1(_04201_),
    .A2(_05260_),
    .B1(_08607_),
    .C1(_08608_),
    .D1(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__o2111ai_4 _18902_ (.A1(_04201_),
    .A2(_05260_),
    .B1(_08607_),
    .C1(_08608_),
    .D1(_08609_),
    .Y(_08611_));
 sky130_fd_sc_hd__a22oi_4 _18903_ (.A1(_08606_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_08609_),
    .Y(_08613_));
 sky130_fd_sc_hd__a22o_1 _18904_ (.A1(_08606_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_08609_),
    .X(_08614_));
 sky130_fd_sc_hd__a32o_1 _18905_ (.A1(net201),
    .A2(_06221_),
    .A3(net292),
    .B1(_06848_),
    .B2(net17),
    .X(_08615_));
 sky130_fd_sc_hd__o21bai_4 _18906_ (.A1(_08610_),
    .A2(_08613_),
    .B1_N(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__nand2_1 _18907_ (.A(_08611_),
    .B(_08615_),
    .Y(_08617_));
 sky130_fd_sc_hd__nand3_2 _18908_ (.A(_08611_),
    .B(_08614_),
    .C(_08615_),
    .Y(_08618_));
 sky130_fd_sc_hd__a21oi_4 _18909_ (.A1(_08616_),
    .A2(_08618_),
    .B1(_08605_),
    .Y(_08619_));
 sky130_fd_sc_hd__a21o_1 _18910_ (.A1(_08616_),
    .A2(_08618_),
    .B1(_08605_),
    .X(_08620_));
 sky130_fd_sc_hd__o211a_1 _18911_ (.A1(_08613_),
    .A2(_08617_),
    .B1(_08616_),
    .C1(_08605_),
    .X(_08621_));
 sky130_fd_sc_hd__o211ai_4 _18912_ (.A1(_08613_),
    .A2(_08617_),
    .B1(_08616_),
    .C1(_08605_),
    .Y(_08622_));
 sky130_fd_sc_hd__o21a_1 _18913_ (.A1(_08619_),
    .A2(_08621_),
    .B1(_08604_),
    .X(_08624_));
 sky130_fd_sc_hd__o211a_1 _18914_ (.A1(_08154_),
    .A2(_08161_),
    .B1(_08620_),
    .C1(_08622_),
    .X(_08625_));
 sky130_fd_sc_hd__and3_2 _18915_ (.A(_08620_),
    .B(_08622_),
    .C(_08604_),
    .X(_08626_));
 sky130_fd_sc_hd__o2111ai_4 _18916_ (.A1(_08160_),
    .A2(_08156_),
    .B1(_08155_),
    .C1(_08622_),
    .D1(_08620_),
    .Y(_08627_));
 sky130_fd_sc_hd__o22a_2 _18917_ (.A1(_08154_),
    .A2(_08161_),
    .B1(_08619_),
    .B2(_08621_),
    .X(_08628_));
 sky130_fd_sc_hd__o22ai_2 _18918_ (.A1(_08154_),
    .A2(_08161_),
    .B1(_08619_),
    .B2(_08621_),
    .Y(_08629_));
 sky130_fd_sc_hd__nand2_1 _18919_ (.A(_08627_),
    .B(_08629_),
    .Y(_08630_));
 sky130_fd_sc_hd__o21ai_2 _18920_ (.A1(_08218_),
    .A2(_08222_),
    .B1(_08199_),
    .Y(_08631_));
 sky130_fd_sc_hd__a21oi_4 _18921_ (.A1(_08226_),
    .A2(_08198_),
    .B1(_08223_),
    .Y(_08632_));
 sky130_fd_sc_hd__and3b_1 _18922_ (.A_N(net59),
    .B(net20),
    .C(net58),
    .X(_08633_));
 sky130_fd_sc_hd__o311a_1 _18923_ (.A1(net245),
    .A2(net241),
    .A3(_07074_),
    .B1(_04889_),
    .C1(_07072_),
    .X(_08635_));
 sky130_fd_sc_hd__a31o_1 _18924_ (.A1(_07072_),
    .A2(net168),
    .A3(_04889_),
    .B1(_08633_),
    .X(_08636_));
 sky130_fd_sc_hd__nor2_1 _18925_ (.A(_04223_),
    .B(net316),
    .Y(_08637_));
 sky130_fd_sc_hd__a31oi_4 _18926_ (.A1(_07499_),
    .A2(net167),
    .A3(_04627_),
    .B1(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__a31o_1 _18927_ (.A1(_07499_),
    .A2(net167),
    .A3(_04627_),
    .B1(_08637_),
    .X(_08639_));
 sky130_fd_sc_hd__nor2_1 _18928_ (.A(_04245_),
    .B(_04375_),
    .Y(_08640_));
 sky130_fd_sc_hd__a31oi_4 _18929_ (.A1(_07771_),
    .A2(_04342_),
    .A3(_07769_),
    .B1(_08640_),
    .Y(_08641_));
 sky130_fd_sc_hd__a31o_1 _18930_ (.A1(_07771_),
    .A2(_04342_),
    .A3(_07769_),
    .B1(_08640_),
    .X(_08642_));
 sky130_fd_sc_hd__nor2_2 _18931_ (.A(_08638_),
    .B(_08641_),
    .Y(_08643_));
 sky130_fd_sc_hd__nand2_2 _18932_ (.A(_08639_),
    .B(_08642_),
    .Y(_08644_));
 sky130_fd_sc_hd__nand2_2 _18933_ (.A(_08638_),
    .B(_08641_),
    .Y(_08646_));
 sky130_fd_sc_hd__a211o_1 _18934_ (.A1(_08644_),
    .A2(_08646_),
    .B1(_08633_),
    .C1(_08635_),
    .X(_08647_));
 sky130_fd_sc_hd__o211ai_2 _18935_ (.A1(_08633_),
    .A2(_08635_),
    .B1(_08644_),
    .C1(_08646_),
    .Y(_08648_));
 sky130_fd_sc_hd__nand3b_4 _18936_ (.A_N(_08636_),
    .B(_08644_),
    .C(_08646_),
    .Y(_08649_));
 sky130_fd_sc_hd__a21bo_2 _18937_ (.A1(_08644_),
    .A2(_08646_),
    .B1_N(_08636_),
    .X(_08650_));
 sky130_fd_sc_hd__a21o_1 _18938_ (.A1(_08202_),
    .A2(_08213_),
    .B1(_08214_),
    .X(_08651_));
 sky130_fd_sc_hd__a21oi_4 _18939_ (.A1(_08202_),
    .A2(_08213_),
    .B1(_08214_),
    .Y(_08652_));
 sky130_fd_sc_hd__o311a_1 _18940_ (.A1(net175),
    .A2(_07074_),
    .A3(_08206_),
    .B1(_04484_),
    .C1(_08204_),
    .X(_08653_));
 sky130_fd_sc_hd__nor2_1 _18941_ (.A(_04256_),
    .B(_04331_),
    .Y(_08654_));
 sky130_fd_sc_hd__o32a_2 _18942_ (.A1(_04495_),
    .A2(_08203_),
    .A3(_08207_),
    .B1(_04331_),
    .B2(_04256_),
    .X(_08655_));
 sky130_fd_sc_hd__and2_4 _18943_ (.A(_04266_),
    .B(net57),
    .X(_08657_));
 sky130_fd_sc_hd__nand2_8 _18944_ (.A(_04266_),
    .B(net57),
    .Y(_08658_));
 sky130_fd_sc_hd__nor2_2 _18945_ (.A(net57),
    .B(_04266_),
    .Y(_08659_));
 sky130_fd_sc_hd__nand2b_4 _18946_ (.A_N(net57),
    .B(net56),
    .Y(_08660_));
 sky130_fd_sc_hd__nor2_1 _18947_ (.A(_08657_),
    .B(_08659_),
    .Y(_08661_));
 sky130_fd_sc_hd__nand2_1 _18948_ (.A(_08658_),
    .B(_08660_),
    .Y(_08662_));
 sky130_fd_sc_hd__a21o_1 _18949_ (.A1(_08658_),
    .A2(_08660_),
    .B1(_03176_),
    .X(_08663_));
 sky130_fd_sc_hd__a31oi_4 _18950_ (.A1(_05930_),
    .A2(_07766_),
    .A3(_04256_),
    .B1(net25),
    .Y(_08664_));
 sky130_fd_sc_hd__o21bai_4 _18951_ (.A1(_07076_),
    .A2(net268),
    .B1_N(net25),
    .Y(_08665_));
 sky130_fd_sc_hd__and4_4 _18952_ (.A(net204),
    .B(_04256_),
    .C(net25),
    .D(_07766_),
    .X(_08666_));
 sky130_fd_sc_hd__nand4_4 _18953_ (.A(_05930_),
    .B(_04256_),
    .C(net25),
    .D(_07766_),
    .Y(_08668_));
 sky130_fd_sc_hd__nor2_8 _18954_ (.A(net160),
    .B(_08666_),
    .Y(_08669_));
 sky130_fd_sc_hd__nand2_8 _18955_ (.A(_08665_),
    .B(net158),
    .Y(_08670_));
 sky130_fd_sc_hd__o21ai_2 _18956_ (.A1(net160),
    .A2(_08666_),
    .B1(net33),
    .Y(_08671_));
 sky130_fd_sc_hd__a211oi_2 _18957_ (.A1(net151),
    .A2(net158),
    .B1(_03286_),
    .C1(_08663_),
    .Y(_08672_));
 sky130_fd_sc_hd__a211o_1 _18958_ (.A1(net151),
    .A2(net158),
    .B1(_03286_),
    .C1(_08663_),
    .X(_08673_));
 sky130_fd_sc_hd__a22oi_4 _18959_ (.A1(net1),
    .A2(_08662_),
    .B1(_08670_),
    .B2(net33),
    .Y(_08674_));
 sky130_fd_sc_hd__o21ai_4 _18960_ (.A1(_03176_),
    .A2(_08661_),
    .B1(_08671_),
    .Y(_08675_));
 sky130_fd_sc_hd__o211ai_2 _18961_ (.A1(_08653_),
    .A2(_08654_),
    .B1(_08673_),
    .C1(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__o21ai_1 _18962_ (.A1(_08672_),
    .A2(_08674_),
    .B1(_08655_),
    .Y(_08677_));
 sky130_fd_sc_hd__o22ai_4 _18963_ (.A1(_08653_),
    .A2(_08654_),
    .B1(_08672_),
    .B2(_08674_),
    .Y(_08679_));
 sky130_fd_sc_hd__nand3_4 _18964_ (.A(_08675_),
    .B(_08655_),
    .C(_08673_),
    .Y(_08680_));
 sky130_fd_sc_hd__a21oi_4 _18965_ (.A1(_08679_),
    .A2(_08680_),
    .B1(_08652_),
    .Y(_08681_));
 sky130_fd_sc_hd__nand3_4 _18966_ (.A(_08677_),
    .B(_08651_),
    .C(_08676_),
    .Y(_08682_));
 sky130_fd_sc_hd__nand3_4 _18967_ (.A(_08652_),
    .B(_08679_),
    .C(_08680_),
    .Y(_08683_));
 sky130_fd_sc_hd__a32oi_4 _18968_ (.A1(_08652_),
    .A2(_08679_),
    .A3(_08680_),
    .B1(_08650_),
    .B2(_08649_),
    .Y(_08684_));
 sky130_fd_sc_hd__nand2_2 _18969_ (.A(_08684_),
    .B(_08682_),
    .Y(_08685_));
 sky130_fd_sc_hd__a22o_2 _18970_ (.A1(_08647_),
    .A2(_08648_),
    .B1(_08682_),
    .B2(_08683_),
    .X(_08686_));
 sky130_fd_sc_hd__a22o_2 _18971_ (.A1(_08649_),
    .A2(_08650_),
    .B1(_08682_),
    .B2(_08683_),
    .X(_08687_));
 sky130_fd_sc_hd__nand4_4 _18972_ (.A(_08649_),
    .B(_08650_),
    .C(_08682_),
    .D(_08683_),
    .Y(_08688_));
 sky130_fd_sc_hd__a22oi_4 _18973_ (.A1(_08224_),
    .A2(_08229_),
    .B1(_08687_),
    .B2(_08688_),
    .Y(_08690_));
 sky130_fd_sc_hd__nand4_4 _18974_ (.A(_08226_),
    .B(_08631_),
    .C(_08685_),
    .D(_08686_),
    .Y(_08691_));
 sky130_fd_sc_hd__a22oi_4 _18975_ (.A1(_08226_),
    .A2(_08631_),
    .B1(_08685_),
    .B2(_08686_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand3_4 _18976_ (.A(_08632_),
    .B(_08687_),
    .C(_08688_),
    .Y(_08693_));
 sky130_fd_sc_hd__o211ai_4 _18977_ (.A1(_08624_),
    .A2(_08625_),
    .B1(_08691_),
    .C1(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__o22ai_4 _18978_ (.A1(_08626_),
    .A2(_08628_),
    .B1(_08690_),
    .B2(_08692_),
    .Y(_08695_));
 sky130_fd_sc_hd__a32oi_4 _18979_ (.A1(_08632_),
    .A2(_08687_),
    .A3(_08688_),
    .B1(_08629_),
    .B2(_08627_),
    .Y(_08696_));
 sky130_fd_sc_hd__o211ai_4 _18980_ (.A1(_08626_),
    .A2(_08628_),
    .B1(_08691_),
    .C1(_08693_),
    .Y(_08697_));
 sky130_fd_sc_hd__o22ai_4 _18981_ (.A1(_08624_),
    .A2(_08625_),
    .B1(_08690_),
    .B2(_08692_),
    .Y(_08698_));
 sky130_fd_sc_hd__o211a_1 _18982_ (.A1(_08235_),
    .A2(_08241_),
    .B1(_08697_),
    .C1(_08698_),
    .X(_08699_));
 sky130_fd_sc_hd__o211ai_4 _18983_ (.A1(_08235_),
    .A2(_08241_),
    .B1(_08697_),
    .C1(_08698_),
    .Y(_08701_));
 sky130_fd_sc_hd__a21boi_2 _18984_ (.A1(_08697_),
    .A2(_08698_),
    .B1_N(_08602_),
    .Y(_08702_));
 sky130_fd_sc_hd__nand3_4 _18985_ (.A(_08695_),
    .B(_08602_),
    .C(_08694_),
    .Y(_08703_));
 sky130_fd_sc_hd__nand4_2 _18986_ (.A(_08598_),
    .B(_08599_),
    .C(_08701_),
    .D(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__a22o_1 _18987_ (.A1(_08598_),
    .A2(_08599_),
    .B1(_08701_),
    .B2(_08703_),
    .X(_08705_));
 sky130_fd_sc_hd__a32oi_4 _18988_ (.A1(_08695_),
    .A2(_08602_),
    .A3(_08694_),
    .B1(_08599_),
    .B2(_08598_),
    .Y(_08706_));
 sky130_fd_sc_hd__and4_1 _18989_ (.A(_08596_),
    .B(_08597_),
    .C(_08701_),
    .D(_08703_),
    .X(_08707_));
 sky130_fd_sc_hd__o2111ai_4 _18990_ (.A1(_08591_),
    .A2(_08595_),
    .B1(_08597_),
    .C1(_08701_),
    .D1(_08703_),
    .Y(_08708_));
 sky130_fd_sc_hd__a22oi_2 _18991_ (.A1(_08596_),
    .A2(_08597_),
    .B1(_08701_),
    .B2(_08703_),
    .Y(_08709_));
 sky130_fd_sc_hd__a22o_1 _18992_ (.A1(_08596_),
    .A2(_08597_),
    .B1(_08701_),
    .B2(_08703_),
    .X(_08710_));
 sky130_fd_sc_hd__nand2_1 _18993_ (.A(_08710_),
    .B(_08539_),
    .Y(_08712_));
 sky130_fd_sc_hd__a221oi_4 _18994_ (.A1(_08706_),
    .A2(_08701_),
    .B1(_08311_),
    .B2(_08245_),
    .C1(_08709_),
    .Y(_08713_));
 sky130_fd_sc_hd__nand3_2 _18995_ (.A(_08710_),
    .B(_08539_),
    .C(_08708_),
    .Y(_08714_));
 sky130_fd_sc_hd__o211a_2 _18996_ (.A1(_08246_),
    .A2(_08538_),
    .B1(_08704_),
    .C1(_08705_),
    .X(_08715_));
 sky130_fd_sc_hd__o211ai_4 _18997_ (.A1(_08246_),
    .A2(_08538_),
    .B1(_08704_),
    .C1(_08705_),
    .Y(_08716_));
 sky130_fd_sc_hd__nand3_4 _18998_ (.A(_08537_),
    .B(_08714_),
    .C(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__o22ai_4 _18999_ (.A1(_08531_),
    .A2(_08534_),
    .B1(_08713_),
    .B2(_08715_),
    .Y(_08718_));
 sky130_fd_sc_hd__nand4_2 _19000_ (.A(_08528_),
    .B(_08530_),
    .C(_08714_),
    .D(_08716_),
    .Y(_08719_));
 sky130_fd_sc_hd__a22o_1 _19001_ (.A1(_08528_),
    .A2(_08530_),
    .B1(_08714_),
    .B2(_08716_),
    .X(_08720_));
 sky130_fd_sc_hd__a2bb2oi_4 _19002_ (.A1_N(_08313_),
    .A2_N(_08318_),
    .B1(_08717_),
    .B2(_08718_),
    .Y(_08721_));
 sky130_fd_sc_hd__o211ai_4 _19003_ (.A1(_08313_),
    .A2(_08318_),
    .B1(_08719_),
    .C1(_08720_),
    .Y(_08723_));
 sky130_fd_sc_hd__a2bb2oi_2 _19004_ (.A1_N(_08315_),
    .A2_N(_08450_),
    .B1(_08719_),
    .B2(_08720_),
    .Y(_08724_));
 sky130_fd_sc_hd__o2111ai_4 _19005_ (.A1(_08134_),
    .A2(_08315_),
    .B1(_08717_),
    .C1(_08718_),
    .D1(_08314_),
    .Y(_08725_));
 sky130_fd_sc_hd__o211ai_2 _19006_ (.A1(_08439_),
    .A2(_08443_),
    .B1(_08723_),
    .C1(_08725_),
    .Y(_08726_));
 sky130_fd_sc_hd__o22ai_2 _19007_ (.A1(_08444_),
    .A2(_08446_),
    .B1(_08721_),
    .B2(_08724_),
    .Y(_08727_));
 sky130_fd_sc_hd__a32oi_4 _19008_ (.A1(_08451_),
    .A2(_08717_),
    .A3(_08718_),
    .B1(_08448_),
    .B2(_08445_),
    .Y(_08728_));
 sky130_fd_sc_hd__o21ai_1 _19009_ (.A1(_08444_),
    .A2(_08446_),
    .B1(_08725_),
    .Y(_08729_));
 sky130_fd_sc_hd__o211a_1 _19010_ (.A1(_08444_),
    .A2(_08446_),
    .B1(_08723_),
    .C1(_08725_),
    .X(_08730_));
 sky130_fd_sc_hd__o22ai_2 _19011_ (.A1(_08439_),
    .A2(_08443_),
    .B1(_08721_),
    .B2(_08724_),
    .Y(_08731_));
 sky130_fd_sc_hd__nand2_1 _19012_ (.A(_08363_),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__o211ai_2 _19013_ (.A1(_08721_),
    .A2(_08729_),
    .B1(_08731_),
    .C1(_08363_),
    .Y(_08734_));
 sky130_fd_sc_hd__o211ai_4 _19014_ (.A1(_08325_),
    .A2(_08362_),
    .B1(_08726_),
    .C1(_08727_),
    .Y(_08735_));
 sky130_fd_sc_hd__o211ai_2 _19015_ (.A1(_08730_),
    .A2(_08732_),
    .B1(_08735_),
    .C1(_08361_),
    .Y(_08736_));
 sky130_fd_sc_hd__a21o_1 _19016_ (.A1(_08734_),
    .A2(_08735_),
    .B1(_08361_),
    .X(_08737_));
 sky130_fd_sc_hd__a21o_1 _19017_ (.A1(_08734_),
    .A2(_08735_),
    .B1(_08360_),
    .X(_08738_));
 sky130_fd_sc_hd__o211ai_2 _19018_ (.A1(_08730_),
    .A2(_08732_),
    .B1(_08735_),
    .C1(_08360_),
    .Y(_08739_));
 sky130_fd_sc_hd__a21oi_1 _19019_ (.A1(_08738_),
    .A2(_08739_),
    .B1(_08358_),
    .Y(_08740_));
 sky130_fd_sc_hd__nand3_4 _19020_ (.A(_08737_),
    .B(_08357_),
    .C(_08736_),
    .Y(_08741_));
 sky130_fd_sc_hd__and3_1 _19021_ (.A(_08358_),
    .B(_08738_),
    .C(_08739_),
    .X(_08742_));
 sky130_fd_sc_hd__nand3_2 _19022_ (.A(_08358_),
    .B(_08738_),
    .C(_08739_),
    .Y(_08743_));
 sky130_fd_sc_hd__a31oi_1 _19023_ (.A1(_08358_),
    .A2(_08738_),
    .A3(_08739_),
    .B1(_08029_),
    .Y(_08745_));
 sky130_fd_sc_hd__and4bb_2 _19024_ (.A_N(_07654_),
    .B_N(_08028_),
    .C(_08741_),
    .D(_08743_),
    .X(_08746_));
 sky130_fd_sc_hd__nand3b_4 _19025_ (.A_N(_08029_),
    .B(_08741_),
    .C(_08743_),
    .Y(_08747_));
 sky130_fd_sc_hd__o2bb2ai_4 _19026_ (.A1_N(_08741_),
    .A2_N(_08743_),
    .B1(_07654_),
    .B2(_08028_),
    .Y(_08748_));
 sky130_fd_sc_hd__o2bb2ai_2 _19027_ (.A1_N(_08747_),
    .A2_N(_08748_),
    .B1(_07961_),
    .B2(_08344_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand2_1 _19028_ (.A(_08748_),
    .B(_08346_),
    .Y(_08750_));
 sky130_fd_sc_hd__nand3_1 _19029_ (.A(_08748_),
    .B(_08346_),
    .C(_08747_),
    .Y(_08751_));
 sky130_fd_sc_hd__a22o_1 _19030_ (.A1(_08352_),
    .A2(_08356_),
    .B1(_08749_),
    .B2(_08751_),
    .X(_08752_));
 sky130_fd_sc_hd__o2111ai_1 _19031_ (.A1(_08746_),
    .A2(_08750_),
    .B1(_08749_),
    .C1(_08352_),
    .D1(_08356_),
    .Y(_08753_));
 sky130_fd_sc_hd__nand2_1 _19032_ (.A(_08752_),
    .B(_08753_),
    .Y(net89));
 sky130_fd_sc_hd__o2bb2ai_1 _19033_ (.A1_N(_08361_),
    .A2_N(_08735_),
    .B1(_08730_),
    .B2(_08732_),
    .Y(_08755_));
 sky130_fd_sc_hd__a21boi_1 _19034_ (.A1(_08361_),
    .A2(_08735_),
    .B1_N(_08734_),
    .Y(_08756_));
 sky130_fd_sc_hd__o22a_1 _19035_ (.A1(_08002_),
    .A2(_08437_),
    .B1(_08364_),
    .B2(_08431_),
    .X(_08757_));
 sky130_fd_sc_hd__a31o_1 _19036_ (.A1(_08365_),
    .A2(_08429_),
    .A3(_08430_),
    .B1(_08441_),
    .X(_08758_));
 sky130_fd_sc_hd__a21o_1 _19037_ (.A1(_08449_),
    .A2(_08723_),
    .B1(_08724_),
    .X(_08759_));
 sky130_fd_sc_hd__a21oi_1 _19038_ (.A1(_08449_),
    .A2(_08723_),
    .B1(_08724_),
    .Y(_08760_));
 sky130_fd_sc_hd__a21boi_4 _19039_ (.A1(_08387_),
    .A2(_08389_),
    .B1_N(_08388_),
    .Y(_08761_));
 sky130_fd_sc_hd__a22oi_4 _19040_ (.A1(_06541_),
    .A2(net273),
    .B1(_06326_),
    .B2(net30),
    .Y(_08762_));
 sky130_fd_sc_hd__a32o_1 _19041_ (.A1(_06486_),
    .A2(net260),
    .A3(net273),
    .B1(_06326_),
    .B2(net30),
    .X(_08763_));
 sky130_fd_sc_hd__a32oi_4 _19042_ (.A1(_07242_),
    .A2(net257),
    .A3(net274),
    .B1(_06029_),
    .B2(net31),
    .Y(_08764_));
 sky130_fd_sc_hd__or3b_1 _19043_ (.A(_03949_),
    .B(net48),
    .C_N(net47),
    .X(_08766_));
 sky130_fd_sc_hd__o211ai_2 _19044_ (.A1(net260),
    .A2(_08656_),
    .B1(net275),
    .C1(_08700_),
    .Y(_08767_));
 sky130_fd_sc_hd__a21oi_2 _19045_ (.A1(_08766_),
    .A2(_08767_),
    .B1(_08764_),
    .Y(_08768_));
 sky130_fd_sc_hd__a21o_2 _19046_ (.A1(_08766_),
    .A2(_08767_),
    .B1(_08764_),
    .X(_08769_));
 sky130_fd_sc_hd__o211a_1 _19047_ (.A1(_03949_),
    .A2(_05766_),
    .B1(_08767_),
    .C1(_08764_),
    .X(_08770_));
 sky130_fd_sc_hd__o221ai_2 _19048_ (.A1(_08711_),
    .A2(_05763_),
    .B1(_05766_),
    .B2(_03949_),
    .C1(_08764_),
    .Y(_08771_));
 sky130_fd_sc_hd__and3_1 _19049_ (.A(_08763_),
    .B(_08769_),
    .C(_08771_),
    .X(_08772_));
 sky130_fd_sc_hd__nand3_2 _19050_ (.A(_08763_),
    .B(_08769_),
    .C(_08771_),
    .Y(_08773_));
 sky130_fd_sc_hd__o21ai_2 _19051_ (.A1(_08768_),
    .A2(_08770_),
    .B1(_08762_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand2_1 _19052_ (.A(_08773_),
    .B(_08774_),
    .Y(_08775_));
 sky130_fd_sc_hd__nor2_1 _19053_ (.A(_08504_),
    .B(_08509_),
    .Y(_08777_));
 sky130_fd_sc_hd__a21o_1 _19054_ (.A1(_08504_),
    .A2(_08512_),
    .B1(_08509_),
    .X(_08778_));
 sky130_fd_sc_hd__a31o_1 _19055_ (.A1(_08506_),
    .A2(_08507_),
    .A3(_08508_),
    .B1(_08777_),
    .X(_08779_));
 sky130_fd_sc_hd__o2bb2ai_2 _19056_ (.A1_N(_08773_),
    .A2_N(_08774_),
    .B1(_08777_),
    .B2(_08511_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand3_2 _19057_ (.A(_08778_),
    .B(_08774_),
    .C(_08773_),
    .Y(_08781_));
 sky130_fd_sc_hd__a21o_1 _19058_ (.A1(_08372_),
    .A2(_08375_),
    .B1(_08373_),
    .X(_08782_));
 sky130_fd_sc_hd__a21oi_1 _19059_ (.A1(_08780_),
    .A2(_08781_),
    .B1(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__a21o_1 _19060_ (.A1(_08780_),
    .A2(_08781_),
    .B1(_08782_),
    .X(_08784_));
 sky130_fd_sc_hd__and3_1 _19061_ (.A(_08780_),
    .B(_08781_),
    .C(_08782_),
    .X(_08785_));
 sky130_fd_sc_hd__nand3_4 _19062_ (.A(_08780_),
    .B(_08781_),
    .C(_08782_),
    .Y(_08786_));
 sky130_fd_sc_hd__nand2_1 _19063_ (.A(_08784_),
    .B(_08786_),
    .Y(_08788_));
 sky130_fd_sc_hd__o2bb2ai_2 _19064_ (.A1_N(_08516_),
    .A2_N(_08500_),
    .B1(_08497_),
    .B2(_08501_),
    .Y(_08789_));
 sky130_fd_sc_hd__o2bb2a_2 _19065_ (.A1_N(_08516_),
    .A2_N(_08500_),
    .B1(_08497_),
    .B2(_08501_),
    .X(_08790_));
 sky130_fd_sc_hd__o21ai_2 _19066_ (.A1(_08783_),
    .A2(_08785_),
    .B1(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__and3_1 _19067_ (.A(_08784_),
    .B(_08789_),
    .C(_08786_),
    .X(_08792_));
 sky130_fd_sc_hd__nand3_2 _19068_ (.A(_08789_),
    .B(_08786_),
    .C(_08784_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand2_1 _19069_ (.A(_08380_),
    .B(_08385_),
    .Y(_08794_));
 sky130_fd_sc_hd__a21oi_1 _19070_ (.A1(_08791_),
    .A2(_08793_),
    .B1(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__a21o_1 _19071_ (.A1(_08791_),
    .A2(_08793_),
    .B1(_08794_),
    .X(_08796_));
 sky130_fd_sc_hd__a22oi_4 _19072_ (.A1(_08380_),
    .A2(_08385_),
    .B1(_08788_),
    .B2(_08790_),
    .Y(_08797_));
 sky130_fd_sc_hd__and3_1 _19073_ (.A(_08791_),
    .B(_08793_),
    .C(_08794_),
    .X(_08799_));
 sky130_fd_sc_hd__o21ai_1 _19074_ (.A1(_08788_),
    .A2(_08790_),
    .B1(_08797_),
    .Y(_08800_));
 sky130_fd_sc_hd__nand4_2 _19075_ (.A(_08380_),
    .B(_08385_),
    .C(_08791_),
    .D(_08793_),
    .Y(_08801_));
 sky130_fd_sc_hd__a22o_1 _19076_ (.A1(_08380_),
    .A2(_08385_),
    .B1(_08791_),
    .B2(_08793_),
    .X(_08802_));
 sky130_fd_sc_hd__o21ai_1 _19077_ (.A1(_08795_),
    .A2(_08799_),
    .B1(_08761_),
    .Y(_08803_));
 sky130_fd_sc_hd__a21oi_2 _19078_ (.A1(_08801_),
    .A2(_08802_),
    .B1(_08761_),
    .Y(_08804_));
 sky130_fd_sc_hd__nand3b_4 _19079_ (.A_N(_08761_),
    .B(_08796_),
    .C(_08800_),
    .Y(_08805_));
 sky130_fd_sc_hd__o2bb2a_1 _19080_ (.A1_N(_04463_),
    .A2_N(_08005_),
    .B1(_08007_),
    .B2(_03396_),
    .X(_08806_));
 sky130_fd_sc_hd__nand2_1 _19081_ (.A(_08418_),
    .B(_08401_),
    .Y(_08807_));
 sky130_fd_sc_hd__a21o_1 _19082_ (.A1(_08404_),
    .A2(_08411_),
    .B1(_08409_),
    .X(_08808_));
 sky130_fd_sc_hd__a32oi_2 _19083_ (.A1(net266),
    .A2(net301),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net27),
    .Y(_08810_));
 sky130_fd_sc_hd__a32o_1 _19084_ (.A1(net266),
    .A2(net301),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net27),
    .X(_08811_));
 sky130_fd_sc_hd__or3b_1 _19085_ (.A(_03725_),
    .B(net52),
    .C_N(net51),
    .X(_08812_));
 sky130_fd_sc_hd__o211ai_2 _19086_ (.A1(_04747_),
    .A2(_05436_),
    .B1(_07223_),
    .C1(_05414_),
    .Y(_08813_));
 sky130_fd_sc_hd__or3_1 _19087_ (.A(net51),
    .B(_04190_),
    .C(_03835_),
    .X(_08814_));
 sky130_fd_sc_hd__nand4_2 _19088_ (.A(_04190_),
    .B(_05841_),
    .C(net265),
    .D(net51),
    .Y(_08815_));
 sky130_fd_sc_hd__a22oi_1 _19089_ (.A1(_08812_),
    .A2(_08813_),
    .B1(_08814_),
    .B2(_08815_),
    .Y(_08816_));
 sky130_fd_sc_hd__a22o_1 _19090_ (.A1(_08812_),
    .A2(_08813_),
    .B1(_08814_),
    .B2(_08815_),
    .X(_08817_));
 sky130_fd_sc_hd__o2111a_1 _19091_ (.A1(_03725_),
    .A2(_07226_),
    .B1(_08813_),
    .C1(_08814_),
    .D1(_08815_),
    .X(_08818_));
 sky130_fd_sc_hd__o2111ai_1 _19092_ (.A1(_03725_),
    .A2(_07226_),
    .B1(_08813_),
    .C1(_08814_),
    .D1(_08815_),
    .Y(_08819_));
 sky130_fd_sc_hd__o21ai_1 _19093_ (.A1(_08816_),
    .A2(_08818_),
    .B1(_08810_),
    .Y(_08821_));
 sky130_fd_sc_hd__nand3_1 _19094_ (.A(_08811_),
    .B(_08817_),
    .C(_08819_),
    .Y(_08822_));
 sky130_fd_sc_hd__nand3_1 _19095_ (.A(_08808_),
    .B(_08821_),
    .C(_08822_),
    .Y(_08823_));
 sky130_fd_sc_hd__a21o_1 _19096_ (.A1(_08821_),
    .A2(_08822_),
    .B1(_08808_),
    .X(_08824_));
 sky130_fd_sc_hd__a32o_1 _19097_ (.A1(_07642_),
    .A2(_04747_),
    .A3(net313),
    .B1(net26),
    .B2(_07643_),
    .X(_08825_));
 sky130_fd_sc_hd__a21o_1 _19098_ (.A1(_08823_),
    .A2(_08824_),
    .B1(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__nand3_2 _19099_ (.A(_08823_),
    .B(_08824_),
    .C(_08825_),
    .Y(_08827_));
 sky130_fd_sc_hd__a22oi_4 _19100_ (.A1(_08417_),
    .A2(_08807_),
    .B1(_08826_),
    .B2(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__and4_2 _19101_ (.A(_08417_),
    .B(_08807_),
    .C(_08826_),
    .D(_08827_),
    .X(_08829_));
 sky130_fd_sc_hd__nor3_2 _19102_ (.A(_08806_),
    .B(_08828_),
    .C(_08829_),
    .Y(_08830_));
 sky130_fd_sc_hd__o21a_1 _19103_ (.A1(_08828_),
    .A2(_08829_),
    .B1(_08806_),
    .X(_08832_));
 sky130_fd_sc_hd__nor2_1 _19104_ (.A(_08830_),
    .B(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__o2bb2ai_2 _19105_ (.A1_N(_08803_),
    .A2_N(_08805_),
    .B1(_08830_),
    .B2(_08832_),
    .Y(_08834_));
 sky130_fd_sc_hd__a311o_4 _19106_ (.A1(_08802_),
    .A2(_08761_),
    .A3(_08801_),
    .B1(_08830_),
    .C1(_08832_),
    .X(_08835_));
 sky130_fd_sc_hd__nand3_1 _19107_ (.A(_08833_),
    .B(_08805_),
    .C(_08803_),
    .Y(_08836_));
 sky130_fd_sc_hd__a22oi_1 _19108_ (.A1(_08526_),
    .A2(_08533_),
    .B1(_08834_),
    .B2(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__a22o_1 _19109_ (.A1(_08526_),
    .A2(_08533_),
    .B1(_08834_),
    .B2(_08836_),
    .X(_08838_));
 sky130_fd_sc_hd__o2111a_1 _19110_ (.A1(_08804_),
    .A2(_08835_),
    .B1(_08834_),
    .C1(_08526_),
    .D1(_08533_),
    .X(_08839_));
 sky130_fd_sc_hd__o2111ai_4 _19111_ (.A1(_08804_),
    .A2(_08835_),
    .B1(_08834_),
    .C1(_08526_),
    .D1(_08533_),
    .Y(_08840_));
 sky130_fd_sc_hd__a21o_1 _19112_ (.A1(_08395_),
    .A2(_08427_),
    .B1(_08396_),
    .X(_08841_));
 sky130_fd_sc_hd__a21oi_2 _19113_ (.A1(_08838_),
    .A2(_08840_),
    .B1(_08841_),
    .Y(_08843_));
 sky130_fd_sc_hd__o21bai_1 _19114_ (.A1(_08837_),
    .A2(_08839_),
    .B1_N(_08841_),
    .Y(_08844_));
 sky130_fd_sc_hd__and3_2 _19115_ (.A(_08838_),
    .B(_08840_),
    .C(_08841_),
    .X(_08845_));
 sky130_fd_sc_hd__nand3_1 _19116_ (.A(_08838_),
    .B(_08840_),
    .C(_08841_),
    .Y(_08846_));
 sky130_fd_sc_hd__nand2_1 _19117_ (.A(_08844_),
    .B(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__a31oi_2 _19118_ (.A1(_08539_),
    .A2(_08708_),
    .A3(_08710_),
    .B1(_08536_),
    .Y(_08848_));
 sky130_fd_sc_hd__nand2_1 _19119_ (.A(_08537_),
    .B(_08714_),
    .Y(_08849_));
 sky130_fd_sc_hd__o2bb2ai_2 _19120_ (.A1_N(_08536_),
    .A2_N(_08716_),
    .B1(_08707_),
    .B2(_08712_),
    .Y(_08850_));
 sky130_fd_sc_hd__o22a_1 _19121_ (.A1(_08707_),
    .A2(_08712_),
    .B1(_08537_),
    .B2(_08715_),
    .X(_08851_));
 sky130_fd_sc_hd__a31oi_4 _19122_ (.A1(_08647_),
    .A2(_08648_),
    .A3(_08683_),
    .B1(_08681_),
    .Y(_08852_));
 sky130_fd_sc_hd__o211ai_1 _19123_ (.A1(net168),
    .A2(_07765_),
    .B1(_04627_),
    .C1(_07771_),
    .Y(_08854_));
 sky130_fd_sc_hd__or3b_1 _19124_ (.A(net58),
    .B(_04245_),
    .C_N(net55),
    .X(_08855_));
 sky130_fd_sc_hd__a32oi_4 _19125_ (.A1(_07771_),
    .A2(_04627_),
    .A3(_07769_),
    .B1(_04649_),
    .B2(net22),
    .Y(_08856_));
 sky130_fd_sc_hd__o211ai_4 _19126_ (.A1(net168),
    .A2(_08206_),
    .B1(_04342_),
    .C1(_08204_),
    .Y(_08857_));
 sky130_fd_sc_hd__or3b_1 _19127_ (.A(net55),
    .B(_04256_),
    .C_N(net44),
    .X(_08858_));
 sky130_fd_sc_hd__a21oi_2 _19128_ (.A1(_08857_),
    .A2(_08858_),
    .B1(_08856_),
    .Y(_08859_));
 sky130_fd_sc_hd__a22o_1 _19129_ (.A1(_08854_),
    .A2(_08855_),
    .B1(_08857_),
    .B2(_08858_),
    .X(_08860_));
 sky130_fd_sc_hd__o311a_2 _19130_ (.A1(_04353_),
    .A2(_08203_),
    .A3(net154),
    .B1(_08858_),
    .C1(_08856_),
    .X(_08861_));
 sky130_fd_sc_hd__o211ai_4 _19131_ (.A1(_04256_),
    .A2(_04375_),
    .B1(_08857_),
    .C1(_08856_),
    .Y(_08862_));
 sky130_fd_sc_hd__and3b_1 _19132_ (.A_N(net59),
    .B(net21),
    .C(net58),
    .X(_08863_));
 sky130_fd_sc_hd__o311a_1 _19133_ (.A1(net245),
    .A2(_05928_),
    .A3(_07501_),
    .B1(_04889_),
    .C1(_07499_),
    .X(_08865_));
 sky130_fd_sc_hd__a31o_1 _19134_ (.A1(_07499_),
    .A2(net167),
    .A3(_04889_),
    .B1(_08863_),
    .X(_08866_));
 sky130_fd_sc_hd__a21oi_2 _19135_ (.A1(_08860_),
    .A2(_08862_),
    .B1(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__o21bai_2 _19136_ (.A1(_08859_),
    .A2(_08861_),
    .B1_N(_08866_),
    .Y(_08868_));
 sky130_fd_sc_hd__o21ai_2 _19137_ (.A1(_08863_),
    .A2(_08865_),
    .B1(_08860_),
    .Y(_08869_));
 sky130_fd_sc_hd__o211a_1 _19138_ (.A1(_08863_),
    .A2(_08865_),
    .B1(_08860_),
    .C1(_08862_),
    .X(_08870_));
 sky130_fd_sc_hd__o21ai_1 _19139_ (.A1(_08861_),
    .A2(_08869_),
    .B1(_08868_),
    .Y(_08871_));
 sky130_fd_sc_hd__o21ai_4 _19140_ (.A1(_08663_),
    .A2(_08671_),
    .B1(_08655_),
    .Y(_08872_));
 sky130_fd_sc_hd__o2bb2a_2 _19141_ (.A1_N(net12),
    .A2_N(_08659_),
    .B1(_08658_),
    .B2(_04528_),
    .X(_08873_));
 sky130_fd_sc_hd__a22o_1 _19142_ (.A1(net12),
    .A2(_08659_),
    .B1(_04539_),
    .B2(_08657_),
    .X(_08874_));
 sky130_fd_sc_hd__a31oi_4 _19143_ (.A1(net204),
    .A2(_07766_),
    .A3(_04256_),
    .B1(_03286_),
    .Y(_08876_));
 sky130_fd_sc_hd__a311oi_4 _19144_ (.A1(_05930_),
    .A2(_07766_),
    .A3(_04256_),
    .B1(net25),
    .C1(_03286_),
    .Y(_08877_));
 sky130_fd_sc_hd__nand3_4 _19145_ (.A(net163),
    .B(net33),
    .C(net319),
    .Y(_08878_));
 sky130_fd_sc_hd__and3_2 _19146_ (.A(_08874_),
    .B(net33),
    .C(_04277_),
    .X(_08879_));
 sky130_fd_sc_hd__a31oi_2 _19147_ (.A1(net163),
    .A2(net33),
    .A3(_04277_),
    .B1(_08874_),
    .Y(_08880_));
 sky130_fd_sc_hd__nor2_8 _19148_ (.A(net319),
    .B(_04331_),
    .Y(_08881_));
 sky130_fd_sc_hd__or3_4 _19149_ (.A(net44),
    .B(net319),
    .C(_03286_),
    .X(_08882_));
 sky130_fd_sc_hd__o21ai_4 _19150_ (.A1(net160),
    .A2(_08666_),
    .B1(_04484_),
    .Y(_08883_));
 sky130_fd_sc_hd__o221a_1 _19151_ (.A1(_04277_),
    .A2(_04331_),
    .B1(_08879_),
    .B2(_08880_),
    .C1(_08883_),
    .X(_08884_));
 sky130_fd_sc_hd__o221ai_4 _19152_ (.A1(_04277_),
    .A2(_04331_),
    .B1(_08879_),
    .B2(_08880_),
    .C1(_08883_),
    .Y(_08885_));
 sky130_fd_sc_hd__a22oi_4 _19153_ (.A1(_08878_),
    .A2(_08873_),
    .B1(_08883_),
    .B2(_08882_),
    .Y(_08887_));
 sky130_fd_sc_hd__o2bb2ai_4 _19154_ (.A1_N(_08882_),
    .A2_N(_08883_),
    .B1(_08874_),
    .B2(_08877_),
    .Y(_08888_));
 sky130_fd_sc_hd__nand4_4 _19155_ (.A(_08675_),
    .B(_08872_),
    .C(_08885_),
    .D(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__a22oi_4 _19156_ (.A1(_08675_),
    .A2(_08872_),
    .B1(_08885_),
    .B2(_08888_),
    .Y(_08890_));
 sky130_fd_sc_hd__o2bb2ai_2 _19157_ (.A1_N(_08675_),
    .A2_N(_08872_),
    .B1(_08884_),
    .B2(_08887_),
    .Y(_08891_));
 sky130_fd_sc_hd__a2bb2oi_4 _19158_ (.A1_N(_08867_),
    .A2_N(_08870_),
    .B1(_08889_),
    .B2(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__a2bb2o_1 _19159_ (.A1_N(_08867_),
    .A2_N(_08870_),
    .B1(_08889_),
    .B2(_08891_),
    .X(_08893_));
 sky130_fd_sc_hd__o211ai_4 _19160_ (.A1(_08869_),
    .A2(_08861_),
    .B1(_08868_),
    .C1(_08889_),
    .Y(_08894_));
 sky130_fd_sc_hd__o2111a_1 _19161_ (.A1(_08869_),
    .A2(_08861_),
    .B1(_08868_),
    .C1(_08889_),
    .D1(_08891_),
    .X(_08895_));
 sky130_fd_sc_hd__o21a_2 _19162_ (.A1(_08892_),
    .A2(_08895_),
    .B1(_08852_),
    .X(_08896_));
 sky130_fd_sc_hd__o21ai_4 _19163_ (.A1(_08892_),
    .A2(_08895_),
    .B1(_08852_),
    .Y(_08898_));
 sky130_fd_sc_hd__o22ai_4 _19164_ (.A1(_08890_),
    .A2(_08894_),
    .B1(_08681_),
    .B2(_08684_),
    .Y(_08899_));
 sky130_fd_sc_hd__o221ai_4 _19165_ (.A1(_08681_),
    .A2(_08684_),
    .B1(_08890_),
    .B2(_08894_),
    .C1(_08893_),
    .Y(_08900_));
 sky130_fd_sc_hd__a21oi_2 _19166_ (.A1(_08611_),
    .A2(_08615_),
    .B1(_08613_),
    .Y(_08901_));
 sky130_fd_sc_hd__inv_2 _19167_ (.A(_08901_),
    .Y(_08902_));
 sky130_fd_sc_hd__o211ai_4 _19168_ (.A1(net175),
    .A2(_06759_),
    .B1(_05688_),
    .C1(net196),
    .Y(_08903_));
 sky130_fd_sc_hd__or3b_2 _19169_ (.A(net61),
    .B(_04201_),
    .C_N(net60),
    .X(_08904_));
 sky130_fd_sc_hd__a221oi_2 _19170_ (.A1(net205),
    .A2(_07073_),
    .B1(net171),
    .B2(net20),
    .C1(_05238_),
    .Y(_08905_));
 sky130_fd_sc_hd__nor2_1 _19171_ (.A(_04212_),
    .B(_05260_),
    .Y(_08906_));
 sky130_fd_sc_hd__a31oi_1 _19172_ (.A1(_07072_),
    .A2(net168),
    .A3(_05227_),
    .B1(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__o2bb2ai_4 _19173_ (.A1_N(_08903_),
    .A2_N(_08904_),
    .B1(_08905_),
    .B2(_08906_),
    .Y(_08909_));
 sky130_fd_sc_hd__nand3_2 _19174_ (.A(_08907_),
    .B(_08904_),
    .C(_08903_),
    .Y(_08910_));
 sky130_fd_sc_hd__a32o_1 _19175_ (.A1(net199),
    .A2(net172),
    .A3(net292),
    .B1(_06848_),
    .B2(net18),
    .X(_08911_));
 sky130_fd_sc_hd__a21oi_1 _19176_ (.A1(_08909_),
    .A2(_08910_),
    .B1(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__a21o_2 _19177_ (.A1(_08909_),
    .A2(_08910_),
    .B1(_08911_),
    .X(_08913_));
 sky130_fd_sc_hd__and3_2 _19178_ (.A(_08909_),
    .B(_08910_),
    .C(_08911_),
    .X(_08914_));
 sky130_fd_sc_hd__nand3_4 _19179_ (.A(_08909_),
    .B(_08910_),
    .C(_08911_),
    .Y(_08915_));
 sky130_fd_sc_hd__o22a_2 _19180_ (.A1(_08633_),
    .A2(_08635_),
    .B1(_08639_),
    .B2(_08642_),
    .X(_08916_));
 sky130_fd_sc_hd__o21ai_1 _19181_ (.A1(_08639_),
    .A2(_08642_),
    .B1(_08636_),
    .Y(_08917_));
 sky130_fd_sc_hd__o21ai_2 _19182_ (.A1(_08638_),
    .A2(_08641_),
    .B1(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__a21oi_4 _19183_ (.A1(_08913_),
    .A2(_08915_),
    .B1(_08918_),
    .Y(_08920_));
 sky130_fd_sc_hd__o21bai_4 _19184_ (.A1(_08912_),
    .A2(_08914_),
    .B1_N(_08918_),
    .Y(_08921_));
 sky130_fd_sc_hd__o21ai_4 _19185_ (.A1(_08643_),
    .A2(_08916_),
    .B1(_08913_),
    .Y(_08922_));
 sky130_fd_sc_hd__o211a_1 _19186_ (.A1(_08643_),
    .A2(_08916_),
    .B1(_08915_),
    .C1(_08913_),
    .X(_08923_));
 sky130_fd_sc_hd__o211ai_2 _19187_ (.A1(_08643_),
    .A2(_08916_),
    .B1(_08915_),
    .C1(_08913_),
    .Y(_08924_));
 sky130_fd_sc_hd__a21oi_4 _19188_ (.A1(_08921_),
    .A2(_08924_),
    .B1(_08902_),
    .Y(_08925_));
 sky130_fd_sc_hd__o21ai_2 _19189_ (.A1(_08920_),
    .A2(_08923_),
    .B1(_08901_),
    .Y(_08926_));
 sky130_fd_sc_hd__o211a_2 _19190_ (.A1(_08914_),
    .A2(_08922_),
    .B1(_08921_),
    .C1(_08902_),
    .X(_08927_));
 sky130_fd_sc_hd__o211ai_4 _19191_ (.A1(_08914_),
    .A2(_08922_),
    .B1(_08921_),
    .C1(_08902_),
    .Y(_08928_));
 sky130_fd_sc_hd__nand2_2 _19192_ (.A(_08926_),
    .B(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__a21o_1 _19193_ (.A1(_08898_),
    .A2(_08900_),
    .B1(_08929_),
    .X(_08931_));
 sky130_fd_sc_hd__o21ai_4 _19194_ (.A1(_08925_),
    .A2(_08927_),
    .B1(_08900_),
    .Y(_08932_));
 sky130_fd_sc_hd__o221ai_4 _19195_ (.A1(_08892_),
    .A2(_08899_),
    .B1(_08925_),
    .B2(_08927_),
    .C1(_08898_),
    .Y(_08933_));
 sky130_fd_sc_hd__o2bb2ai_1 _19196_ (.A1_N(_08898_),
    .A2_N(_08900_),
    .B1(_08925_),
    .B2(_08927_),
    .Y(_08934_));
 sky130_fd_sc_hd__o2111ai_4 _19197_ (.A1(_08892_),
    .A2(_08899_),
    .B1(_08926_),
    .C1(_08928_),
    .D1(_08898_),
    .Y(_08935_));
 sky130_fd_sc_hd__a21oi_4 _19198_ (.A1(_08630_),
    .A2(_08693_),
    .B1(_08690_),
    .Y(_08936_));
 sky130_fd_sc_hd__and3_1 _19199_ (.A(_08931_),
    .B(_08936_),
    .C(_08933_),
    .X(_08937_));
 sky130_fd_sc_hd__o211ai_4 _19200_ (.A1(_08896_),
    .A2(_08932_),
    .B1(_08936_),
    .C1(_08931_),
    .Y(_08938_));
 sky130_fd_sc_hd__a2bb2o_4 _19201_ (.A1_N(_08563_),
    .A2_N(_08558_),
    .B1(_08584_),
    .B2(_08566_),
    .X(_08939_));
 sky130_fd_sc_hd__o21ai_2 _19202_ (.A1(_08604_),
    .A2(_08619_),
    .B1(_08622_),
    .Y(_08940_));
 sky130_fd_sc_hd__o22a_2 _19203_ (.A1(_04091_),
    .A2(_01326_),
    .B1(_04793_),
    .B2(_01304_),
    .X(_08942_));
 sky130_fd_sc_hd__nor2_1 _19204_ (.A(_04113_),
    .B(_12363_),
    .Y(_08943_));
 sky130_fd_sc_hd__a31oi_4 _19205_ (.A1(net211),
    .A2(net183),
    .A3(_12330_),
    .B1(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__nand3_1 _19206_ (.A(net181),
    .B(net179),
    .C(net252),
    .Y(_08945_));
 sky130_fd_sc_hd__or3_1 _19207_ (.A(net35),
    .B(_04135_),
    .C(_03971_),
    .X(_08946_));
 sky130_fd_sc_hd__a21oi_1 _19208_ (.A1(_08945_),
    .A2(_08946_),
    .B1(_08944_),
    .Y(_08947_));
 sky130_fd_sc_hd__a21o_1 _19209_ (.A1(_08945_),
    .A2(_08946_),
    .B1(_08944_),
    .X(_08948_));
 sky130_fd_sc_hd__o211a_1 _19210_ (.A1(_04135_),
    .A2(_11804_),
    .B1(_08945_),
    .C1(_08944_),
    .X(_08949_));
 sky130_fd_sc_hd__o221ai_4 _19211_ (.A1(_04135_),
    .A2(_11804_),
    .B1(_05294_),
    .B2(_11782_),
    .C1(_08944_),
    .Y(_08950_));
 sky130_fd_sc_hd__o21a_1 _19212_ (.A1(_08947_),
    .A2(_08949_),
    .B1(_08942_),
    .X(_08951_));
 sky130_fd_sc_hd__nor3_2 _19213_ (.A(_08942_),
    .B(_08947_),
    .C(_08949_),
    .Y(_08953_));
 sky130_fd_sc_hd__a21oi_2 _19214_ (.A1(_08948_),
    .A2(_08950_),
    .B1(_08942_),
    .Y(_08954_));
 sky130_fd_sc_hd__a21o_1 _19215_ (.A1(_08948_),
    .A2(_08950_),
    .B1(_08942_),
    .X(_08955_));
 sky130_fd_sc_hd__and3_1 _19216_ (.A(_08948_),
    .B(_08950_),
    .C(_08942_),
    .X(_08956_));
 sky130_fd_sc_hd__nand3_1 _19217_ (.A(_08950_),
    .B(_08942_),
    .C(_08948_),
    .Y(_08957_));
 sky130_fd_sc_hd__o21a_1 _19218_ (.A1(_08549_),
    .A2(_08553_),
    .B1(_08545_),
    .X(_08958_));
 sky130_fd_sc_hd__o21ai_1 _19219_ (.A1(_08545_),
    .A2(_08555_),
    .B1(_08554_),
    .Y(_08959_));
 sky130_fd_sc_hd__a21boi_2 _19220_ (.A1(_08547_),
    .A2(_08556_),
    .B1_N(_08554_),
    .Y(_08960_));
 sky130_fd_sc_hd__o32a_4 _19221_ (.A1(_10324_),
    .A2(_05548_),
    .A3(net206),
    .B1(_10346_),
    .B2(_04146_),
    .X(_08961_));
 sky130_fd_sc_hd__o211ai_2 _19222_ (.A1(net231),
    .A2(_05927_),
    .B1(net291),
    .C1(_05933_),
    .Y(_08962_));
 sky130_fd_sc_hd__or3b_2 _19223_ (.A(net64),
    .B(_04157_),
    .C_N(net63),
    .X(_08964_));
 sky130_fd_sc_hd__o31a_1 _19224_ (.A1(_08261_),
    .A2(net205),
    .A3(_05932_),
    .B1(_08964_),
    .X(_08965_));
 sky130_fd_sc_hd__a32oi_4 _19225_ (.A1(net201),
    .A2(_06221_),
    .A3(_07658_),
    .B1(_07680_),
    .B2(net17),
    .Y(_08966_));
 sky130_fd_sc_hd__o211a_2 _19226_ (.A1(_04157_),
    .A2(_08283_),
    .B1(_08962_),
    .C1(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__nand2_2 _19227_ (.A(_08965_),
    .B(_08966_),
    .Y(_08968_));
 sky130_fd_sc_hd__a21oi_4 _19228_ (.A1(_08962_),
    .A2(_08964_),
    .B1(_08966_),
    .Y(_08969_));
 sky130_fd_sc_hd__o21a_1 _19229_ (.A1(_08965_),
    .A2(_08966_),
    .B1(_08961_),
    .X(_08970_));
 sky130_fd_sc_hd__o21ai_2 _19230_ (.A1(_08965_),
    .A2(_08966_),
    .B1(_08961_),
    .Y(_08971_));
 sky130_fd_sc_hd__o21bai_4 _19231_ (.A1(_08967_),
    .A2(_08969_),
    .B1_N(_08961_),
    .Y(_08972_));
 sky130_fd_sc_hd__nand3b_2 _19232_ (.A_N(_08969_),
    .B(_08961_),
    .C(_08968_),
    .Y(_08973_));
 sky130_fd_sc_hd__o21ai_1 _19233_ (.A1(_08967_),
    .A2(_08969_),
    .B1(_08961_),
    .Y(_08975_));
 sky130_fd_sc_hd__a21oi_4 _19234_ (.A1(_08972_),
    .A2(_08973_),
    .B1(_08960_),
    .Y(_08976_));
 sky130_fd_sc_hd__o311ai_4 _19235_ (.A1(_08961_),
    .A2(_08967_),
    .A3(_08969_),
    .B1(_08975_),
    .C1(_08959_),
    .Y(_08977_));
 sky130_fd_sc_hd__o211a_2 _19236_ (.A1(_08555_),
    .A2(_08958_),
    .B1(_08972_),
    .C1(_08973_),
    .X(_08978_));
 sky130_fd_sc_hd__o211ai_2 _19237_ (.A1(_08555_),
    .A2(_08958_),
    .B1(_08972_),
    .C1(_08973_),
    .Y(_08979_));
 sky130_fd_sc_hd__a32o_2 _19238_ (.A1(_08960_),
    .A2(_08972_),
    .A3(_08973_),
    .B1(_08957_),
    .B2(_08955_),
    .X(_08980_));
 sky130_fd_sc_hd__o211ai_2 _19239_ (.A1(_08954_),
    .A2(_08956_),
    .B1(_08977_),
    .C1(_08979_),
    .Y(_08981_));
 sky130_fd_sc_hd__inv_2 _19240_ (.A(_08981_),
    .Y(_08982_));
 sky130_fd_sc_hd__o22ai_4 _19241_ (.A1(_08951_),
    .A2(_08953_),
    .B1(_08976_),
    .B2(_08978_),
    .Y(_08983_));
 sky130_fd_sc_hd__o211ai_2 _19242_ (.A1(_08951_),
    .A2(_08953_),
    .B1(_08977_),
    .C1(_08979_),
    .Y(_08984_));
 sky130_fd_sc_hd__o22ai_2 _19243_ (.A1(_08954_),
    .A2(_08956_),
    .B1(_08976_),
    .B2(_08978_),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_1 _19244_ (.A(_08940_),
    .B(_08983_),
    .Y(_08987_));
 sky130_fd_sc_hd__and3_1 _19245_ (.A(_08940_),
    .B(_08981_),
    .C(_08983_),
    .X(_08988_));
 sky130_fd_sc_hd__o211ai_2 _19246_ (.A1(_08976_),
    .A2(_08980_),
    .B1(_08983_),
    .C1(_08940_),
    .Y(_08989_));
 sky130_fd_sc_hd__o2111a_1 _19247_ (.A1(_08604_),
    .A2(_08619_),
    .B1(_08622_),
    .C1(_08984_),
    .D1(_08986_),
    .X(_08990_));
 sky130_fd_sc_hd__o2111ai_4 _19248_ (.A1(_08604_),
    .A2(_08619_),
    .B1(_08622_),
    .C1(_08984_),
    .D1(_08986_),
    .Y(_08991_));
 sky130_fd_sc_hd__nor2_1 _19249_ (.A(_08939_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__a31oi_2 _19250_ (.A1(_08940_),
    .A2(_08981_),
    .A3(_08983_),
    .B1(_08939_),
    .Y(_08993_));
 sky130_fd_sc_hd__o2bb2ai_4 _19251_ (.A1_N(_08939_),
    .A2_N(_08991_),
    .B1(_08982_),
    .B2(_08987_),
    .Y(_08994_));
 sky130_fd_sc_hd__a21oi_2 _19252_ (.A1(_08989_),
    .A2(_08991_),
    .B1(_08939_),
    .Y(_08995_));
 sky130_fd_sc_hd__a21o_1 _19253_ (.A1(_08989_),
    .A2(_08991_),
    .B1(_08939_),
    .X(_08997_));
 sky130_fd_sc_hd__and3_1 _19254_ (.A(_08939_),
    .B(_08989_),
    .C(_08991_),
    .X(_08998_));
 sky130_fd_sc_hd__o211ai_2 _19255_ (.A1(_08982_),
    .A2(_08987_),
    .B1(_08991_),
    .C1(_08939_),
    .Y(_08999_));
 sky130_fd_sc_hd__nand2_2 _19256_ (.A(_08997_),
    .B(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__o2bb2ai_2 _19257_ (.A1_N(_08939_),
    .A2_N(_08988_),
    .B1(_08992_),
    .B2(_08994_),
    .Y(_09001_));
 sky130_fd_sc_hd__o211ai_4 _19258_ (.A1(_08690_),
    .A2(_08696_),
    .B1(_08934_),
    .C1(_08935_),
    .Y(_09002_));
 sky130_fd_sc_hd__o21ai_2 _19259_ (.A1(_08995_),
    .A2(_08998_),
    .B1(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__o211ai_4 _19260_ (.A1(_08995_),
    .A2(_08998_),
    .B1(_09002_),
    .C1(_08938_),
    .Y(_09004_));
 sky130_fd_sc_hd__a21o_2 _19261_ (.A1(_08938_),
    .A2(_09002_),
    .B1(_09000_),
    .X(_09005_));
 sky130_fd_sc_hd__a21oi_2 _19262_ (.A1(_08938_),
    .A2(_09002_),
    .B1(_09001_),
    .Y(_09006_));
 sky130_fd_sc_hd__a22o_1 _19263_ (.A1(_08997_),
    .A2(_08999_),
    .B1(_09002_),
    .B2(_08938_),
    .X(_09008_));
 sky130_fd_sc_hd__nand4_2 _19264_ (.A(_08938_),
    .B(_08997_),
    .C(_08999_),
    .D(_09002_),
    .Y(_09009_));
 sky130_fd_sc_hd__a32oi_4 _19265_ (.A1(_08603_),
    .A2(_08697_),
    .A3(_08698_),
    .B1(_08597_),
    .B2(_08596_),
    .Y(_09010_));
 sky130_fd_sc_hd__a21o_2 _19266_ (.A1(_08600_),
    .A2(_08701_),
    .B1(_08702_),
    .X(_09011_));
 sky130_fd_sc_hd__a21boi_1 _19267_ (.A1(_08600_),
    .A2(_08701_),
    .B1_N(_08703_),
    .Y(_09012_));
 sky130_fd_sc_hd__o221ai_4 _19268_ (.A1(_09003_),
    .A2(_08937_),
    .B1(_08702_),
    .B2(_09010_),
    .C1(_09005_),
    .Y(_09013_));
 sky130_fd_sc_hd__o21ai_2 _19269_ (.A1(_08699_),
    .A2(_08706_),
    .B1(_09009_),
    .Y(_09014_));
 sky130_fd_sc_hd__a21oi_2 _19270_ (.A1(_09004_),
    .A2(_09005_),
    .B1(_09011_),
    .Y(_09015_));
 sky130_fd_sc_hd__nand3_4 _19271_ (.A(_09008_),
    .B(_09009_),
    .C(_09012_),
    .Y(_09016_));
 sky130_fd_sc_hd__o21ai_2 _19272_ (.A1(_08456_),
    .A2(_08475_),
    .B1(_08474_),
    .Y(_09017_));
 sky130_fd_sc_hd__o21a_1 _19273_ (.A1(_08456_),
    .A2(_08475_),
    .B1(_08474_),
    .X(_09019_));
 sky130_fd_sc_hd__a21oi_1 _19274_ (.A1(_08460_),
    .A2(_08468_),
    .B1(_08465_),
    .Y(_09020_));
 sky130_fd_sc_hd__a21o_1 _19275_ (.A1(_08460_),
    .A2(_08468_),
    .B1(_08465_),
    .X(_09021_));
 sky130_fd_sc_hd__nor2_1 _19276_ (.A(_04059_),
    .B(_04218_),
    .Y(_09022_));
 sky130_fd_sc_hd__and3_1 _19277_ (.A(net230),
    .B(net228),
    .C(net281),
    .X(_09023_));
 sky130_fd_sc_hd__a31oi_4 _19278_ (.A1(net230),
    .A2(net228),
    .A3(net281),
    .B1(_09022_),
    .Y(_09024_));
 sky130_fd_sc_hd__o31ai_1 _19279_ (.A1(net259),
    .A2(_03956_),
    .A3(_04407_),
    .B1(net285),
    .Y(_09025_));
 sky130_fd_sc_hd__o32a_1 _19280_ (.A1(_04037_),
    .A2(net39),
    .A3(_04069_),
    .B1(_04410_),
    .B2(_09025_),
    .X(_09026_));
 sky130_fd_sc_hd__o22ai_2 _19281_ (.A1(_04069_),
    .A2(_03737_),
    .B1(_04410_),
    .B2(_09025_),
    .Y(_09027_));
 sky130_fd_sc_hd__or3b_1 _19282_ (.A(net38),
    .B(_04080_),
    .C_N(net37),
    .X(_09028_));
 sky130_fd_sc_hd__o31ai_1 _19283_ (.A1(_04557_),
    .A2(net7),
    .A3(net248),
    .B1(_02858_),
    .Y(_09030_));
 sky130_fd_sc_hd__o211ai_2 _19284_ (.A1(net231),
    .A2(_04557_),
    .B1(_02858_),
    .C1(net218),
    .Y(_09031_));
 sky130_fd_sc_hd__o22ai_2 _19285_ (.A1(_04080_),
    .A2(_02891_),
    .B1(_04554_),
    .B2(_09030_),
    .Y(_09032_));
 sky130_fd_sc_hd__o221a_2 _19286_ (.A1(_04080_),
    .A2(_02891_),
    .B1(_04562_),
    .B2(_02869_),
    .C1(_09026_),
    .X(_09033_));
 sky130_fd_sc_hd__nand2_2 _19287_ (.A(_09027_),
    .B(_09032_),
    .Y(_09034_));
 sky130_fd_sc_hd__o2111ai_1 _19288_ (.A1(_04080_),
    .A2(_02891_),
    .B1(_09024_),
    .C1(_09031_),
    .D1(_09026_),
    .Y(_09035_));
 sky130_fd_sc_hd__o221a_2 _19289_ (.A1(_04133_),
    .A2(_04216_),
    .B1(_04218_),
    .B2(_04059_),
    .C1(_09034_),
    .X(_09036_));
 sky130_fd_sc_hd__o22ai_1 _19290_ (.A1(_09022_),
    .A2(_09023_),
    .B1(_09027_),
    .B2(_09032_),
    .Y(_09037_));
 sky130_fd_sc_hd__o21ai_1 _19291_ (.A1(_09024_),
    .A2(_09033_),
    .B1(_09034_),
    .Y(_09038_));
 sky130_fd_sc_hd__a31o_1 _19292_ (.A1(_09026_),
    .A2(_09028_),
    .A3(_09031_),
    .B1(_09036_),
    .X(_09039_));
 sky130_fd_sc_hd__nand3_2 _19293_ (.A(_09034_),
    .B(_09035_),
    .C(_09037_),
    .Y(_09041_));
 sky130_fd_sc_hd__a211o_1 _19294_ (.A1(_09028_),
    .A2(_09031_),
    .B1(_09024_),
    .C1(_09026_),
    .X(_09042_));
 sky130_fd_sc_hd__o211a_1 _19295_ (.A1(_09024_),
    .A2(_09034_),
    .B1(_09041_),
    .C1(_08577_),
    .X(_09043_));
 sky130_fd_sc_hd__o211ai_2 _19296_ (.A1(_09024_),
    .A2(_09034_),
    .B1(_09041_),
    .C1(_08577_),
    .Y(_09044_));
 sky130_fd_sc_hd__a21oi_4 _19297_ (.A1(_09041_),
    .A2(_09042_),
    .B1(_08577_),
    .Y(_09045_));
 sky130_fd_sc_hd__o22ai_2 _19298_ (.A1(_08465_),
    .A2(_08471_),
    .B1(_09043_),
    .B2(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__nand3b_1 _19299_ (.A_N(_09045_),
    .B(_09020_),
    .C(_09044_),
    .Y(_09047_));
 sky130_fd_sc_hd__o21ai_1 _19300_ (.A1(_09043_),
    .A2(_09045_),
    .B1(_09020_),
    .Y(_09048_));
 sky130_fd_sc_hd__o21a_1 _19301_ (.A1(_08465_),
    .A2(_08471_),
    .B1(_09044_),
    .X(_09049_));
 sky130_fd_sc_hd__a31o_1 _19302_ (.A1(_08577_),
    .A2(_09041_),
    .A3(_09042_),
    .B1(_09020_),
    .X(_09050_));
 sky130_fd_sc_hd__nand3_4 _19303_ (.A(_09019_),
    .B(_09046_),
    .C(_09047_),
    .Y(_09052_));
 sky130_fd_sc_hd__inv_2 _19304_ (.A(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__o211ai_4 _19305_ (.A1(_09045_),
    .A2(_09050_),
    .B1(_09017_),
    .C1(_09048_),
    .Y(_09054_));
 sky130_fd_sc_hd__or3b_1 _19306_ (.A(_04026_),
    .B(net42),
    .C_N(net41),
    .X(_09055_));
 sky130_fd_sc_hd__nand2_1 _19307_ (.A(_02453_),
    .B(net279),
    .Y(_09056_));
 sky130_fd_sc_hd__nand3_1 _19308_ (.A(_02421_),
    .B(_02453_),
    .C(net279),
    .Y(_09057_));
 sky130_fd_sc_hd__o22ai_1 _19309_ (.A1(_04026_),
    .A2(_04483_),
    .B1(_02410_),
    .B2(_09056_),
    .Y(_09058_));
 sky130_fd_sc_hd__o211ai_2 _19310_ (.A1(net253),
    .A2(_03954_),
    .B1(net280),
    .C1(_03952_),
    .Y(_09059_));
 sky130_fd_sc_hd__nor2_1 _19311_ (.A(_04048_),
    .B(_04270_),
    .Y(_09060_));
 sky130_fd_sc_hd__or3b_2 _19312_ (.A(_04048_),
    .B(net41),
    .C_N(net40),
    .X(_09061_));
 sky130_fd_sc_hd__a22oi_2 _19313_ (.A1(_09055_),
    .A2(_09057_),
    .B1(_09059_),
    .B2(_09061_),
    .Y(_09063_));
 sky130_fd_sc_hd__a22o_2 _19314_ (.A1(_09055_),
    .A2(_09057_),
    .B1(_09059_),
    .B2(_09061_),
    .X(_09064_));
 sky130_fd_sc_hd__a211oi_1 _19315_ (.A1(_03959_),
    .A2(net280),
    .B1(_09060_),
    .C1(_09058_),
    .Y(_09065_));
 sky130_fd_sc_hd__nand3b_2 _19316_ (.A_N(_09058_),
    .B(_09059_),
    .C(_09061_),
    .Y(_09066_));
 sky130_fd_sc_hd__a32o_1 _19317_ (.A1(_00625_),
    .A2(net250),
    .A3(net243),
    .B1(_04897_),
    .B2(net5),
    .X(_09067_));
 sky130_fd_sc_hd__o21bai_2 _19318_ (.A1(_09063_),
    .A2(_09065_),
    .B1_N(_09067_),
    .Y(_09068_));
 sky130_fd_sc_hd__nand3_4 _19319_ (.A(_09064_),
    .B(_09066_),
    .C(_09067_),
    .Y(_09069_));
 sky130_fd_sc_hd__o21ai_4 _19320_ (.A1(_08486_),
    .A2(_08495_),
    .B1(_08494_),
    .Y(_09070_));
 sky130_fd_sc_hd__a21oi_2 _19321_ (.A1(_09068_),
    .A2(_09069_),
    .B1(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__a21o_1 _19322_ (.A1(_09068_),
    .A2(_09069_),
    .B1(_09070_),
    .X(_09072_));
 sky130_fd_sc_hd__nand3_4 _19323_ (.A(_09068_),
    .B(_09070_),
    .C(_09069_),
    .Y(_09074_));
 sky130_fd_sc_hd__nand2_1 _19324_ (.A(_09072_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__a32o_1 _19325_ (.A1(net255),
    .A2(_09698_),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net2),
    .X(_09076_));
 sky130_fd_sc_hd__and3_1 _19326_ (.A(_04124_),
    .B(net43),
    .C(net4),
    .X(_09077_));
 sky130_fd_sc_hd__a31oi_2 _19327_ (.A1(net234),
    .A2(net251),
    .A3(_04985_),
    .B1(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__a31o_1 _19328_ (.A1(net234),
    .A2(net251),
    .A3(_04985_),
    .B1(_09077_),
    .X(_09079_));
 sky130_fd_sc_hd__o32a_1 _19329_ (.A1(_05226_),
    .A2(_11420_),
    .A3(_11343_),
    .B1(_03982_),
    .B2(_05229_),
    .X(_09080_));
 sky130_fd_sc_hd__a32o_1 _19330_ (.A1(_11354_),
    .A2(net253),
    .A3(net276),
    .B1(_05228_),
    .B2(net3),
    .X(_09081_));
 sky130_fd_sc_hd__nand2_1 _19331_ (.A(_09079_),
    .B(_09081_),
    .Y(_09082_));
 sky130_fd_sc_hd__o221a_1 _19332_ (.A1(_11453_),
    .A2(_05226_),
    .B1(_05229_),
    .B2(_03982_),
    .C1(_09078_),
    .X(_09083_));
 sky130_fd_sc_hd__nand2_1 _19333_ (.A(_09078_),
    .B(_09080_),
    .Y(_09085_));
 sky130_fd_sc_hd__a21oi_1 _19334_ (.A1(_09082_),
    .A2(_09085_),
    .B1(_09076_),
    .Y(_09086_));
 sky130_fd_sc_hd__a21o_1 _19335_ (.A1(_09082_),
    .A2(_09085_),
    .B1(_09076_),
    .X(_09087_));
 sky130_fd_sc_hd__and3_1 _19336_ (.A(_09076_),
    .B(_09082_),
    .C(_09085_),
    .X(_09088_));
 sky130_fd_sc_hd__nand3_1 _19337_ (.A(_09076_),
    .B(_09082_),
    .C(_09085_),
    .Y(_09089_));
 sky130_fd_sc_hd__nand2_1 _19338_ (.A(_09087_),
    .B(_09089_),
    .Y(_09090_));
 sky130_fd_sc_hd__and4_1 _19339_ (.A(_09072_),
    .B(_09074_),
    .C(_09087_),
    .D(_09089_),
    .X(_09091_));
 sky130_fd_sc_hd__o2bb2a_1 _19340_ (.A1_N(_09072_),
    .A2_N(_09074_),
    .B1(_09086_),
    .B2(_09088_),
    .X(_09092_));
 sky130_fd_sc_hd__and3_1 _19341_ (.A(_09075_),
    .B(_09087_),
    .C(_09089_),
    .X(_09093_));
 sky130_fd_sc_hd__a211o_1 _19342_ (.A1(_09072_),
    .A2(_09074_),
    .B1(_09086_),
    .C1(_09088_),
    .X(_09094_));
 sky130_fd_sc_hd__and3_1 _19343_ (.A(_09072_),
    .B(_09074_),
    .C(_09090_),
    .X(_09096_));
 sky130_fd_sc_hd__a21o_1 _19344_ (.A1(_09087_),
    .A2(_09089_),
    .B1(_09075_),
    .X(_09097_));
 sky130_fd_sc_hd__o2bb2a_1 _19345_ (.A1_N(_09052_),
    .A2_N(_09054_),
    .B1(_09091_),
    .B2(_09092_),
    .X(_09098_));
 sky130_fd_sc_hd__o2bb2ai_2 _19346_ (.A1_N(_09052_),
    .A2_N(_09054_),
    .B1(_09091_),
    .B2(_09092_),
    .Y(_09099_));
 sky130_fd_sc_hd__o211ai_4 _19347_ (.A1(_09093_),
    .A2(_09096_),
    .B1(_09052_),
    .C1(_09054_),
    .Y(_09100_));
 sky130_fd_sc_hd__o2bb2ai_2 _19348_ (.A1_N(_09052_),
    .A2_N(_09054_),
    .B1(_09093_),
    .B2(_09096_),
    .Y(_09101_));
 sky130_fd_sc_hd__o211ai_4 _19349_ (.A1(_09091_),
    .A2(_09092_),
    .B1(_09052_),
    .C1(_09054_),
    .Y(_09102_));
 sky130_fd_sc_hd__nand4_4 _19350_ (.A(_08592_),
    .B(_08595_),
    .C(_09101_),
    .D(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__o21ai_1 _19351_ (.A1(_08591_),
    .A2(_08594_),
    .B1(_09100_),
    .Y(_09104_));
 sky130_fd_sc_hd__o211a_1 _19352_ (.A1(_08591_),
    .A2(_08594_),
    .B1(_09099_),
    .C1(_09100_),
    .X(_09105_));
 sky130_fd_sc_hd__o211ai_4 _19353_ (.A1(_08591_),
    .A2(_08594_),
    .B1(_09099_),
    .C1(_09100_),
    .Y(_09107_));
 sky130_fd_sc_hd__a31o_2 _19354_ (.A1(_08482_),
    .A2(_08517_),
    .A3(_08518_),
    .B1(_08483_),
    .X(_09108_));
 sky130_fd_sc_hd__o2bb2a_2 _19355_ (.A1_N(_08477_),
    .A2_N(_08479_),
    .B1(_08519_),
    .B2(_08481_),
    .X(_09109_));
 sky130_fd_sc_hd__a21oi_2 _19356_ (.A1(_09103_),
    .A2(_09107_),
    .B1(_09109_),
    .Y(_09110_));
 sky130_fd_sc_hd__and3_1 _19357_ (.A(_09103_),
    .B(_09107_),
    .C(_09109_),
    .X(_09111_));
 sky130_fd_sc_hd__a21oi_2 _19358_ (.A1(_09103_),
    .A2(_09107_),
    .B1(_09108_),
    .Y(_09112_));
 sky130_fd_sc_hd__a21o_1 _19359_ (.A1(_09103_),
    .A2(_09107_),
    .B1(_09108_),
    .X(_09113_));
 sky130_fd_sc_hd__a41oi_4 _19360_ (.A1(_08592_),
    .A2(_08595_),
    .A3(_09101_),
    .A4(_09102_),
    .B1(_09109_),
    .Y(_09114_));
 sky130_fd_sc_hd__nand2_1 _19361_ (.A(_09103_),
    .B(_09108_),
    .Y(_09115_));
 sky130_fd_sc_hd__and3_1 _19362_ (.A(_09103_),
    .B(_09107_),
    .C(_09108_),
    .X(_09116_));
 sky130_fd_sc_hd__o21ai_2 _19363_ (.A1(_09105_),
    .A2(_09115_),
    .B1(_09113_),
    .Y(_09118_));
 sky130_fd_sc_hd__a21oi_1 _19364_ (.A1(_09107_),
    .A2(_09114_),
    .B1(_09112_),
    .Y(_09119_));
 sky130_fd_sc_hd__o221ai_4 _19365_ (.A1(_09112_),
    .A2(_09116_),
    .B1(_09006_),
    .B2(_09014_),
    .C1(_09013_),
    .Y(_09120_));
 sky130_fd_sc_hd__o2bb2ai_2 _19366_ (.A1_N(_09013_),
    .A2_N(_09016_),
    .B1(_09110_),
    .B2(_09111_),
    .Y(_09121_));
 sky130_fd_sc_hd__o2bb2ai_2 _19367_ (.A1_N(_09013_),
    .A2_N(_09016_),
    .B1(_09112_),
    .B2(_09116_),
    .Y(_09122_));
 sky130_fd_sc_hd__a31oi_2 _19368_ (.A1(_09011_),
    .A2(_09005_),
    .A3(_09004_),
    .B1(_09118_),
    .Y(_09123_));
 sky130_fd_sc_hd__o21ai_1 _19369_ (.A1(_09110_),
    .A2(_09111_),
    .B1(_09013_),
    .Y(_09124_));
 sky130_fd_sc_hd__o211ai_4 _19370_ (.A1(_09110_),
    .A2(_09111_),
    .B1(_09013_),
    .C1(_09016_),
    .Y(_09125_));
 sky130_fd_sc_hd__a22oi_2 _19371_ (.A1(_08716_),
    .A2(_08849_),
    .B1(_09122_),
    .B2(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__o211ai_4 _19372_ (.A1(_08715_),
    .A2(_08848_),
    .B1(_09120_),
    .C1(_09121_),
    .Y(_09127_));
 sky130_fd_sc_hd__o211a_1 _19373_ (.A1(_09015_),
    .A2(_09124_),
    .B1(_08850_),
    .C1(_09122_),
    .X(_09129_));
 sky130_fd_sc_hd__nand3_4 _19374_ (.A(_09122_),
    .B(_09125_),
    .C(_08850_),
    .Y(_09130_));
 sky130_fd_sc_hd__o211ai_2 _19375_ (.A1(_08843_),
    .A2(_08845_),
    .B1(_09127_),
    .C1(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__a21o_1 _19376_ (.A1(_09127_),
    .A2(_09130_),
    .B1(_08847_),
    .X(_09132_));
 sky130_fd_sc_hd__o21ai_2 _19377_ (.A1(_08843_),
    .A2(_08845_),
    .B1(_09130_),
    .Y(_09133_));
 sky130_fd_sc_hd__a32oi_4 _19378_ (.A1(_08851_),
    .A2(_09120_),
    .A3(_09121_),
    .B1(_09130_),
    .B2(_08847_),
    .Y(_09134_));
 sky130_fd_sc_hd__nand4_2 _19379_ (.A(_08844_),
    .B(_08846_),
    .C(_09127_),
    .D(_09130_),
    .Y(_09135_));
 sky130_fd_sc_hd__inv_2 _19380_ (.A(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__o22ai_2 _19381_ (.A1(_08843_),
    .A2(_08845_),
    .B1(_09126_),
    .B2(_09129_),
    .Y(_09137_));
 sky130_fd_sc_hd__o21ai_1 _19382_ (.A1(_08721_),
    .A2(_08728_),
    .B1(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__a2bb2oi_2 _19383_ (.A1_N(_08721_),
    .A2_N(_08728_),
    .B1(_09131_),
    .B2(_09132_),
    .Y(_09140_));
 sky130_fd_sc_hd__o211ai_2 _19384_ (.A1(_08721_),
    .A2(_08728_),
    .B1(_09135_),
    .C1(_09137_),
    .Y(_09141_));
 sky130_fd_sc_hd__a21oi_1 _19385_ (.A1(_09135_),
    .A2(_09137_),
    .B1(_08760_),
    .Y(_09142_));
 sky130_fd_sc_hd__nand3_2 _19386_ (.A(_08759_),
    .B(_09131_),
    .C(_09132_),
    .Y(_09143_));
 sky130_fd_sc_hd__o22ai_2 _19387_ (.A1(_08435_),
    .A2(_08441_),
    .B1(_09140_),
    .B2(_09142_),
    .Y(_09144_));
 sky130_fd_sc_hd__o2111ai_4 _19388_ (.A1(_08364_),
    .A2(_08431_),
    .B1(_08442_),
    .C1(_09141_),
    .D1(_09143_),
    .Y(_09145_));
 sky130_fd_sc_hd__o22ai_1 _19389_ (.A1(_08432_),
    .A2(_08757_),
    .B1(_09140_),
    .B2(_09142_),
    .Y(_09146_));
 sky130_fd_sc_hd__o211ai_1 _19390_ (.A1(_08435_),
    .A2(_08441_),
    .B1(_09141_),
    .C1(_09143_),
    .Y(_09147_));
 sky130_fd_sc_hd__a21oi_1 _19391_ (.A1(_09146_),
    .A2(_09147_),
    .B1(_08755_),
    .Y(_09148_));
 sky130_fd_sc_hd__nand3_1 _19392_ (.A(_08756_),
    .B(_09144_),
    .C(_09145_),
    .Y(_09149_));
 sky130_fd_sc_hd__a21oi_1 _19393_ (.A1(_09144_),
    .A2(_09145_),
    .B1(_08756_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand3_1 _19394_ (.A(_09146_),
    .B(_09147_),
    .C(_08755_),
    .Y(_09152_));
 sky130_fd_sc_hd__nor2_1 _19395_ (.A(_08399_),
    .B(_08421_),
    .Y(_09153_));
 sky130_fd_sc_hd__a21oi_1 _19396_ (.A1(_08399_),
    .A2(_08422_),
    .B1(_08421_),
    .Y(_09154_));
 sky130_fd_sc_hd__a31oi_1 _19397_ (.A1(_08756_),
    .A2(_09144_),
    .A3(_09145_),
    .B1(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__nand3b_1 _19398_ (.A_N(_09154_),
    .B(_09152_),
    .C(_09149_),
    .Y(_09156_));
 sky130_fd_sc_hd__o2bb2ai_1 _19399_ (.A1_N(_09149_),
    .A2_N(_09152_),
    .B1(_09153_),
    .B2(_08423_),
    .Y(_09157_));
 sky130_fd_sc_hd__o21a_1 _19400_ (.A1(_07654_),
    .A2(_08028_),
    .B1(_08741_),
    .X(_09158_));
 sky130_fd_sc_hd__o2bb2ai_1 _19401_ (.A1_N(_09156_),
    .A2_N(_09157_),
    .B1(_09158_),
    .B2(_08742_),
    .Y(_09159_));
 sky130_fd_sc_hd__o211ai_2 _19402_ (.A1(_08740_),
    .A2(_08745_),
    .B1(_09156_),
    .C1(_09157_),
    .Y(_09160_));
 sky130_fd_sc_hd__nand2_1 _19403_ (.A(_09159_),
    .B(_09160_),
    .Y(_09162_));
 sky130_fd_sc_hd__o2111a_2 _19404_ (.A1(_08746_),
    .A2(_08750_),
    .B1(_08353_),
    .C1(_08749_),
    .D1(_07959_),
    .X(_09163_));
 sky130_fd_sc_hd__nand4_1 _19405_ (.A(_08749_),
    .B(_08751_),
    .C(_08353_),
    .D(_08354_),
    .Y(_09164_));
 sky130_fd_sc_hd__o211ai_1 _19406_ (.A1(_08346_),
    .A2(_08351_),
    .B1(_08747_),
    .C1(_08748_),
    .Y(_09165_));
 sky130_fd_sc_hd__nand2_1 _19407_ (.A(_09164_),
    .B(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__a21oi_4 _19408_ (.A1(_09163_),
    .A2(_07598_),
    .B1(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__nand2_1 _19409_ (.A(_07599_),
    .B(_09163_),
    .Y(_09168_));
 sky130_fd_sc_hd__o211ai_4 _19410_ (.A1(_06315_),
    .A2(_06318_),
    .B1(_07599_),
    .C1(_09163_),
    .Y(_09169_));
 sky130_fd_sc_hd__o21a_2 _19411_ (.A1(_06319_),
    .A2(_09168_),
    .B1(_09167_),
    .X(_09170_));
 sky130_fd_sc_hd__o21ai_4 _19412_ (.A1(_06319_),
    .A2(_09168_),
    .B1(_09167_),
    .Y(_09171_));
 sky130_fd_sc_hd__xnor2_1 _19413_ (.A(_09162_),
    .B(_09171_),
    .Y(net90));
 sky130_fd_sc_hd__o2bb2ai_1 _19414_ (.A1_N(_08758_),
    .A2_N(_09143_),
    .B1(_09138_),
    .B2(_09136_),
    .Y(_09173_));
 sky130_fd_sc_hd__a21oi_2 _19415_ (.A1(_09143_),
    .A2(_08758_),
    .B1(_09140_),
    .Y(_09174_));
 sky130_fd_sc_hd__a32oi_4 _19416_ (.A1(_09004_),
    .A2(_09005_),
    .A3(_09011_),
    .B1(_09016_),
    .B2(_09118_),
    .Y(_09175_));
 sky130_fd_sc_hd__a2bb2oi_2 _19417_ (.A1_N(_09006_),
    .A2_N(_09014_),
    .B1(_09119_),
    .B2(_09013_),
    .Y(_09176_));
 sky130_fd_sc_hd__a21oi_1 _19418_ (.A1(_09066_),
    .A2(_09067_),
    .B1(_09063_),
    .Y(_09177_));
 sky130_fd_sc_hd__and3_1 _19419_ (.A(_04102_),
    .B(net42),
    .C(net6),
    .X(_09178_));
 sky130_fd_sc_hd__o311a_1 _19420_ (.A1(net259),
    .A2(_11387_),
    .A3(_02442_),
    .B1(net243),
    .C1(_02421_),
    .X(_09179_));
 sky130_fd_sc_hd__a31oi_4 _19421_ (.A1(_02421_),
    .A2(net248),
    .A3(net243),
    .B1(_09178_),
    .Y(_09180_));
 sky130_fd_sc_hd__nor2_1 _19422_ (.A(_04059_),
    .B(_04270_),
    .Y(_09181_));
 sky130_fd_sc_hd__a31oi_4 _19423_ (.A1(net230),
    .A2(net228),
    .A3(net280),
    .B1(_09181_),
    .Y(_09183_));
 sky130_fd_sc_hd__a311o_1 _19424_ (.A1(_06519_),
    .A2(net286),
    .A3(net283),
    .B1(_04481_),
    .C1(_03951_),
    .X(_09184_));
 sky130_fd_sc_hd__or3b_2 _19425_ (.A(_04048_),
    .B(net42),
    .C_N(net41),
    .X(_09185_));
 sky130_fd_sc_hd__a32oi_4 _19426_ (.A1(_03952_),
    .A2(net231),
    .A3(net279),
    .B1(_04482_),
    .B2(net7),
    .Y(_09186_));
 sky130_fd_sc_hd__a21oi_2 _19427_ (.A1(_09184_),
    .A2(_09185_),
    .B1(_09183_),
    .Y(_09187_));
 sky130_fd_sc_hd__a21o_1 _19428_ (.A1(_09184_),
    .A2(_09185_),
    .B1(_09183_),
    .X(_09188_));
 sky130_fd_sc_hd__o2111ai_4 _19429_ (.A1(_03961_),
    .A2(_04481_),
    .B1(_09180_),
    .C1(_09185_),
    .D1(_09183_),
    .Y(_09189_));
 sky130_fd_sc_hd__o2bb2a_1 _19430_ (.A1_N(_09183_),
    .A2_N(_09186_),
    .B1(_09178_),
    .B2(_09179_),
    .X(_09190_));
 sky130_fd_sc_hd__o2bb2ai_2 _19431_ (.A1_N(_09183_),
    .A2_N(_09186_),
    .B1(_09178_),
    .B2(_09179_),
    .Y(_09191_));
 sky130_fd_sc_hd__o211ai_4 _19432_ (.A1(_09183_),
    .A2(_09186_),
    .B1(_09189_),
    .C1(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__a211o_1 _19433_ (.A1(_09184_),
    .A2(_09185_),
    .B1(_09180_),
    .C1(_09183_),
    .X(_09194_));
 sky130_fd_sc_hd__a22oi_4 _19434_ (.A1(_09064_),
    .A2(_09069_),
    .B1(_09192_),
    .B2(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__o211a_1 _19435_ (.A1(_09180_),
    .A2(_09188_),
    .B1(_09177_),
    .C1(_09192_),
    .X(_09196_));
 sky130_fd_sc_hd__o211ai_2 _19436_ (.A1(_09180_),
    .A2(_09188_),
    .B1(_09177_),
    .C1(_09192_),
    .Y(_09197_));
 sky130_fd_sc_hd__o32a_1 _19437_ (.A1(_05463_),
    .A2(_11420_),
    .A3(_11343_),
    .B1(_03982_),
    .B2(_05465_),
    .X(_09198_));
 sky130_fd_sc_hd__a32o_1 _19438_ (.A1(_11354_),
    .A2(net253),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net3),
    .X(_09199_));
 sky130_fd_sc_hd__a41oi_4 _19439_ (.A1(net307),
    .A2(net296),
    .A3(net287),
    .A4(_00635_),
    .B1(_04986_),
    .Y(_09200_));
 sky130_fd_sc_hd__a22oi_2 _19440_ (.A1(net5),
    .A2(_04988_),
    .B1(_00625_),
    .B2(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__a32oi_2 _19441_ (.A1(net234),
    .A2(net251),
    .A3(net276),
    .B1(_05228_),
    .B2(net4),
    .Y(_09202_));
 sky130_fd_sc_hd__nor2_1 _19442_ (.A(_09201_),
    .B(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__o221a_1 _19443_ (.A1(_13021_),
    .A2(_05226_),
    .B1(_05229_),
    .B2(_04004_),
    .C1(_09201_),
    .X(_09205_));
 sky130_fd_sc_hd__nand2_1 _19444_ (.A(_09201_),
    .B(_09202_),
    .Y(_09206_));
 sky130_fd_sc_hd__o21ai_1 _19445_ (.A1(_09203_),
    .A2(_09205_),
    .B1(_09199_),
    .Y(_09207_));
 sky130_fd_sc_hd__nand3b_1 _19446_ (.A_N(_09203_),
    .B(_09206_),
    .C(_09198_),
    .Y(_09208_));
 sky130_fd_sc_hd__nand2_1 _19447_ (.A(_09207_),
    .B(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__o211ai_2 _19448_ (.A1(_09195_),
    .A2(_09196_),
    .B1(_09207_),
    .C1(_09208_),
    .Y(_09210_));
 sky130_fd_sc_hd__nand3b_1 _19449_ (.A_N(_09195_),
    .B(_09197_),
    .C(_09209_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand2_1 _19450_ (.A(_09210_),
    .B(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__nor2_1 _19451_ (.A(_04080_),
    .B(_03737_),
    .Y(_09213_));
 sky130_fd_sc_hd__a31o_1 _19452_ (.A1(_11420_),
    .A2(net283),
    .A3(_04556_),
    .B1(_03714_),
    .X(_09214_));
 sky130_fd_sc_hd__nor3_1 _19453_ (.A(net216),
    .B(_03714_),
    .C(_04554_),
    .Y(_09216_));
 sky130_fd_sc_hd__o32a_1 _19454_ (.A1(_04037_),
    .A2(net39),
    .A3(_04080_),
    .B1(_04554_),
    .B2(_09214_),
    .X(_09217_));
 sky130_fd_sc_hd__o311a_1 _19455_ (.A1(net7),
    .A2(net248),
    .A3(_04787_),
    .B1(_02858_),
    .C1(net214),
    .X(_09218_));
 sky130_fd_sc_hd__and3_1 _19456_ (.A(_04037_),
    .B(net11),
    .C(net37),
    .X(_09219_));
 sky130_fd_sc_hd__or3b_1 _19457_ (.A(net38),
    .B(_04091_),
    .C_N(net37),
    .X(_09220_));
 sky130_fd_sc_hd__a31o_1 _19458_ (.A1(net214),
    .A2(_02858_),
    .A3(net184),
    .B1(_09219_),
    .X(_09221_));
 sky130_fd_sc_hd__o221ai_4 _19459_ (.A1(_04080_),
    .A2(_03737_),
    .B1(_04554_),
    .B2(_09214_),
    .C1(_09220_),
    .Y(_09222_));
 sky130_fd_sc_hd__o221ai_2 _19460_ (.A1(_04091_),
    .A2(_02891_),
    .B1(_04793_),
    .B2(_02869_),
    .C1(_09217_),
    .Y(_09223_));
 sky130_fd_sc_hd__o22a_2 _19461_ (.A1(_09213_),
    .A2(_09216_),
    .B1(_09218_),
    .B2(_09219_),
    .X(_09224_));
 sky130_fd_sc_hd__o21ai_1 _19462_ (.A1(_09213_),
    .A2(_09216_),
    .B1(_09221_),
    .Y(_09225_));
 sky130_fd_sc_hd__o21ai_1 _19463_ (.A1(_09218_),
    .A2(_09222_),
    .B1(_09225_),
    .Y(_09227_));
 sky130_fd_sc_hd__o22a_1 _19464_ (.A1(_04069_),
    .A2(_04218_),
    .B1(net187),
    .B2(_04216_),
    .X(_09228_));
 sky130_fd_sc_hd__a32o_1 _19465_ (.A1(net222),
    .A2(net281),
    .A3(net188),
    .B1(_04217_),
    .B2(net9),
    .X(_09229_));
 sky130_fd_sc_hd__nand2_2 _19466_ (.A(_09227_),
    .B(_09228_),
    .Y(_09230_));
 sky130_fd_sc_hd__o21ai_1 _19467_ (.A1(_09218_),
    .A2(_09222_),
    .B1(_09229_),
    .Y(_09231_));
 sky130_fd_sc_hd__and3_4 _19468_ (.A(_09223_),
    .B(_09225_),
    .C(_09229_),
    .X(_09232_));
 sky130_fd_sc_hd__o211ai_2 _19469_ (.A1(_09222_),
    .A2(_09218_),
    .B1(_09229_),
    .C1(_09225_),
    .Y(_09233_));
 sky130_fd_sc_hd__o21ai_4 _19470_ (.A1(_08942_),
    .A2(_08949_),
    .B1(_08948_),
    .Y(_09234_));
 sky130_fd_sc_hd__a21oi_4 _19471_ (.A1(_09230_),
    .A2(_09233_),
    .B1(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__a21o_1 _19472_ (.A1(_09230_),
    .A2(_09233_),
    .B1(_09234_),
    .X(_09236_));
 sky130_fd_sc_hd__nand2_2 _19473_ (.A(_09230_),
    .B(_09234_),
    .Y(_09238_));
 sky130_fd_sc_hd__o211a_1 _19474_ (.A1(_09224_),
    .A2(_09231_),
    .B1(_09234_),
    .C1(_09230_),
    .X(_09239_));
 sky130_fd_sc_hd__o211ai_2 _19475_ (.A1(_09232_),
    .A2(_09238_),
    .B1(_09038_),
    .C1(_09236_),
    .Y(_09240_));
 sky130_fd_sc_hd__o22ai_2 _19476_ (.A1(_09033_),
    .A2(_09036_),
    .B1(_09235_),
    .B2(_09239_),
    .Y(_09241_));
 sky130_fd_sc_hd__o21ai_2 _19477_ (.A1(_09235_),
    .A2(_09239_),
    .B1(_09038_),
    .Y(_09242_));
 sky130_fd_sc_hd__o221ai_4 _19478_ (.A1(_09033_),
    .A2(_09036_),
    .B1(_09232_),
    .B2(_09238_),
    .C1(_09236_),
    .Y(_09243_));
 sky130_fd_sc_hd__a21oi_2 _19479_ (.A1(_09021_),
    .A2(_09044_),
    .B1(_09045_),
    .Y(_09244_));
 sky130_fd_sc_hd__and3_1 _19480_ (.A(_09242_),
    .B(_09243_),
    .C(_09244_),
    .X(_09245_));
 sky130_fd_sc_hd__nand3_1 _19481_ (.A(_09242_),
    .B(_09243_),
    .C(_09244_),
    .Y(_09246_));
 sky130_fd_sc_hd__o211a_1 _19482_ (.A1(_09045_),
    .A2(_09049_),
    .B1(_09240_),
    .C1(_09241_),
    .X(_09247_));
 sky130_fd_sc_hd__o211ai_4 _19483_ (.A1(_09045_),
    .A2(_09049_),
    .B1(_09240_),
    .C1(_09241_),
    .Y(_09249_));
 sky130_fd_sc_hd__nand3_1 _19484_ (.A(_09212_),
    .B(_09246_),
    .C(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__a21o_1 _19485_ (.A1(_09246_),
    .A2(_09249_),
    .B1(_09212_),
    .X(_09251_));
 sky130_fd_sc_hd__a22o_1 _19486_ (.A1(_09210_),
    .A2(_09211_),
    .B1(_09246_),
    .B2(_09249_),
    .X(_09252_));
 sky130_fd_sc_hd__a31oi_2 _19487_ (.A1(_09242_),
    .A2(_09243_),
    .A3(_09244_),
    .B1(_09212_),
    .Y(_09253_));
 sky130_fd_sc_hd__nand2_1 _19488_ (.A(_09253_),
    .B(_09249_),
    .Y(_09254_));
 sky130_fd_sc_hd__o211ai_4 _19489_ (.A1(_08990_),
    .A2(_08993_),
    .B1(_09250_),
    .C1(_09251_),
    .Y(_09255_));
 sky130_fd_sc_hd__nand3_4 _19490_ (.A(_09252_),
    .B(_09254_),
    .C(_08994_),
    .Y(_09256_));
 sky130_fd_sc_hd__and3_1 _19491_ (.A(_09054_),
    .B(_09094_),
    .C(_09097_),
    .X(_09257_));
 sky130_fd_sc_hd__a31oi_4 _19492_ (.A1(_09054_),
    .A2(_09094_),
    .A3(_09097_),
    .B1(_09053_),
    .Y(_09258_));
 sky130_fd_sc_hd__and3_2 _19493_ (.A(_09255_),
    .B(_09256_),
    .C(_09258_),
    .X(_09260_));
 sky130_fd_sc_hd__nand3_2 _19494_ (.A(_09255_),
    .B(_09256_),
    .C(_09258_),
    .Y(_09261_));
 sky130_fd_sc_hd__a21oi_2 _19495_ (.A1(_09255_),
    .A2(_09256_),
    .B1(_09258_),
    .Y(_09262_));
 sky130_fd_sc_hd__o2bb2ai_2 _19496_ (.A1_N(_09255_),
    .A2_N(_09256_),
    .B1(_09257_),
    .B2(_09053_),
    .Y(_09263_));
 sky130_fd_sc_hd__nand2_2 _19497_ (.A(_09261_),
    .B(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__a32oi_4 _19498_ (.A1(_08931_),
    .A2(_08933_),
    .A3(_08936_),
    .B1(_09000_),
    .B2(_09002_),
    .Y(_09265_));
 sky130_fd_sc_hd__a21boi_4 _19499_ (.A1(_08938_),
    .A2(_09001_),
    .B1_N(_09002_),
    .Y(_09266_));
 sky130_fd_sc_hd__o22ai_4 _19500_ (.A1(_08892_),
    .A2(_08899_),
    .B1(_08929_),
    .B2(_08896_),
    .Y(_09267_));
 sky130_fd_sc_hd__and3b_2 _19501_ (.A_N(net59),
    .B(net22),
    .C(net58),
    .X(_09268_));
 sky130_fd_sc_hd__o311a_2 _19502_ (.A1(_03958_),
    .A2(_05927_),
    .A3(_07767_),
    .B1(_07771_),
    .C1(_04889_),
    .X(_09269_));
 sky130_fd_sc_hd__a31o_1 _19503_ (.A1(_07771_),
    .A2(_04889_),
    .A3(_07769_),
    .B1(_09268_),
    .X(_09271_));
 sky130_fd_sc_hd__nor2_1 _19504_ (.A(_04277_),
    .B(_04375_),
    .Y(_09272_));
 sky130_fd_sc_hd__or3b_2 _19505_ (.A(net55),
    .B(_04277_),
    .C_N(net44),
    .X(_09273_));
 sky130_fd_sc_hd__a21oi_4 _19506_ (.A1(net151),
    .A2(net158),
    .B1(_04353_),
    .Y(_09274_));
 sky130_fd_sc_hd__o21ai_1 _19507_ (.A1(net160),
    .A2(_08666_),
    .B1(_04342_),
    .Y(_09275_));
 sky130_fd_sc_hd__o21ai_1 _19508_ (.A1(_07076_),
    .A2(_08206_),
    .B1(_04627_),
    .Y(_09276_));
 sky130_fd_sc_hd__a32oi_1 _19509_ (.A1(_08204_),
    .A2(net163),
    .A3(_04627_),
    .B1(_04649_),
    .B2(net24),
    .Y(_09277_));
 sky130_fd_sc_hd__a32o_1 _19510_ (.A1(_08204_),
    .A2(net163),
    .A3(_04627_),
    .B1(_04649_),
    .B2(net24),
    .X(_09278_));
 sky130_fd_sc_hd__o21ai_4 _19511_ (.A1(_09272_),
    .A2(_09274_),
    .B1(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__o221ai_4 _19512_ (.A1(_04256_),
    .A2(net316),
    .B1(_08203_),
    .B2(_09276_),
    .C1(_09273_),
    .Y(_09280_));
 sky130_fd_sc_hd__o211ai_2 _19513_ (.A1(_04277_),
    .A2(_04375_),
    .B1(_09277_),
    .C1(_09275_),
    .Y(_09282_));
 sky130_fd_sc_hd__o22ai_4 _19514_ (.A1(_09268_),
    .A2(_09269_),
    .B1(_09274_),
    .B2(_09280_),
    .Y(_09283_));
 sky130_fd_sc_hd__nand2_1 _19515_ (.A(_09279_),
    .B(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__a21oi_2 _19516_ (.A1(_09279_),
    .A2(_09282_),
    .B1(_09271_),
    .Y(_09285_));
 sky130_fd_sc_hd__a21o_1 _19517_ (.A1(_09279_),
    .A2(_09282_),
    .B1(_09271_),
    .X(_09286_));
 sky130_fd_sc_hd__o221a_2 _19518_ (.A1(_09268_),
    .A2(_09269_),
    .B1(_09274_),
    .B2(_09280_),
    .C1(_09279_),
    .X(_09287_));
 sky130_fd_sc_hd__o221ai_4 _19519_ (.A1(_09268_),
    .A2(_09269_),
    .B1(_09274_),
    .B2(_09280_),
    .C1(_09279_),
    .Y(_09288_));
 sky130_fd_sc_hd__o32a_1 _19520_ (.A1(_04408_),
    .A2(_04441_),
    .A3(_08658_),
    .B1(_08660_),
    .B2(_03396_),
    .X(_09289_));
 sky130_fd_sc_hd__a32o_1 _19521_ (.A1(_08657_),
    .A2(_04452_),
    .A3(_04419_),
    .B1(net23),
    .B2(_08659_),
    .X(_09290_));
 sky130_fd_sc_hd__a31o_1 _19522_ (.A1(net163),
    .A2(net33),
    .A3(net319),
    .B1(_09290_),
    .X(_09291_));
 sky130_fd_sc_hd__and4_2 _19523_ (.A(net163),
    .B(net33),
    .C(net319),
    .D(_09290_),
    .X(_09293_));
 sky130_fd_sc_hd__o2111ai_4 _19524_ (.A1(_07076_),
    .A2(_08206_),
    .B1(_09290_),
    .C1(net319),
    .D1(net33),
    .Y(_09294_));
 sky130_fd_sc_hd__and3_2 _19525_ (.A(_03286_),
    .B(net319),
    .C(net44),
    .X(_09295_));
 sky130_fd_sc_hd__or3b_1 _19526_ (.A(net33),
    .B(net25),
    .C_N(net44),
    .X(_09296_));
 sky130_fd_sc_hd__o21a_4 _19527_ (.A1(net169),
    .A2(net268),
    .B1(_09295_),
    .X(_09297_));
 sky130_fd_sc_hd__o21ai_4 _19528_ (.A1(net169),
    .A2(net268),
    .B1(_09295_),
    .Y(_09298_));
 sky130_fd_sc_hd__a22oi_4 _19529_ (.A1(net25),
    .A2(_04320_),
    .B1(net163),
    .B2(_09295_),
    .Y(_09299_));
 sky130_fd_sc_hd__o2bb2ai_4 _19530_ (.A1_N(_09295_),
    .A2_N(net163),
    .B1(_04331_),
    .B2(net319),
    .Y(_09300_));
 sky130_fd_sc_hd__a21oi_2 _19531_ (.A1(_09291_),
    .A2(_09294_),
    .B1(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__a21oi_4 _19532_ (.A1(_08878_),
    .A2(_09289_),
    .B1(net148),
    .Y(_09302_));
 sky130_fd_sc_hd__a21oi_2 _19533_ (.A1(_09291_),
    .A2(_09294_),
    .B1(net148),
    .Y(_09304_));
 sky130_fd_sc_hd__and3_1 _19534_ (.A(_09291_),
    .B(_09294_),
    .C(net148),
    .X(_09305_));
 sky130_fd_sc_hd__o221a_1 _19535_ (.A1(_08878_),
    .A2(_08873_),
    .B1(_09302_),
    .B2(_09301_),
    .C1(_08888_),
    .X(_09306_));
 sky130_fd_sc_hd__o221ai_4 _19536_ (.A1(_08878_),
    .A2(_08873_),
    .B1(_09302_),
    .B2(_09301_),
    .C1(_08888_),
    .Y(_09307_));
 sky130_fd_sc_hd__o22a_1 _19537_ (.A1(_08879_),
    .A2(_08887_),
    .B1(_09304_),
    .B2(_09305_),
    .X(_09308_));
 sky130_fd_sc_hd__o22ai_4 _19538_ (.A1(_08879_),
    .A2(_08887_),
    .B1(_09304_),
    .B2(_09305_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand4_4 _19539_ (.A(_09286_),
    .B(_09288_),
    .C(_09307_),
    .D(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__o22ai_4 _19540_ (.A1(_09285_),
    .A2(_09287_),
    .B1(_09306_),
    .B2(_09308_),
    .Y(_09311_));
 sky130_fd_sc_hd__o21a_1 _19541_ (.A1(_08867_),
    .A2(_08870_),
    .B1(_08889_),
    .X(_09312_));
 sky130_fd_sc_hd__o21ai_2 _19542_ (.A1(_08890_),
    .A2(_08871_),
    .B1(_08889_),
    .Y(_09313_));
 sky130_fd_sc_hd__nand3_4 _19543_ (.A(_09313_),
    .B(_09311_),
    .C(_09310_),
    .Y(_09315_));
 sky130_fd_sc_hd__a21oi_4 _19544_ (.A1(_09310_),
    .A2(_09311_),
    .B1(_09313_),
    .Y(_09316_));
 sky130_fd_sc_hd__o2bb2ai_4 _19545_ (.A1_N(_09310_),
    .A2_N(_09311_),
    .B1(_09312_),
    .B2(_08890_),
    .Y(_09317_));
 sky130_fd_sc_hd__and2_2 _19546_ (.A(_08909_),
    .B(_08915_),
    .X(_09318_));
 sky130_fd_sc_hd__nand2_1 _19547_ (.A(_08909_),
    .B(_08915_),
    .Y(_09319_));
 sky130_fd_sc_hd__o311a_1 _19548_ (.A1(net246),
    .A2(_05928_),
    .A3(_06759_),
    .B1(net292),
    .C1(net195),
    .X(_09320_));
 sky130_fd_sc_hd__and3_1 _19549_ (.A(_03927_),
    .B(net19),
    .C(net61),
    .X(_09321_));
 sky130_fd_sc_hd__a31o_1 _19550_ (.A1(net195),
    .A2(net171),
    .A3(net292),
    .B1(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__o211ai_4 _19551_ (.A1(net175),
    .A2(_07501_),
    .B1(_05227_),
    .C1(_07499_),
    .Y(_09323_));
 sky130_fd_sc_hd__or3b_1 _19552_ (.A(net60),
    .B(_04223_),
    .C_N(net59),
    .X(_09324_));
 sky130_fd_sc_hd__a221oi_4 _19553_ (.A1(net205),
    .A2(_07073_),
    .B1(net171),
    .B2(net20),
    .C1(_05699_),
    .Y(_09326_));
 sky130_fd_sc_hd__o221ai_4 _19554_ (.A1(net175),
    .A2(_07074_),
    .B1(_04212_),
    .B2(net189),
    .C1(_05688_),
    .Y(_09327_));
 sky130_fd_sc_hd__nor2_1 _19555_ (.A(_04212_),
    .B(_05720_),
    .Y(_09328_));
 sky130_fd_sc_hd__or3b_1 _19556_ (.A(net61),
    .B(_04212_),
    .C_N(net60),
    .X(_09329_));
 sky130_fd_sc_hd__o2bb2a_2 _19557_ (.A1_N(_09323_),
    .A2_N(_09324_),
    .B1(_09326_),
    .B2(_09328_),
    .X(_09330_));
 sky130_fd_sc_hd__o2bb2ai_4 _19558_ (.A1_N(_09323_),
    .A2_N(_09324_),
    .B1(_09326_),
    .B2(_09328_),
    .Y(_09331_));
 sky130_fd_sc_hd__o2111ai_4 _19559_ (.A1(_04223_),
    .A2(_05260_),
    .B1(_09323_),
    .C1(_09327_),
    .D1(_09329_),
    .Y(_09332_));
 sky130_fd_sc_hd__a21oi_2 _19560_ (.A1(_09331_),
    .A2(_09332_),
    .B1(_09322_),
    .Y(_09333_));
 sky130_fd_sc_hd__a21o_1 _19561_ (.A1(_09331_),
    .A2(_09332_),
    .B1(_09322_),
    .X(_09334_));
 sky130_fd_sc_hd__o211a_4 _19562_ (.A1(_09320_),
    .A2(_09321_),
    .B1(_09331_),
    .C1(_09332_),
    .X(_09335_));
 sky130_fd_sc_hd__o211ai_4 _19563_ (.A1(_09320_),
    .A2(_09321_),
    .B1(_09331_),
    .C1(_09332_),
    .Y(_09337_));
 sky130_fd_sc_hd__a21oi_2 _19564_ (.A1(_08862_),
    .A2(_08866_),
    .B1(_08859_),
    .Y(_09338_));
 sky130_fd_sc_hd__a21o_1 _19565_ (.A1(_08862_),
    .A2(_08866_),
    .B1(_08859_),
    .X(_09339_));
 sky130_fd_sc_hd__a21oi_2 _19566_ (.A1(_09334_),
    .A2(_09337_),
    .B1(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__o21ai_4 _19567_ (.A1(_09333_),
    .A2(_09335_),
    .B1(_09338_),
    .Y(_09341_));
 sky130_fd_sc_hd__nand3_4 _19568_ (.A(_09334_),
    .B(_09337_),
    .C(_09339_),
    .Y(_09342_));
 sky130_fd_sc_hd__a21oi_2 _19569_ (.A1(_09341_),
    .A2(_09342_),
    .B1(_09319_),
    .Y(_09343_));
 sky130_fd_sc_hd__a21o_1 _19570_ (.A1(_09341_),
    .A2(_09342_),
    .B1(_09319_),
    .X(_09344_));
 sky130_fd_sc_hd__and3_1 _19571_ (.A(_09319_),
    .B(_09341_),
    .C(_09342_),
    .X(_09345_));
 sky130_fd_sc_hd__nand3_1 _19572_ (.A(_09319_),
    .B(_09341_),
    .C(_09342_),
    .Y(_09346_));
 sky130_fd_sc_hd__a21oi_2 _19573_ (.A1(_09341_),
    .A2(_09342_),
    .B1(_09318_),
    .Y(_09348_));
 sky130_fd_sc_hd__a22o_1 _19574_ (.A1(_08909_),
    .A2(_08915_),
    .B1(_09341_),
    .B2(_09342_),
    .X(_09349_));
 sky130_fd_sc_hd__and3_1 _19575_ (.A(_09341_),
    .B(_09342_),
    .C(_09318_),
    .X(_09350_));
 sky130_fd_sc_hd__nand4_2 _19576_ (.A(_08909_),
    .B(_08915_),
    .C(_09341_),
    .D(_09342_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand2_1 _19577_ (.A(_09344_),
    .B(_09346_),
    .Y(_09352_));
 sky130_fd_sc_hd__o211ai_2 _19578_ (.A1(_09343_),
    .A2(_09345_),
    .B1(_09315_),
    .C1(_09317_),
    .Y(_09353_));
 sky130_fd_sc_hd__o2bb2ai_1 _19579_ (.A1_N(_09315_),
    .A2_N(_09317_),
    .B1(_09348_),
    .B2(_09350_),
    .Y(_09354_));
 sky130_fd_sc_hd__o2bb2a_1 _19580_ (.A1_N(_09315_),
    .A2_N(_09317_),
    .B1(_09343_),
    .B2(_09345_),
    .X(_09355_));
 sky130_fd_sc_hd__o2bb2ai_4 _19581_ (.A1_N(_09315_),
    .A2_N(_09317_),
    .B1(_09343_),
    .B2(_09345_),
    .Y(_09356_));
 sky130_fd_sc_hd__o211ai_4 _19582_ (.A1(_09348_),
    .A2(_09350_),
    .B1(_09315_),
    .C1(_09317_),
    .Y(_09357_));
 sky130_fd_sc_hd__nand3_2 _19583_ (.A(_08898_),
    .B(_08932_),
    .C(_09357_),
    .Y(_09359_));
 sky130_fd_sc_hd__nand3_4 _19584_ (.A(_09267_),
    .B(_09356_),
    .C(_09357_),
    .Y(_09360_));
 sky130_fd_sc_hd__a22oi_4 _19585_ (.A1(_08898_),
    .A2(_08932_),
    .B1(_09356_),
    .B2(_09357_),
    .Y(_09361_));
 sky130_fd_sc_hd__o2111ai_4 _19586_ (.A1(_08929_),
    .A2(_08896_),
    .B1(_08900_),
    .C1(_09353_),
    .D1(_09354_),
    .Y(_09362_));
 sky130_fd_sc_hd__nor2_2 _19587_ (.A(_04168_),
    .B(_08283_),
    .Y(_09363_));
 sky130_fd_sc_hd__a31oi_2 _19588_ (.A1(net201),
    .A2(_06221_),
    .A3(net291),
    .B1(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__nand3_2 _19589_ (.A(net199),
    .B(net172),
    .C(_07658_),
    .Y(_09365_));
 sky130_fd_sc_hd__or3_1 _19590_ (.A(net63),
    .B(_04179_),
    .C(_03927_),
    .X(_09366_));
 sky130_fd_sc_hd__a21oi_1 _19591_ (.A1(_09365_),
    .A2(_09366_),
    .B1(_09364_),
    .Y(_09367_));
 sky130_fd_sc_hd__a21o_2 _19592_ (.A1(_09365_),
    .A2(_09366_),
    .B1(_09364_),
    .X(_09368_));
 sky130_fd_sc_hd__o221ai_4 _19593_ (.A1(_04179_),
    .A2(_07691_),
    .B1(_08261_),
    .B2(_06222_),
    .C1(_09365_),
    .Y(_09370_));
 sky130_fd_sc_hd__o211a_1 _19594_ (.A1(_04179_),
    .A2(_07691_),
    .B1(_09365_),
    .C1(_09364_),
    .X(_09371_));
 sky130_fd_sc_hd__o211ai_1 _19595_ (.A1(_04179_),
    .A2(_07691_),
    .B1(_09365_),
    .C1(_09364_),
    .Y(_09372_));
 sky130_fd_sc_hd__a32o_1 _19596_ (.A1(_05933_),
    .A2(net289),
    .A3(net175),
    .B1(_10335_),
    .B2(net16),
    .X(_09373_));
 sky130_fd_sc_hd__a21oi_1 _19597_ (.A1(_09368_),
    .A2(_09372_),
    .B1(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__o21bai_2 _19598_ (.A1(_09367_),
    .A2(_09371_),
    .B1_N(_09373_),
    .Y(_09375_));
 sky130_fd_sc_hd__o211a_1 _19599_ (.A1(_09363_),
    .A2(_09370_),
    .B1(_09373_),
    .C1(_09368_),
    .X(_09376_));
 sky130_fd_sc_hd__o211ai_4 _19600_ (.A1(_09363_),
    .A2(_09370_),
    .B1(_09373_),
    .C1(_09368_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand4_4 _19601_ (.A(_08968_),
    .B(_08971_),
    .C(_09375_),
    .D(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__o22ai_4 _19602_ (.A1(_08967_),
    .A2(_08970_),
    .B1(_09374_),
    .B2(_09376_),
    .Y(_09379_));
 sky130_fd_sc_hd__nor2_1 _19603_ (.A(_04113_),
    .B(_01326_),
    .Y(_09381_));
 sky130_fd_sc_hd__o311a_1 _19604_ (.A1(net11),
    .A2(_04557_),
    .A3(net208),
    .B1(_01293_),
    .C1(net211),
    .X(_09382_));
 sky130_fd_sc_hd__a31o_1 _19605_ (.A1(net211),
    .A2(net183),
    .A3(_01293_),
    .B1(_09381_),
    .X(_09383_));
 sky130_fd_sc_hd__nand4_1 _19606_ (.A(_03993_),
    .B(net181),
    .C(net179),
    .D(net36),
    .Y(_09384_));
 sky130_fd_sc_hd__nor2_1 _19607_ (.A(_04135_),
    .B(_12363_),
    .Y(_09385_));
 sky130_fd_sc_hd__or3_1 _19608_ (.A(net36),
    .B(_04135_),
    .C(_03993_),
    .X(_09386_));
 sky130_fd_sc_hd__a31oi_4 _19609_ (.A1(net181),
    .A2(net179),
    .A3(_12330_),
    .B1(_09385_),
    .Y(_09387_));
 sky130_fd_sc_hd__or3_1 _19610_ (.A(net35),
    .B(_04146_),
    .C(_03971_),
    .X(_09388_));
 sky130_fd_sc_hd__o2111ai_4 _19611_ (.A1(_04789_),
    .A2(_05551_),
    .B1(net35),
    .C1(net178),
    .D1(_03971_),
    .Y(_09389_));
 sky130_fd_sc_hd__a32oi_4 _19612_ (.A1(net178),
    .A2(net177),
    .A3(net252),
    .B1(_11793_),
    .B2(net15),
    .Y(_09390_));
 sky130_fd_sc_hd__o2111a_1 _19613_ (.A1(_04146_),
    .A2(_11804_),
    .B1(_09384_),
    .C1(_09386_),
    .D1(_09389_),
    .X(_09392_));
 sky130_fd_sc_hd__nand2_1 _19614_ (.A(_09387_),
    .B(_09390_),
    .Y(_09393_));
 sky130_fd_sc_hd__a21oi_4 _19615_ (.A1(_09388_),
    .A2(_09389_),
    .B1(_09387_),
    .Y(_09394_));
 sky130_fd_sc_hd__a22o_1 _19616_ (.A1(_09384_),
    .A2(_09386_),
    .B1(_09388_),
    .B2(_09389_),
    .X(_09395_));
 sky130_fd_sc_hd__o21ai_1 _19617_ (.A1(_09392_),
    .A2(_09394_),
    .B1(_09383_),
    .Y(_09396_));
 sky130_fd_sc_hd__o21bai_2 _19618_ (.A1(_09387_),
    .A2(_09390_),
    .B1_N(_09383_),
    .Y(_09397_));
 sky130_fd_sc_hd__a2bb2oi_1 _19619_ (.A1_N(_09381_),
    .A2_N(_09382_),
    .B1(_09387_),
    .B2(_09390_),
    .Y(_09398_));
 sky130_fd_sc_hd__and3_1 _19620_ (.A(_09383_),
    .B(_09393_),
    .C(_09395_),
    .X(_09399_));
 sky130_fd_sc_hd__a21oi_1 _19621_ (.A1(_09393_),
    .A2(_09395_),
    .B1(_09383_),
    .Y(_09400_));
 sky130_fd_sc_hd__o41ai_4 _19622_ (.A1(_09381_),
    .A2(_09382_),
    .A3(_09392_),
    .A4(_09394_),
    .B1(_09396_),
    .Y(_09401_));
 sky130_fd_sc_hd__nand3_4 _19623_ (.A(_09378_),
    .B(_09379_),
    .C(_09401_),
    .Y(_09403_));
 sky130_fd_sc_hd__o2bb2ai_4 _19624_ (.A1_N(_09378_),
    .A2_N(_09379_),
    .B1(_09399_),
    .B2(_09400_),
    .Y(_09404_));
 sky130_fd_sc_hd__a41o_1 _19625_ (.A1(_08968_),
    .A2(_08971_),
    .A3(_09375_),
    .A4(_09377_),
    .B1(_09401_),
    .X(_09405_));
 sky130_fd_sc_hd__a21boi_1 _19626_ (.A1(_09379_),
    .A2(_09401_),
    .B1_N(_09378_),
    .Y(_09406_));
 sky130_fd_sc_hd__nand2_1 _19627_ (.A(_09403_),
    .B(_09404_),
    .Y(_09407_));
 sky130_fd_sc_hd__a31oi_2 _19628_ (.A1(_08913_),
    .A2(_08915_),
    .A3(_08918_),
    .B1(_08902_),
    .Y(_09408_));
 sky130_fd_sc_hd__o22ai_4 _19629_ (.A1(_08922_),
    .A2(_08914_),
    .B1(_08901_),
    .B2(_08920_),
    .Y(_09409_));
 sky130_fd_sc_hd__a31o_1 _19630_ (.A1(_08614_),
    .A2(_08618_),
    .A3(_08924_),
    .B1(_08920_),
    .X(_09410_));
 sky130_fd_sc_hd__a21oi_1 _19631_ (.A1(_09403_),
    .A2(_09404_),
    .B1(_09409_),
    .Y(_09411_));
 sky130_fd_sc_hd__o2bb2ai_4 _19632_ (.A1_N(_09403_),
    .A2_N(_09404_),
    .B1(_09408_),
    .B2(_08920_),
    .Y(_09412_));
 sky130_fd_sc_hd__and3_2 _19633_ (.A(_09409_),
    .B(_09404_),
    .C(_09403_),
    .X(_09414_));
 sky130_fd_sc_hd__nand3_4 _19634_ (.A(_09409_),
    .B(_09404_),
    .C(_09403_),
    .Y(_09415_));
 sky130_fd_sc_hd__and3_1 _19635_ (.A(_08955_),
    .B(_08957_),
    .C(_08977_),
    .X(_09416_));
 sky130_fd_sc_hd__o31a_1 _19636_ (.A1(_08954_),
    .A2(_08956_),
    .A3(_08976_),
    .B1(_08979_),
    .X(_09417_));
 sky130_fd_sc_hd__a31o_1 _19637_ (.A1(_08955_),
    .A2(_08957_),
    .A3(_08977_),
    .B1(_08978_),
    .X(_09418_));
 sky130_fd_sc_hd__o22a_1 _19638_ (.A1(_09411_),
    .A2(_09414_),
    .B1(_09416_),
    .B2(_08978_),
    .X(_09419_));
 sky130_fd_sc_hd__o2bb2ai_4 _19639_ (.A1_N(_09412_),
    .A2_N(_09415_),
    .B1(_09416_),
    .B2(_08978_),
    .Y(_09420_));
 sky130_fd_sc_hd__a22oi_4 _19640_ (.A1(_08977_),
    .A2(_08980_),
    .B1(_09407_),
    .B2(_09410_),
    .Y(_09421_));
 sky130_fd_sc_hd__nand3_4 _19641_ (.A(_09412_),
    .B(_09415_),
    .C(_09417_),
    .Y(_09422_));
 sky130_fd_sc_hd__inv_2 _19642_ (.A(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__o2bb2a_1 _19643_ (.A1_N(_08977_),
    .A2_N(_08980_),
    .B1(_09411_),
    .B2(_09414_),
    .X(_09425_));
 sky130_fd_sc_hd__and3_1 _19644_ (.A(_09412_),
    .B(_09415_),
    .C(_09418_),
    .X(_09426_));
 sky130_fd_sc_hd__nand2_2 _19645_ (.A(_09420_),
    .B(_09422_),
    .Y(_09427_));
 sky130_fd_sc_hd__o2bb2ai_4 _19646_ (.A1_N(_09360_),
    .A2_N(_09362_),
    .B1(_09425_),
    .B2(_09426_),
    .Y(_09428_));
 sky130_fd_sc_hd__o211ai_4 _19647_ (.A1(_09355_),
    .A2(_09359_),
    .B1(_09362_),
    .C1(_09427_),
    .Y(_09429_));
 sky130_fd_sc_hd__o2bb2ai_2 _19648_ (.A1_N(_09360_),
    .A2_N(_09362_),
    .B1(_09419_),
    .B2(_09423_),
    .Y(_09430_));
 sky130_fd_sc_hd__nand4_4 _19649_ (.A(_09360_),
    .B(_09362_),
    .C(_09420_),
    .D(_09422_),
    .Y(_09431_));
 sky130_fd_sc_hd__a21oi_4 _19650_ (.A1(_09430_),
    .A2(_09431_),
    .B1(_09265_),
    .Y(_09432_));
 sky130_fd_sc_hd__nand3_2 _19651_ (.A(_09266_),
    .B(_09428_),
    .C(_09429_),
    .Y(_09433_));
 sky130_fd_sc_hd__a21oi_2 _19652_ (.A1(_09428_),
    .A2(_09429_),
    .B1(_09266_),
    .Y(_09434_));
 sky130_fd_sc_hd__nand3_4 _19653_ (.A(_09265_),
    .B(_09430_),
    .C(_09431_),
    .Y(_09436_));
 sky130_fd_sc_hd__a21o_1 _19654_ (.A1(_09433_),
    .A2(_09436_),
    .B1(_09264_),
    .X(_09437_));
 sky130_fd_sc_hd__o21ai_2 _19655_ (.A1(_09260_),
    .A2(_09262_),
    .B1(_09436_),
    .Y(_09438_));
 sky130_fd_sc_hd__a311oi_2 _19656_ (.A1(_09266_),
    .A2(_09428_),
    .A3(_09429_),
    .B1(_09262_),
    .C1(_09260_),
    .Y(_09439_));
 sky130_fd_sc_hd__nand4_4 _19657_ (.A(_09261_),
    .B(_09263_),
    .C(_09433_),
    .D(_09436_),
    .Y(_09440_));
 sky130_fd_sc_hd__inv_2 _19658_ (.A(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__o22ai_4 _19659_ (.A1(_09260_),
    .A2(_09262_),
    .B1(_09432_),
    .B2(_09434_),
    .Y(_09442_));
 sky130_fd_sc_hd__o21ai_1 _19660_ (.A1(_09015_),
    .A2(_09123_),
    .B1(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__and3_1 _19661_ (.A(_09442_),
    .B(_09175_),
    .C(_09440_),
    .X(_09444_));
 sky130_fd_sc_hd__o211ai_4 _19662_ (.A1(_09015_),
    .A2(_09123_),
    .B1(_09440_),
    .C1(_09442_),
    .Y(_09445_));
 sky130_fd_sc_hd__o211a_1 _19663_ (.A1(_09438_),
    .A2(_09432_),
    .B1(_09176_),
    .C1(_09437_),
    .X(_09447_));
 sky130_fd_sc_hd__o211ai_4 _19664_ (.A1(_09438_),
    .A2(_09432_),
    .B1(_09176_),
    .C1(_09437_),
    .Y(_09448_));
 sky130_fd_sc_hd__o21ai_2 _19665_ (.A1(_08775_),
    .A2(_08779_),
    .B1(_08786_),
    .Y(_09449_));
 sky130_fd_sc_hd__o21ai_1 _19666_ (.A1(_08762_),
    .A2(_08770_),
    .B1(_08769_),
    .Y(_09450_));
 sky130_fd_sc_hd__a21oi_2 _19667_ (.A1(_09079_),
    .A2(_09081_),
    .B1(_09076_),
    .Y(_09451_));
 sky130_fd_sc_hd__o21ai_1 _19668_ (.A1(_09079_),
    .A2(_09081_),
    .B1(_09076_),
    .Y(_09452_));
 sky130_fd_sc_hd__o21ai_1 _19669_ (.A1(_09078_),
    .A2(_09080_),
    .B1(_09452_),
    .Y(_09453_));
 sky130_fd_sc_hd__and3_1 _19670_ (.A(_04190_),
    .B(net49),
    .C(net31),
    .X(_09454_));
 sky130_fd_sc_hd__and3_2 _19671_ (.A(_07242_),
    .B(net257),
    .C(net273),
    .X(_09455_));
 sky130_fd_sc_hd__a21oi_2 _19672_ (.A1(net31),
    .A2(_06326_),
    .B1(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__a31o_1 _19673_ (.A1(_07242_),
    .A2(net257),
    .A3(net273),
    .B1(_09454_),
    .X(_09458_));
 sky130_fd_sc_hd__o211ai_4 _19674_ (.A1(net259),
    .A2(_09665_),
    .B1(net275),
    .C1(_09698_),
    .Y(_09459_));
 sky130_fd_sc_hd__or3b_1 _19675_ (.A(_03960_),
    .B(net48),
    .C_N(net47),
    .X(_09460_));
 sky130_fd_sc_hd__o21ai_1 _19676_ (.A1(_03960_),
    .A2(_05766_),
    .B1(_09459_),
    .Y(_09461_));
 sky130_fd_sc_hd__o211ai_1 _19677_ (.A1(net259),
    .A2(_08656_),
    .B1(net274),
    .C1(_08700_),
    .Y(_09462_));
 sky130_fd_sc_hd__nor2_1 _19678_ (.A(_03949_),
    .B(_06030_),
    .Y(_09463_));
 sky130_fd_sc_hd__a31oi_4 _19679_ (.A1(net256),
    .A2(_08700_),
    .A3(net274),
    .B1(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__o21ai_1 _19680_ (.A1(_03949_),
    .A2(_06030_),
    .B1(_09462_),
    .Y(_09465_));
 sky130_fd_sc_hd__a21oi_2 _19681_ (.A1(_09459_),
    .A2(_09460_),
    .B1(_09464_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand2_2 _19682_ (.A(_09461_),
    .B(_09465_),
    .Y(_09467_));
 sky130_fd_sc_hd__o221a_2 _19683_ (.A1(_09720_),
    .A2(_05763_),
    .B1(_05766_),
    .B2(_03960_),
    .C1(_09464_),
    .X(_09469_));
 sky130_fd_sc_hd__o211ai_4 _19684_ (.A1(_03960_),
    .A2(_05766_),
    .B1(_09459_),
    .C1(_09464_),
    .Y(_09470_));
 sky130_fd_sc_hd__o211ai_2 _19685_ (.A1(_09454_),
    .A2(_09455_),
    .B1(_09467_),
    .C1(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__a21o_1 _19686_ (.A1(_09467_),
    .A2(_09470_),
    .B1(_09458_),
    .X(_09472_));
 sky130_fd_sc_hd__o22ai_4 _19687_ (.A1(_09454_),
    .A2(_09455_),
    .B1(_09466_),
    .B2(_09469_),
    .Y(_09473_));
 sky130_fd_sc_hd__nand3_2 _19688_ (.A(_09467_),
    .B(_09470_),
    .C(_09456_),
    .Y(_09474_));
 sky130_fd_sc_hd__a22oi_2 _19689_ (.A1(_09082_),
    .A2(_09452_),
    .B1(_09473_),
    .B2(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__nand3_2 _19690_ (.A(_09472_),
    .B(_09453_),
    .C(_09471_),
    .Y(_09476_));
 sky130_fd_sc_hd__a2bb2oi_2 _19691_ (.A1_N(_09083_),
    .A2_N(_09451_),
    .B1(_09471_),
    .B2(_09472_),
    .Y(_09477_));
 sky130_fd_sc_hd__o211ai_4 _19692_ (.A1(_09083_),
    .A2(_09451_),
    .B1(_09473_),
    .C1(_09474_),
    .Y(_09478_));
 sky130_fd_sc_hd__a21oi_2 _19693_ (.A1(_09476_),
    .A2(_09478_),
    .B1(_09450_),
    .Y(_09480_));
 sky130_fd_sc_hd__o211ai_1 _19694_ (.A1(_08768_),
    .A2(_08772_),
    .B1(_09476_),
    .C1(_09478_),
    .Y(_09481_));
 sky130_fd_sc_hd__o2111ai_4 _19695_ (.A1(_08762_),
    .A2(_08770_),
    .B1(_09476_),
    .C1(_09478_),
    .D1(_08769_),
    .Y(_09482_));
 sky130_fd_sc_hd__o22ai_2 _19696_ (.A1(_08768_),
    .A2(_08772_),
    .B1(_09475_),
    .B2(_09477_),
    .Y(_09483_));
 sky130_fd_sc_hd__o21ai_1 _19697_ (.A1(_09086_),
    .A2(_09088_),
    .B1(_09074_),
    .Y(_09484_));
 sky130_fd_sc_hd__o2111a_1 _19698_ (.A1(_09090_),
    .A2(_09071_),
    .B1(_09074_),
    .C1(_09482_),
    .D1(_09483_),
    .X(_09485_));
 sky130_fd_sc_hd__o2111ai_4 _19699_ (.A1(_09090_),
    .A2(_09071_),
    .B1(_09074_),
    .C1(_09482_),
    .D1(_09483_),
    .Y(_09486_));
 sky130_fd_sc_hd__nand3_2 _19700_ (.A(_09072_),
    .B(_09481_),
    .C(_09484_),
    .Y(_09487_));
 sky130_fd_sc_hd__o21ai_1 _19701_ (.A1(_09480_),
    .A2(_09487_),
    .B1(_09486_),
    .Y(_09488_));
 sky130_fd_sc_hd__o211ai_4 _19702_ (.A1(_08775_),
    .A2(_08779_),
    .B1(_08786_),
    .C1(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__o211ai_4 _19703_ (.A1(_09480_),
    .A2(_09487_),
    .B1(_09486_),
    .C1(_09449_),
    .Y(_09491_));
 sky130_fd_sc_hd__a31oi_1 _19704_ (.A1(_08784_),
    .A2(_08789_),
    .A3(_08786_),
    .B1(_08794_),
    .Y(_09492_));
 sky130_fd_sc_hd__a21oi_1 _19705_ (.A1(_08788_),
    .A2(_08790_),
    .B1(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__a21oi_2 _19706_ (.A1(_09489_),
    .A2(_09491_),
    .B1(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__a21o_1 _19707_ (.A1(_09489_),
    .A2(_09491_),
    .B1(_09493_),
    .X(_09495_));
 sky130_fd_sc_hd__o211a_1 _19708_ (.A1(_08792_),
    .A2(_08797_),
    .B1(_09489_),
    .C1(_09491_),
    .X(_09496_));
 sky130_fd_sc_hd__o211ai_4 _19709_ (.A1(_08792_),
    .A2(_08797_),
    .B1(_09489_),
    .C1(_09491_),
    .Y(_09497_));
 sky130_fd_sc_hd__a32oi_4 _19710_ (.A1(_08005_),
    .A2(_04747_),
    .A3(net313),
    .B1(net26),
    .B2(_08006_),
    .Y(_09498_));
 sky130_fd_sc_hd__a32o_1 _19711_ (.A1(net313),
    .A2(_04747_),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net26),
    .X(_09499_));
 sky130_fd_sc_hd__a32o_1 _19712_ (.A1(net266),
    .A2(net301),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net27),
    .X(_09500_));
 sky130_fd_sc_hd__o21ai_1 _19713_ (.A1(_08810_),
    .A2(_08818_),
    .B1(_08817_),
    .Y(_09502_));
 sky130_fd_sc_hd__a21oi_1 _19714_ (.A1(_08811_),
    .A2(_08819_),
    .B1(_08816_),
    .Y(_09503_));
 sky130_fd_sc_hd__and3_1 _19715_ (.A(_04234_),
    .B(net52),
    .C(net28),
    .X(_09504_));
 sky130_fd_sc_hd__o311a_1 _19716_ (.A1(net26),
    .A2(_04452_),
    .A3(_05436_),
    .B1(_07305_),
    .C1(_05414_),
    .X(_09505_));
 sky130_fd_sc_hd__a21oi_1 _19717_ (.A1(net28),
    .A2(_07308_),
    .B1(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__or3b_2 _19718_ (.A(_03835_),
    .B(net52),
    .C_N(net51),
    .X(_09507_));
 sky130_fd_sc_hd__nand3_2 _19719_ (.A(_05841_),
    .B(net265),
    .C(_07223_),
    .Y(_09508_));
 sky130_fd_sc_hd__or3_2 _19720_ (.A(net51),
    .B(_04190_),
    .C(_03916_),
    .X(_09509_));
 sky130_fd_sc_hd__o211ai_4 _19721_ (.A1(_04747_),
    .A2(net264),
    .B1(_06863_),
    .C1(_06486_),
    .Y(_09510_));
 sky130_fd_sc_hd__a22oi_4 _19722_ (.A1(_09507_),
    .A2(_09508_),
    .B1(_09509_),
    .B2(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__a22o_1 _19723_ (.A1(_09507_),
    .A2(_09508_),
    .B1(_09509_),
    .B2(_09510_),
    .X(_09513_));
 sky130_fd_sc_hd__o2111a_1 _19724_ (.A1(_03835_),
    .A2(_07226_),
    .B1(_09508_),
    .C1(_09509_),
    .D1(_09510_),
    .X(_09514_));
 sky130_fd_sc_hd__o2111ai_2 _19725_ (.A1(_03835_),
    .A2(_07226_),
    .B1(_09508_),
    .C1(_09509_),
    .D1(_09510_),
    .Y(_09515_));
 sky130_fd_sc_hd__nor3_1 _19726_ (.A(_09504_),
    .B(_09505_),
    .C(_09511_),
    .Y(_09516_));
 sky130_fd_sc_hd__o21a_1 _19727_ (.A1(_09504_),
    .A2(_09505_),
    .B1(_09515_),
    .X(_09517_));
 sky130_fd_sc_hd__nand3_1 _19728_ (.A(_09513_),
    .B(_09515_),
    .C(_09506_),
    .Y(_09518_));
 sky130_fd_sc_hd__o22ai_1 _19729_ (.A1(_09504_),
    .A2(_09505_),
    .B1(_09511_),
    .B2(_09514_),
    .Y(_09519_));
 sky130_fd_sc_hd__o21ai_1 _19730_ (.A1(_09511_),
    .A2(_09514_),
    .B1(_09506_),
    .Y(_09520_));
 sky130_fd_sc_hd__o211ai_1 _19731_ (.A1(_09504_),
    .A2(_09505_),
    .B1(_09513_),
    .C1(_09515_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand3_1 _19732_ (.A(_09520_),
    .B(_09521_),
    .C(_09502_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand3_1 _19733_ (.A(_09503_),
    .B(_09518_),
    .C(_09519_),
    .Y(_09524_));
 sky130_fd_sc_hd__a21o_1 _19734_ (.A1(_09522_),
    .A2(_09524_),
    .B1(_09500_),
    .X(_09525_));
 sky130_fd_sc_hd__nand2_1 _19735_ (.A(_09500_),
    .B(_09524_),
    .Y(_09526_));
 sky130_fd_sc_hd__nand3_1 _19736_ (.A(_09500_),
    .B(_09522_),
    .C(_09524_),
    .Y(_09527_));
 sky130_fd_sc_hd__nand2b_1 _19737_ (.A_N(_08825_),
    .B(_08823_),
    .Y(_09528_));
 sky130_fd_sc_hd__a22o_1 _19738_ (.A1(_09525_),
    .A2(_09527_),
    .B1(_09528_),
    .B2(_08824_),
    .X(_09529_));
 sky130_fd_sc_hd__inv_2 _19739_ (.A(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__and4_1 _19740_ (.A(_08824_),
    .B(_09525_),
    .C(_09527_),
    .D(_09528_),
    .X(_09531_));
 sky130_fd_sc_hd__nand4_2 _19741_ (.A(_08824_),
    .B(_09525_),
    .C(_09527_),
    .D(_09528_),
    .Y(_09532_));
 sky130_fd_sc_hd__nand2_1 _19742_ (.A(_09529_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__and3_1 _19743_ (.A(_09499_),
    .B(_09529_),
    .C(_09532_),
    .X(_09535_));
 sky130_fd_sc_hd__a21oi_1 _19744_ (.A1(_09529_),
    .A2(_09532_),
    .B1(_09499_),
    .Y(_09536_));
 sky130_fd_sc_hd__nor2_2 _19745_ (.A(_09535_),
    .B(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__or2_2 _19746_ (.A(_09535_),
    .B(_09536_),
    .X(_09538_));
 sky130_fd_sc_hd__o21ai_4 _19747_ (.A1(_09494_),
    .A2(_09496_),
    .B1(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__nand3_4 _19748_ (.A(_09495_),
    .B(_09497_),
    .C(_09537_),
    .Y(_09540_));
 sky130_fd_sc_hd__o2bb2ai_2 _19749_ (.A1_N(_09108_),
    .A2_N(_09103_),
    .B1(_09098_),
    .B2(_09104_),
    .Y(_09541_));
 sky130_fd_sc_hd__a21oi_4 _19750_ (.A1(_09539_),
    .A2(_09540_),
    .B1(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__a21o_1 _19751_ (.A1(_09539_),
    .A2(_09540_),
    .B1(_09541_),
    .X(_09543_));
 sky130_fd_sc_hd__a32oi_4 _19752_ (.A1(_09495_),
    .A2(_09497_),
    .A3(_09537_),
    .B1(_09115_),
    .B2(_09107_),
    .Y(_09544_));
 sky130_fd_sc_hd__o211ai_4 _19753_ (.A1(_09105_),
    .A2(_09114_),
    .B1(_09539_),
    .C1(_09540_),
    .Y(_09546_));
 sky130_fd_sc_hd__inv_2 _19754_ (.A(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__o31a_2 _19755_ (.A1(_08761_),
    .A2(_08795_),
    .A3(_08799_),
    .B1(_08835_),
    .X(_09548_));
 sky130_fd_sc_hd__a221oi_4 _19756_ (.A1(_08805_),
    .A2(_08835_),
    .B1(_09544_),
    .B2(_09539_),
    .C1(_09542_),
    .Y(_09549_));
 sky130_fd_sc_hd__a221o_2 _19757_ (.A1(_08805_),
    .A2(_08835_),
    .B1(_09544_),
    .B2(_09539_),
    .C1(_09542_),
    .X(_09550_));
 sky130_fd_sc_hd__a21boi_2 _19758_ (.A1(_09543_),
    .A2(_09546_),
    .B1_N(_09548_),
    .Y(_09551_));
 sky130_fd_sc_hd__o21ai_4 _19759_ (.A1(_09542_),
    .A2(_09547_),
    .B1(_09548_),
    .Y(_09552_));
 sky130_fd_sc_hd__nor2_1 _19760_ (.A(_09549_),
    .B(_09551_),
    .Y(_09553_));
 sky130_fd_sc_hd__o2bb2ai_4 _19761_ (.A1_N(_09445_),
    .A2_N(_09448_),
    .B1(_09549_),
    .B2(_09551_),
    .Y(_09554_));
 sky130_fd_sc_hd__nand2_1 _19762_ (.A(_09448_),
    .B(_09553_),
    .Y(_09555_));
 sky130_fd_sc_hd__and3_1 _19763_ (.A(_09445_),
    .B(_09448_),
    .C(_09553_),
    .X(_09557_));
 sky130_fd_sc_hd__nand4_4 _19764_ (.A(_09445_),
    .B(_09448_),
    .C(_09550_),
    .D(_09552_),
    .Y(_09558_));
 sky130_fd_sc_hd__a22oi_4 _19765_ (.A1(_09127_),
    .A2(_09133_),
    .B1(_09554_),
    .B2(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__a22o_1 _19766_ (.A1(_09127_),
    .A2(_09133_),
    .B1(_09554_),
    .B2(_09558_),
    .X(_09560_));
 sky130_fd_sc_hd__nand2_1 _19767_ (.A(_09554_),
    .B(_09134_),
    .Y(_09561_));
 sky130_fd_sc_hd__o211a_1 _19768_ (.A1(_09444_),
    .A2(_09555_),
    .B1(_09134_),
    .C1(_09554_),
    .X(_09562_));
 sky130_fd_sc_hd__a21o_1 _19769_ (.A1(_08838_),
    .A2(_08841_),
    .B1(_08839_),
    .X(_09563_));
 sky130_fd_sc_hd__inv_2 _19770_ (.A(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__o21bai_1 _19771_ (.A1(_09559_),
    .A2(_09562_),
    .B1_N(_09563_),
    .Y(_09565_));
 sky130_fd_sc_hd__o221ai_2 _19772_ (.A1(_08839_),
    .A2(_08845_),
    .B1(_09557_),
    .B2(_09561_),
    .C1(_09560_),
    .Y(_09566_));
 sky130_fd_sc_hd__o211ai_2 _19773_ (.A1(_09557_),
    .A2(_09561_),
    .B1(_09564_),
    .C1(_09560_),
    .Y(_09568_));
 sky130_fd_sc_hd__o22ai_2 _19774_ (.A1(_08839_),
    .A2(_08845_),
    .B1(_09559_),
    .B2(_09562_),
    .Y(_09569_));
 sky130_fd_sc_hd__nand3_1 _19775_ (.A(_09174_),
    .B(_09568_),
    .C(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__a21oi_1 _19776_ (.A1(_09568_),
    .A2(_09569_),
    .B1(_09174_),
    .Y(_09571_));
 sky130_fd_sc_hd__nand3_2 _19777_ (.A(_09173_),
    .B(_09565_),
    .C(_09566_),
    .Y(_09572_));
 sky130_fd_sc_hd__a221oi_1 _19778_ (.A1(_04463_),
    .A2(_08005_),
    .B1(_08006_),
    .B2(net23),
    .C1(_08829_),
    .Y(_09573_));
 sky130_fd_sc_hd__nor2_1 _19779_ (.A(_08806_),
    .B(_08828_),
    .Y(_09574_));
 sky130_fd_sc_hd__nor2_1 _19780_ (.A(_08829_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__o2bb2ai_2 _19781_ (.A1_N(_09570_),
    .A2_N(_09572_),
    .B1(_09573_),
    .B2(_08828_),
    .Y(_09576_));
 sky130_fd_sc_hd__a31oi_1 _19782_ (.A1(_09174_),
    .A2(_09568_),
    .A3(_09569_),
    .B1(_09575_),
    .Y(_09577_));
 sky130_fd_sc_hd__a31o_1 _19783_ (.A1(_09174_),
    .A2(_09568_),
    .A3(_09569_),
    .B1(_09575_),
    .X(_09579_));
 sky130_fd_sc_hd__o211ai_2 _19784_ (.A1(_08829_),
    .A2(_09574_),
    .B1(_09572_),
    .C1(_09570_),
    .Y(_09580_));
 sky130_fd_sc_hd__o21a_1 _19785_ (.A1(_08423_),
    .A2(_09153_),
    .B1(_09152_),
    .X(_09581_));
 sky130_fd_sc_hd__a21oi_1 _19786_ (.A1(_09152_),
    .A2(_09154_),
    .B1(_09148_),
    .Y(_09582_));
 sky130_fd_sc_hd__a21oi_1 _19787_ (.A1(_09576_),
    .A2(_09580_),
    .B1(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__o2bb2ai_1 _19788_ (.A1_N(_09576_),
    .A2_N(_09580_),
    .B1(_09581_),
    .B2(_09148_),
    .Y(_09584_));
 sky130_fd_sc_hd__o211ai_2 _19789_ (.A1(_09151_),
    .A2(_09155_),
    .B1(_09576_),
    .C1(_09580_),
    .Y(_09585_));
 sky130_fd_sc_hd__nand2_1 _19790_ (.A(_09584_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__o21ai_1 _19791_ (.A1(_09162_),
    .A2(_09170_),
    .B1(_09160_),
    .Y(_09587_));
 sky130_fd_sc_hd__xnor2_1 _19792_ (.A(_09586_),
    .B(_09587_),
    .Y(net91));
 sky130_fd_sc_hd__a32oi_4 _19793_ (.A1(_09175_),
    .A2(_09440_),
    .A3(_09442_),
    .B1(_09550_),
    .B2(_09552_),
    .Y(_09589_));
 sky130_fd_sc_hd__o2bb2ai_1 _19794_ (.A1_N(_09553_),
    .A2_N(_09448_),
    .B1(_09443_),
    .B2(_09441_),
    .Y(_09590_));
 sky130_fd_sc_hd__o311a_1 _19795_ (.A1(_04747_),
    .A2(net264),
    .A3(_08656_),
    .B1(net273),
    .C1(_08700_),
    .X(_09591_));
 sky130_fd_sc_hd__and3_1 _19796_ (.A(_04190_),
    .B(net49),
    .C(net32),
    .X(_09592_));
 sky130_fd_sc_hd__a31o_1 _19797_ (.A1(net256),
    .A2(_08700_),
    .A3(net273),
    .B1(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__a31oi_2 _19798_ (.A1(net310),
    .A2(net294),
    .A3(net290),
    .B1(_06028_),
    .Y(_09594_));
 sky130_fd_sc_hd__a22oi_2 _19799_ (.A1(net2),
    .A2(_06029_),
    .B1(_09698_),
    .B2(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__a22o_1 _19800_ (.A1(net2),
    .A2(_06029_),
    .B1(_09698_),
    .B2(_09594_),
    .X(_09596_));
 sky130_fd_sc_hd__nor2_1 _19801_ (.A(_03982_),
    .B(_05766_),
    .Y(_09597_));
 sky130_fd_sc_hd__o311a_1 _19802_ (.A1(_04747_),
    .A2(net264),
    .A3(_11387_),
    .B1(net275),
    .C1(_11354_),
    .X(_09598_));
 sky130_fd_sc_hd__o221ai_4 _19803_ (.A1(_11453_),
    .A2(_05763_),
    .B1(_05766_),
    .B2(_03982_),
    .C1(_09595_),
    .Y(_09600_));
 sky130_fd_sc_hd__o21ai_4 _19804_ (.A1(_09597_),
    .A2(_09598_),
    .B1(_09596_),
    .Y(_09601_));
 sky130_fd_sc_hd__o211a_1 _19805_ (.A1(_09591_),
    .A2(_09592_),
    .B1(_09600_),
    .C1(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__o211ai_4 _19806_ (.A1(_09591_),
    .A2(_09592_),
    .B1(_09600_),
    .C1(_09601_),
    .Y(_09603_));
 sky130_fd_sc_hd__a21oi_2 _19807_ (.A1(_09600_),
    .A2(_09601_),
    .B1(_09593_),
    .Y(_09604_));
 sky130_fd_sc_hd__a21o_1 _19808_ (.A1(_09600_),
    .A2(_09601_),
    .B1(_09593_),
    .X(_09605_));
 sky130_fd_sc_hd__a21o_1 _19809_ (.A1(_09199_),
    .A2(_09206_),
    .B1(_09203_),
    .X(_09606_));
 sky130_fd_sc_hd__a21oi_2 _19810_ (.A1(_09199_),
    .A2(_09206_),
    .B1(_09203_),
    .Y(_09607_));
 sky130_fd_sc_hd__o21a_1 _19811_ (.A1(_09602_),
    .A2(_09604_),
    .B1(_09607_),
    .X(_09608_));
 sky130_fd_sc_hd__o21ai_4 _19812_ (.A1(_09602_),
    .A2(_09604_),
    .B1(_09607_),
    .Y(_09609_));
 sky130_fd_sc_hd__and3_1 _19813_ (.A(_09603_),
    .B(_09605_),
    .C(_09606_),
    .X(_09611_));
 sky130_fd_sc_hd__nand3_2 _19814_ (.A(_09603_),
    .B(_09605_),
    .C(_09606_),
    .Y(_09612_));
 sky130_fd_sc_hd__a21oi_1 _19815_ (.A1(_09461_),
    .A2(_09465_),
    .B1(_09458_),
    .Y(_09613_));
 sky130_fd_sc_hd__a21o_1 _19816_ (.A1(_09458_),
    .A2(_09470_),
    .B1(_09466_),
    .X(_09614_));
 sky130_fd_sc_hd__a31o_1 _19817_ (.A1(_09459_),
    .A2(_09460_),
    .A3(_09464_),
    .B1(_09613_),
    .X(_09615_));
 sky130_fd_sc_hd__nor2_1 _19818_ (.A(_09615_),
    .B(_09608_),
    .Y(_09616_));
 sky130_fd_sc_hd__nand2_1 _19819_ (.A(_09609_),
    .B(_09614_),
    .Y(_09617_));
 sky130_fd_sc_hd__nand3_1 _19820_ (.A(_09609_),
    .B(_09612_),
    .C(_09614_),
    .Y(_09618_));
 sky130_fd_sc_hd__o2bb2ai_1 _19821_ (.A1_N(_09609_),
    .A2_N(_09612_),
    .B1(_09613_),
    .B2(_09469_),
    .Y(_09619_));
 sky130_fd_sc_hd__a21o_1 _19822_ (.A1(_09609_),
    .A2(_09612_),
    .B1(_09615_),
    .X(_09620_));
 sky130_fd_sc_hd__o2111ai_4 _19823_ (.A1(_09456_),
    .A2(_09469_),
    .B1(_09609_),
    .C1(_09612_),
    .D1(_09467_),
    .Y(_09622_));
 sky130_fd_sc_hd__a21oi_2 _19824_ (.A1(_09197_),
    .A2(_09209_),
    .B1(_09195_),
    .Y(_09623_));
 sky130_fd_sc_hd__a21o_1 _19825_ (.A1(_09197_),
    .A2(_09209_),
    .B1(_09195_),
    .X(_09624_));
 sky130_fd_sc_hd__nand3_1 _19826_ (.A(_09620_),
    .B(_09622_),
    .C(_09623_),
    .Y(_09625_));
 sky130_fd_sc_hd__and3_1 _19827_ (.A(_09618_),
    .B(_09619_),
    .C(_09624_),
    .X(_09626_));
 sky130_fd_sc_hd__o211ai_2 _19828_ (.A1(_09611_),
    .A2(_09617_),
    .B1(_09619_),
    .C1(_09624_),
    .Y(_09627_));
 sky130_fd_sc_hd__and3_1 _19829_ (.A(_08769_),
    .B(_08773_),
    .C(_09476_),
    .X(_09628_));
 sky130_fd_sc_hd__o31a_1 _19830_ (.A1(_08768_),
    .A2(_08772_),
    .A3(_09475_),
    .B1(_09478_),
    .X(_09629_));
 sky130_fd_sc_hd__a31o_1 _19831_ (.A1(_08769_),
    .A2(_08773_),
    .A3(_09476_),
    .B1(_09477_),
    .X(_09630_));
 sky130_fd_sc_hd__o2bb2ai_2 _19832_ (.A1_N(_09625_),
    .A2_N(_09627_),
    .B1(_09628_),
    .B2(_09477_),
    .Y(_09631_));
 sky130_fd_sc_hd__a31oi_4 _19833_ (.A1(_09620_),
    .A2(_09623_),
    .A3(_09622_),
    .B1(_09630_),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2_1 _19834_ (.A(_09633_),
    .B(_09627_),
    .Y(_09634_));
 sky130_fd_sc_hd__o211a_1 _19835_ (.A1(_09480_),
    .A2(_09487_),
    .B1(_08781_),
    .C1(_08786_),
    .X(_09635_));
 sky130_fd_sc_hd__a2bb2o_1 _19836_ (.A1_N(_09480_),
    .A2_N(_09487_),
    .B1(_09486_),
    .B2(_09449_),
    .X(_09636_));
 sky130_fd_sc_hd__o2bb2a_1 _19837_ (.A1_N(_09631_),
    .A2_N(_09634_),
    .B1(_09635_),
    .B2(_09485_),
    .X(_09637_));
 sky130_fd_sc_hd__o2bb2ai_1 _19838_ (.A1_N(_09631_),
    .A2_N(_09634_),
    .B1(_09635_),
    .B2(_09485_),
    .Y(_09638_));
 sky130_fd_sc_hd__nand3_2 _19839_ (.A(_09636_),
    .B(_09634_),
    .C(_09631_),
    .Y(_09639_));
 sky130_fd_sc_hd__nand2_1 _19840_ (.A(_09638_),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__a32o_2 _19841_ (.A1(net266),
    .A2(net301),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net27),
    .X(_09641_));
 sky130_fd_sc_hd__o311a_2 _19842_ (.A1(net26),
    .A2(_04452_),
    .A3(_05436_),
    .B1(_07642_),
    .C1(_05414_),
    .X(_09642_));
 sky130_fd_sc_hd__and3b_1 _19843_ (.A_N(net54),
    .B(net53),
    .C(net28),
    .X(_09644_));
 sky130_fd_sc_hd__a21oi_1 _19844_ (.A1(net28),
    .A2(_07643_),
    .B1(_09642_),
    .Y(_09645_));
 sky130_fd_sc_hd__or3b_1 _19845_ (.A(_03916_),
    .B(net52),
    .C_N(net51),
    .X(_09646_));
 sky130_fd_sc_hd__o211ai_4 _19846_ (.A1(_04747_),
    .A2(net264),
    .B1(_07223_),
    .C1(_06486_),
    .Y(_09647_));
 sky130_fd_sc_hd__or3_2 _19847_ (.A(net51),
    .B(_04190_),
    .C(_03938_),
    .X(_09648_));
 sky130_fd_sc_hd__nand3_2 _19848_ (.A(_07242_),
    .B(net257),
    .C(_06863_),
    .Y(_09649_));
 sky130_fd_sc_hd__a22oi_2 _19849_ (.A1(_09646_),
    .A2(_09647_),
    .B1(_09648_),
    .B2(_09649_),
    .Y(_09650_));
 sky130_fd_sc_hd__a22o_1 _19850_ (.A1(_09646_),
    .A2(_09647_),
    .B1(_09648_),
    .B2(_09649_),
    .X(_09651_));
 sky130_fd_sc_hd__o2111a_1 _19851_ (.A1(_03916_),
    .A2(_07226_),
    .B1(_09647_),
    .C1(_09648_),
    .D1(_09649_),
    .X(_09652_));
 sky130_fd_sc_hd__o2111ai_4 _19852_ (.A1(_03916_),
    .A2(_07226_),
    .B1(_09647_),
    .C1(_09648_),
    .D1(_09649_),
    .Y(_09653_));
 sky130_fd_sc_hd__a32o_1 _19853_ (.A1(_05841_),
    .A2(net265),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net29),
    .X(_09655_));
 sky130_fd_sc_hd__nand3_1 _19854_ (.A(_09651_),
    .B(_09653_),
    .C(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__a21oi_1 _19855_ (.A1(_09651_),
    .A2(_09653_),
    .B1(_09655_),
    .Y(_09657_));
 sky130_fd_sc_hd__o21bai_1 _19856_ (.A1(_09650_),
    .A2(_09652_),
    .B1_N(_09655_),
    .Y(_09658_));
 sky130_fd_sc_hd__a2bb2oi_1 _19857_ (.A1_N(_09514_),
    .A2_N(_09516_),
    .B1(_09656_),
    .B2(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__a2bb2o_1 _19858_ (.A1_N(_09514_),
    .A2_N(_09516_),
    .B1(_09656_),
    .B2(_09658_),
    .X(_09660_));
 sky130_fd_sc_hd__o21ai_1 _19859_ (.A1(_09511_),
    .A2(_09517_),
    .B1(_09656_),
    .Y(_09661_));
 sky130_fd_sc_hd__o211a_1 _19860_ (.A1(_09511_),
    .A2(_09517_),
    .B1(_09656_),
    .C1(_09658_),
    .X(_09662_));
 sky130_fd_sc_hd__or2_1 _19861_ (.A(_09657_),
    .B(_09661_),
    .X(_09663_));
 sky130_fd_sc_hd__o21ai_1 _19862_ (.A1(_09659_),
    .A2(_09662_),
    .B1(_09645_),
    .Y(_09664_));
 sky130_fd_sc_hd__o221ai_2 _19863_ (.A1(_09642_),
    .A2(_09644_),
    .B1(_09657_),
    .B2(_09661_),
    .C1(_09660_),
    .Y(_09666_));
 sky130_fd_sc_hd__o211ai_1 _19864_ (.A1(_09657_),
    .A2(_09661_),
    .B1(_09645_),
    .C1(_09660_),
    .Y(_09667_));
 sky130_fd_sc_hd__o22ai_1 _19865_ (.A1(_09642_),
    .A2(_09644_),
    .B1(_09659_),
    .B2(_09662_),
    .Y(_09668_));
 sky130_fd_sc_hd__a32o_1 _19866_ (.A1(_09502_),
    .A2(_09520_),
    .A3(_09521_),
    .B1(_09524_),
    .B2(_09500_),
    .X(_09669_));
 sky130_fd_sc_hd__a22oi_2 _19867_ (.A1(_09522_),
    .A2(_09526_),
    .B1(_09667_),
    .B2(_09668_),
    .Y(_09670_));
 sky130_fd_sc_hd__a21oi_1 _19868_ (.A1(_09664_),
    .A2(_09666_),
    .B1(_09669_),
    .Y(_09671_));
 sky130_fd_sc_hd__nor2_1 _19869_ (.A(_09670_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__nor2_1 _19870_ (.A(_09641_),
    .B(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__and2_1 _19871_ (.A(_09672_),
    .B(_09641_),
    .X(_09674_));
 sky130_fd_sc_hd__xnor2_2 _19872_ (.A(_09641_),
    .B(_09672_),
    .Y(_09675_));
 sky130_fd_sc_hd__nor2_2 _19873_ (.A(_09673_),
    .B(_09674_),
    .Y(_09677_));
 sky130_fd_sc_hd__nand2_1 _19874_ (.A(_09640_),
    .B(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__a31oi_2 _19875_ (.A1(_09631_),
    .A2(_09634_),
    .A3(_09636_),
    .B1(_09677_),
    .Y(_09679_));
 sky130_fd_sc_hd__nand3_1 _19876_ (.A(_09675_),
    .B(_09639_),
    .C(_09638_),
    .Y(_09680_));
 sky130_fd_sc_hd__nand2_1 _19877_ (.A(_09640_),
    .B(_09675_),
    .Y(_09681_));
 sky130_fd_sc_hd__nand3_2 _19878_ (.A(_09638_),
    .B(_09639_),
    .C(_09677_),
    .Y(_09682_));
 sky130_fd_sc_hd__nand2_1 _19879_ (.A(_09681_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__a31o_1 _19880_ (.A1(_08994_),
    .A2(_09252_),
    .A3(_09254_),
    .B1(_09258_),
    .X(_09684_));
 sky130_fd_sc_hd__nand2_1 _19881_ (.A(_09255_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__nand4_2 _19882_ (.A(_09256_),
    .B(_09261_),
    .C(_09678_),
    .D(_09680_),
    .Y(_09686_));
 sky130_fd_sc_hd__and4_1 _19883_ (.A(_09255_),
    .B(_09681_),
    .C(_09682_),
    .D(_09684_),
    .X(_09688_));
 sky130_fd_sc_hd__nand4_4 _19884_ (.A(_09255_),
    .B(_09681_),
    .C(_09682_),
    .D(_09684_),
    .Y(_09689_));
 sky130_fd_sc_hd__o21ai_2 _19885_ (.A1(_09494_),
    .A2(_09538_),
    .B1(_09497_),
    .Y(_09690_));
 sky130_fd_sc_hd__a21oi_2 _19886_ (.A1(_09686_),
    .A2(_09689_),
    .B1(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__a21o_1 _19887_ (.A1(_09686_),
    .A2(_09689_),
    .B1(_09690_),
    .X(_09692_));
 sky130_fd_sc_hd__a22oi_1 _19888_ (.A1(_09497_),
    .A2(_09540_),
    .B1(_09685_),
    .B2(_09683_),
    .Y(_09693_));
 sky130_fd_sc_hd__nand2_1 _19889_ (.A(_09686_),
    .B(_09690_),
    .Y(_09694_));
 sky130_fd_sc_hd__and3_1 _19890_ (.A(_09686_),
    .B(_09689_),
    .C(_09690_),
    .X(_09695_));
 sky130_fd_sc_hd__a21oi_1 _19891_ (.A1(_09689_),
    .A2(_09693_),
    .B1(_09691_),
    .Y(_09696_));
 sky130_fd_sc_hd__o21ai_1 _19892_ (.A1(_09688_),
    .A2(_09694_),
    .B1(_09692_),
    .Y(_09697_));
 sky130_fd_sc_hd__a32oi_1 _19893_ (.A1(_09266_),
    .A2(_09428_),
    .A3(_09429_),
    .B1(_09436_),
    .B2(_09264_),
    .Y(_09699_));
 sky130_fd_sc_hd__a32o_1 _19894_ (.A1(_09266_),
    .A2(_09428_),
    .A3(_09429_),
    .B1(_09436_),
    .B2(_09264_),
    .X(_09700_));
 sky130_fd_sc_hd__a32oi_4 _19895_ (.A1(_09267_),
    .A2(_09356_),
    .A3(_09357_),
    .B1(_09420_),
    .B2(_09422_),
    .Y(_09701_));
 sky130_fd_sc_hd__nand2_2 _19896_ (.A(_09360_),
    .B(_09427_),
    .Y(_09702_));
 sky130_fd_sc_hd__o22ai_1 _19897_ (.A1(_09355_),
    .A2(_09359_),
    .B1(_09427_),
    .B2(_09361_),
    .Y(_09703_));
 sky130_fd_sc_hd__a31oi_4 _19898_ (.A1(_09315_),
    .A2(_09349_),
    .A3(_09351_),
    .B1(_09316_),
    .Y(_09704_));
 sky130_fd_sc_hd__o311a_1 _19899_ (.A1(net246),
    .A2(_05928_),
    .A3(_07074_),
    .B1(net292),
    .C1(_07072_),
    .X(_09705_));
 sky130_fd_sc_hd__and3_1 _19900_ (.A(_03927_),
    .B(net20),
    .C(net61),
    .X(_09706_));
 sky130_fd_sc_hd__a31o_2 _19901_ (.A1(_07072_),
    .A2(net168),
    .A3(net292),
    .B1(_09706_),
    .X(_09707_));
 sky130_fd_sc_hd__nand3_2 _19902_ (.A(_07771_),
    .B(_05227_),
    .C(_07769_),
    .Y(_09708_));
 sky130_fd_sc_hd__or3b_2 _19903_ (.A(net60),
    .B(_04245_),
    .C_N(net59),
    .X(_09710_));
 sky130_fd_sc_hd__nor2_1 _19904_ (.A(_04223_),
    .B(_05720_),
    .Y(_09711_));
 sky130_fd_sc_hd__or3b_1 _19905_ (.A(net61),
    .B(_04223_),
    .C_N(net60),
    .X(_09712_));
 sky130_fd_sc_hd__nand2_1 _19906_ (.A(net167),
    .B(_05688_),
    .Y(_09713_));
 sky130_fd_sc_hd__a21oi_1 _19907_ (.A1(net21),
    .A2(net168),
    .B1(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__nand3_1 _19908_ (.A(_07499_),
    .B(net167),
    .C(_05688_),
    .Y(_09715_));
 sky130_fd_sc_hd__o2bb2a_1 _19909_ (.A1_N(_09708_),
    .A2_N(_09710_),
    .B1(_09711_),
    .B2(_09714_),
    .X(_09716_));
 sky130_fd_sc_hd__o2bb2ai_4 _19910_ (.A1_N(_09708_),
    .A2_N(_09710_),
    .B1(_09711_),
    .B2(_09714_),
    .Y(_09717_));
 sky130_fd_sc_hd__nand4_4 _19911_ (.A(_09708_),
    .B(_09710_),
    .C(_09712_),
    .D(_09715_),
    .Y(_09718_));
 sky130_fd_sc_hd__a21oi_4 _19912_ (.A1(_09717_),
    .A2(_09718_),
    .B1(_09707_),
    .Y(_09719_));
 sky130_fd_sc_hd__a21o_1 _19913_ (.A1(_09717_),
    .A2(_09718_),
    .B1(_09707_),
    .X(_09721_));
 sky130_fd_sc_hd__o211a_2 _19914_ (.A1(_09705_),
    .A2(_09706_),
    .B1(_09717_),
    .C1(_09718_),
    .X(_09722_));
 sky130_fd_sc_hd__o211ai_4 _19915_ (.A1(_09705_),
    .A2(_09706_),
    .B1(_09717_),
    .C1(_09718_),
    .Y(_09723_));
 sky130_fd_sc_hd__o211a_1 _19916_ (.A1(_09719_),
    .A2(_09722_),
    .B1(_09279_),
    .C1(_09283_),
    .X(_09724_));
 sky130_fd_sc_hd__o211ai_4 _19917_ (.A1(_09719_),
    .A2(_09722_),
    .B1(_09279_),
    .C1(_09283_),
    .Y(_09725_));
 sky130_fd_sc_hd__a21o_1 _19918_ (.A1(_09279_),
    .A2(_09283_),
    .B1(_09722_),
    .X(_09726_));
 sky130_fd_sc_hd__nand3_2 _19919_ (.A(_09284_),
    .B(_09721_),
    .C(_09723_),
    .Y(_09727_));
 sky130_fd_sc_hd__a21o_1 _19920_ (.A1(_09322_),
    .A2(_09332_),
    .B1(_09330_),
    .X(_09728_));
 sky130_fd_sc_hd__a21oi_4 _19921_ (.A1(_09725_),
    .A2(_09727_),
    .B1(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__a21o_1 _19922_ (.A1(_09725_),
    .A2(_09727_),
    .B1(_09728_),
    .X(_09730_));
 sky130_fd_sc_hd__o211a_2 _19923_ (.A1(_09330_),
    .A2(_09335_),
    .B1(_09725_),
    .C1(_09727_),
    .X(_09732_));
 sky130_fd_sc_hd__o221ai_4 _19924_ (.A1(_09330_),
    .A2(_09335_),
    .B1(_09719_),
    .B2(_09726_),
    .C1(_09725_),
    .Y(_09733_));
 sky130_fd_sc_hd__nor2_1 _19925_ (.A(_09729_),
    .B(_09732_),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_1 _19926_ (.A(_09730_),
    .B(_09733_),
    .Y(_09735_));
 sky130_fd_sc_hd__a32o_2 _19927_ (.A1(_08657_),
    .A2(net267),
    .A3(net314),
    .B1(net26),
    .B2(_08659_),
    .X(_09736_));
 sky130_fd_sc_hd__a31oi_4 _19928_ (.A1(net162),
    .A2(net33),
    .A3(net319),
    .B1(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__and3_1 _19929_ (.A(_09736_),
    .B(net33),
    .C(net319),
    .X(_09738_));
 sky130_fd_sc_hd__nand3_1 _19930_ (.A(_09736_),
    .B(net33),
    .C(net319),
    .Y(_09739_));
 sky130_fd_sc_hd__o221ai_4 _19931_ (.A1(_09296_),
    .A2(_08207_),
    .B1(_09738_),
    .B2(_09737_),
    .C1(_08882_),
    .Y(_09740_));
 sky130_fd_sc_hd__o22a_4 _19932_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_09736_),
    .B2(_08877_),
    .X(_09741_));
 sky130_fd_sc_hd__o21ai_2 _19933_ (.A1(_09737_),
    .A2(_09738_),
    .B1(_09300_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand3b_2 _19934_ (.A_N(_09737_),
    .B(_09739_),
    .C(net148),
    .Y(_09744_));
 sky130_fd_sc_hd__a21oi_2 _19935_ (.A1(_09291_),
    .A2(_09300_),
    .B1(_09293_),
    .Y(_09745_));
 sky130_fd_sc_hd__nand3_4 _19936_ (.A(_09743_),
    .B(_09744_),
    .C(_09745_),
    .Y(_09746_));
 sky130_fd_sc_hd__o21ai_4 _19937_ (.A1(_09293_),
    .A2(_09302_),
    .B1(_09740_),
    .Y(_09747_));
 sky130_fd_sc_hd__o221a_1 _19938_ (.A1(_09293_),
    .A2(_09302_),
    .B1(_09737_),
    .B2(net148),
    .C1(_09740_),
    .X(_09748_));
 sky130_fd_sc_hd__o221ai_1 _19939_ (.A1(_09293_),
    .A2(_09302_),
    .B1(_09737_),
    .B2(net148),
    .C1(_09740_),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_1 _19940_ (.A(_09746_),
    .B(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__nor2_1 _19941_ (.A(net25),
    .B(_04353_),
    .Y(_09751_));
 sky130_fd_sc_hd__or3b_1 _19942_ (.A(net44),
    .B(net25),
    .C_N(net55),
    .X(_09752_));
 sky130_fd_sc_hd__a22oi_4 _19943_ (.A1(net25),
    .A2(_04364_),
    .B1(net163),
    .B2(_09751_),
    .Y(_09754_));
 sky130_fd_sc_hd__a31o_4 _19944_ (.A1(_04277_),
    .A2(net163),
    .A3(_04342_),
    .B1(_09272_),
    .X(_09755_));
 sky130_fd_sc_hd__a21oi_4 _19945_ (.A1(net151),
    .A2(net158),
    .B1(_04638_),
    .Y(_09756_));
 sky130_fd_sc_hd__o21ai_1 _19946_ (.A1(_08664_),
    .A2(_08666_),
    .B1(_04627_),
    .Y(_09757_));
 sky130_fd_sc_hd__nor2_2 _19947_ (.A(net319),
    .B(net316),
    .Y(_09758_));
 sky130_fd_sc_hd__or3b_2 _19948_ (.A(net58),
    .B(net319),
    .C_N(net55),
    .X(_09759_));
 sky130_fd_sc_hd__o221ai_4 _19949_ (.A1(_04277_),
    .A2(net316),
    .B1(_09752_),
    .B2(net154),
    .C1(_09273_),
    .Y(_09760_));
 sky130_fd_sc_hd__a21oi_4 _19950_ (.A1(_08670_),
    .A2(_04627_),
    .B1(_09760_),
    .Y(_09761_));
 sky130_fd_sc_hd__o2bb2a_4 _19951_ (.A1_N(net24),
    .A2_N(_04911_),
    .B1(_08209_),
    .B2(_04900_),
    .X(_09762_));
 sky130_fd_sc_hd__a32o_1 _19952_ (.A1(_08204_),
    .A2(net163),
    .A3(_04889_),
    .B1(_04911_),
    .B2(net24),
    .X(_09763_));
 sky130_fd_sc_hd__a21oi_4 _19953_ (.A1(_09757_),
    .A2(_09759_),
    .B1(_09754_),
    .Y(_09765_));
 sky130_fd_sc_hd__o21ai_4 _19954_ (.A1(_09756_),
    .A2(_09758_),
    .B1(_09755_),
    .Y(_09766_));
 sky130_fd_sc_hd__o211ai_4 _19955_ (.A1(_09756_),
    .A2(_09760_),
    .B1(_09762_),
    .C1(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__o21ai_4 _19956_ (.A1(_09761_),
    .A2(_09765_),
    .B1(_09763_),
    .Y(_09768_));
 sky130_fd_sc_hd__o21a_1 _19957_ (.A1(_09760_),
    .A2(_09756_),
    .B1(_09763_),
    .X(_09769_));
 sky130_fd_sc_hd__o21ai_2 _19958_ (.A1(_09760_),
    .A2(_09756_),
    .B1(_09763_),
    .Y(_09770_));
 sky130_fd_sc_hd__o21ai_4 _19959_ (.A1(_09761_),
    .A2(_09765_),
    .B1(_09762_),
    .Y(_09771_));
 sky130_fd_sc_hd__o211ai_4 _19960_ (.A1(_09761_),
    .A2(_09762_),
    .B1(_09771_),
    .C1(_09750_),
    .Y(_09772_));
 sky130_fd_sc_hd__o2111ai_4 _19961_ (.A1(_09747_),
    .A2(_09741_),
    .B1(_09746_),
    .C1(_09767_),
    .D1(_09768_),
    .Y(_09773_));
 sky130_fd_sc_hd__nand3_2 _19962_ (.A(_09750_),
    .B(_09767_),
    .C(_09768_),
    .Y(_09774_));
 sky130_fd_sc_hd__o2111ai_4 _19963_ (.A1(_09747_),
    .A2(_09741_),
    .B1(_09746_),
    .C1(_09770_),
    .D1(_09771_),
    .Y(_09776_));
 sky130_fd_sc_hd__o21ai_4 _19964_ (.A1(_09285_),
    .A2(_09287_),
    .B1(_09309_),
    .Y(_09777_));
 sky130_fd_sc_hd__nand3_2 _19965_ (.A(_09286_),
    .B(_09288_),
    .C(_09307_),
    .Y(_09778_));
 sky130_fd_sc_hd__a22oi_4 _19966_ (.A1(_09774_),
    .A2(_09776_),
    .B1(_09777_),
    .B2(_09307_),
    .Y(_09779_));
 sky130_fd_sc_hd__nand4_4 _19967_ (.A(_09309_),
    .B(_09772_),
    .C(_09773_),
    .D(_09778_),
    .Y(_09780_));
 sky130_fd_sc_hd__a22oi_4 _19968_ (.A1(_09772_),
    .A2(_09773_),
    .B1(_09778_),
    .B2(_09309_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand4_4 _19969_ (.A(_09307_),
    .B(_09774_),
    .C(_09776_),
    .D(_09777_),
    .Y(_09782_));
 sky130_fd_sc_hd__nand4_4 _19970_ (.A(_09730_),
    .B(_09733_),
    .C(_09780_),
    .D(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__inv_2 _19971_ (.A(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__o22ai_4 _19972_ (.A1(_09729_),
    .A2(_09732_),
    .B1(_09779_),
    .B2(_09781_),
    .Y(_09785_));
 sky130_fd_sc_hd__o21ai_1 _19973_ (.A1(_09779_),
    .A2(_09781_),
    .B1(_09734_),
    .Y(_09787_));
 sky130_fd_sc_hd__o211ai_2 _19974_ (.A1(_09729_),
    .A2(_09732_),
    .B1(_09780_),
    .C1(_09782_),
    .Y(_09788_));
 sky130_fd_sc_hd__nand2_2 _19975_ (.A(_09704_),
    .B(_09785_),
    .Y(_09789_));
 sky130_fd_sc_hd__and3_1 _19976_ (.A(_09704_),
    .B(_09783_),
    .C(_09785_),
    .X(_09790_));
 sky130_fd_sc_hd__nand3_2 _19977_ (.A(_09704_),
    .B(_09783_),
    .C(_09785_),
    .Y(_09791_));
 sky130_fd_sc_hd__a21oi_4 _19978_ (.A1(_09783_),
    .A2(_09785_),
    .B1(_09704_),
    .Y(_09792_));
 sky130_fd_sc_hd__o2111ai_4 _19979_ (.A1(_09352_),
    .A2(_09316_),
    .B1(_09315_),
    .C1(_09788_),
    .D1(_09787_),
    .Y(_09793_));
 sky130_fd_sc_hd__o22a_1 _19980_ (.A1(_04135_),
    .A2(_01326_),
    .B1(_05294_),
    .B2(_01304_),
    .X(_09794_));
 sky130_fd_sc_hd__a32o_1 _19981_ (.A1(net182),
    .A2(net179),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net14),
    .X(_09795_));
 sky130_fd_sc_hd__nor2_1 _19982_ (.A(_04146_),
    .B(_12363_),
    .Y(_09796_));
 sky130_fd_sc_hd__a31oi_4 _19983_ (.A1(net178),
    .A2(net177),
    .A3(_12330_),
    .B1(_09796_),
    .Y(_09798_));
 sky130_fd_sc_hd__a31o_1 _19984_ (.A1(net178),
    .A2(net177),
    .A3(_12330_),
    .B1(_09796_),
    .X(_09799_));
 sky130_fd_sc_hd__o211ai_2 _19985_ (.A1(net231),
    .A2(_05927_),
    .B1(net252),
    .C1(_05933_),
    .Y(_09800_));
 sky130_fd_sc_hd__or3_1 _19986_ (.A(net35),
    .B(_04157_),
    .C(_03971_),
    .X(_09801_));
 sky130_fd_sc_hd__o21ai_2 _19987_ (.A1(_04157_),
    .A2(_11804_),
    .B1(_09800_),
    .Y(_09802_));
 sky130_fd_sc_hd__a21oi_2 _19988_ (.A1(_09800_),
    .A2(_09801_),
    .B1(_09798_),
    .Y(_09803_));
 sky130_fd_sc_hd__nand2_1 _19989_ (.A(_09799_),
    .B(_09802_),
    .Y(_09804_));
 sky130_fd_sc_hd__o311a_2 _19990_ (.A1(_03971_),
    .A2(net35),
    .A3(_04157_),
    .B1(_09800_),
    .C1(_09798_),
    .X(_09805_));
 sky130_fd_sc_hd__o221ai_4 _19991_ (.A1(_04157_),
    .A2(_11804_),
    .B1(net155),
    .B2(_11782_),
    .C1(_09798_),
    .Y(_09806_));
 sky130_fd_sc_hd__a21oi_2 _19992_ (.A1(_09804_),
    .A2(_09806_),
    .B1(_09795_),
    .Y(_09807_));
 sky130_fd_sc_hd__nor3_2 _19993_ (.A(_09794_),
    .B(_09803_),
    .C(_09805_),
    .Y(_09809_));
 sky130_fd_sc_hd__nand3_1 _19994_ (.A(_09795_),
    .B(_09804_),
    .C(_09806_),
    .Y(_09810_));
 sky130_fd_sc_hd__nor2_1 _19995_ (.A(_09807_),
    .B(_09809_),
    .Y(_09811_));
 sky130_fd_sc_hd__and3_1 _19996_ (.A(_03971_),
    .B(net17),
    .C(net64),
    .X(_09812_));
 sky130_fd_sc_hd__and3_1 _19997_ (.A(net201),
    .B(_06221_),
    .C(net289),
    .X(_09813_));
 sky130_fd_sc_hd__a31oi_4 _19998_ (.A1(net201),
    .A2(_06221_),
    .A3(net289),
    .B1(_09812_),
    .Y(_09814_));
 sky130_fd_sc_hd__o211ai_2 _19999_ (.A1(net175),
    .A2(_06451_),
    .B1(net291),
    .C1(net199),
    .Y(_09815_));
 sky130_fd_sc_hd__nor2_1 _20000_ (.A(_04179_),
    .B(_08283_),
    .Y(_09816_));
 sky130_fd_sc_hd__or3b_1 _20001_ (.A(net64),
    .B(_04179_),
    .C_N(net63),
    .X(_09817_));
 sky130_fd_sc_hd__a31oi_4 _20002_ (.A1(net199),
    .A2(net172),
    .A3(net291),
    .B1(_09816_),
    .Y(_09818_));
 sky130_fd_sc_hd__a31o_1 _20003_ (.A1(net199),
    .A2(net172),
    .A3(net291),
    .B1(_09816_),
    .X(_09820_));
 sky130_fd_sc_hd__nor2_1 _20004_ (.A(_04201_),
    .B(_07691_),
    .Y(_09821_));
 sky130_fd_sc_hd__or3_1 _20005_ (.A(net63),
    .B(_04201_),
    .C(_03927_),
    .X(_09822_));
 sky130_fd_sc_hd__o2111ai_4 _20006_ (.A1(net175),
    .A2(_06759_),
    .B1(net63),
    .C1(net195),
    .D1(_03927_),
    .Y(_09823_));
 sky130_fd_sc_hd__o31a_1 _20007_ (.A1(net189),
    .A2(_07669_),
    .A3(_06756_),
    .B1(_09822_),
    .X(_09824_));
 sky130_fd_sc_hd__a31o_1 _20008_ (.A1(net195),
    .A2(net171),
    .A3(_07658_),
    .B1(_09821_),
    .X(_09825_));
 sky130_fd_sc_hd__o311a_1 _20009_ (.A1(_03927_),
    .A2(net63),
    .A3(_04201_),
    .B1(_09823_),
    .C1(_09818_),
    .X(_09826_));
 sky130_fd_sc_hd__a21oi_1 _20010_ (.A1(_09822_),
    .A2(_09823_),
    .B1(_09818_),
    .Y(_09827_));
 sky130_fd_sc_hd__a22o_2 _20011_ (.A1(_09815_),
    .A2(_09817_),
    .B1(_09822_),
    .B2(_09823_),
    .X(_09828_));
 sky130_fd_sc_hd__o2111ai_4 _20012_ (.A1(_04201_),
    .A2(_07691_),
    .B1(_09814_),
    .C1(_09823_),
    .D1(_09818_),
    .Y(_09829_));
 sky130_fd_sc_hd__o21a_1 _20013_ (.A1(_09818_),
    .A2(_09824_),
    .B1(_09814_),
    .X(_09831_));
 sky130_fd_sc_hd__o22a_1 _20014_ (.A1(_09812_),
    .A2(_09813_),
    .B1(_09820_),
    .B2(_09825_),
    .X(_09832_));
 sky130_fd_sc_hd__o22ai_2 _20015_ (.A1(_09812_),
    .A2(_09813_),
    .B1(_09820_),
    .B2(_09825_),
    .Y(_09833_));
 sky130_fd_sc_hd__a32o_1 _20016_ (.A1(_09815_),
    .A2(_09817_),
    .A3(_09824_),
    .B1(_09828_),
    .B2(_09814_),
    .X(_09834_));
 sky130_fd_sc_hd__o211ai_4 _20017_ (.A1(_09818_),
    .A2(_09824_),
    .B1(_09829_),
    .C1(_09833_),
    .Y(_09835_));
 sky130_fd_sc_hd__a221o_1 _20018_ (.A1(_09815_),
    .A2(_09817_),
    .B1(_09822_),
    .B2(_09823_),
    .C1(_09814_),
    .X(_09836_));
 sky130_fd_sc_hd__a22oi_4 _20019_ (.A1(_09368_),
    .A2(_09377_),
    .B1(_09835_),
    .B2(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__a22o_1 _20020_ (.A1(_09368_),
    .A2(_09377_),
    .B1(_09835_),
    .B2(_09836_),
    .X(_09838_));
 sky130_fd_sc_hd__o2111a_1 _20021_ (.A1(_09828_),
    .A2(_09814_),
    .B1(_09377_),
    .C1(_09368_),
    .D1(_09835_),
    .X(_09839_));
 sky130_fd_sc_hd__o2111ai_4 _20022_ (.A1(_09828_),
    .A2(_09814_),
    .B1(_09377_),
    .C1(_09368_),
    .D1(_09835_),
    .Y(_09840_));
 sky130_fd_sc_hd__nand3b_2 _20023_ (.A_N(_09807_),
    .B(_09810_),
    .C(_09840_),
    .Y(_09842_));
 sky130_fd_sc_hd__nand3_1 _20024_ (.A(_09838_),
    .B(_09840_),
    .C(_09811_),
    .Y(_09843_));
 sky130_fd_sc_hd__o22ai_4 _20025_ (.A1(_09807_),
    .A2(_09809_),
    .B1(_09837_),
    .B2(_09839_),
    .Y(_09844_));
 sky130_fd_sc_hd__o21ai_1 _20026_ (.A1(_09837_),
    .A2(_09842_),
    .B1(_09844_),
    .Y(_09845_));
 sky130_fd_sc_hd__o31a_1 _20027_ (.A1(_09333_),
    .A2(_09335_),
    .A3(_09338_),
    .B1(_09318_),
    .X(_09846_));
 sky130_fd_sc_hd__o21ai_2 _20028_ (.A1(_09318_),
    .A2(_09340_),
    .B1(_09342_),
    .Y(_09847_));
 sky130_fd_sc_hd__o21a_1 _20029_ (.A1(_09318_),
    .A2(_09340_),
    .B1(_09342_),
    .X(_09848_));
 sky130_fd_sc_hd__a21oi_1 _20030_ (.A1(_09843_),
    .A2(_09844_),
    .B1(_09847_),
    .Y(_09849_));
 sky130_fd_sc_hd__o2bb2ai_2 _20031_ (.A1_N(_09843_),
    .A2_N(_09844_),
    .B1(_09846_),
    .B2(_09340_),
    .Y(_09850_));
 sky130_fd_sc_hd__o211a_2 _20032_ (.A1(_09837_),
    .A2(_09842_),
    .B1(_09844_),
    .C1(_09847_),
    .X(_09851_));
 sky130_fd_sc_hd__o211ai_4 _20033_ (.A1(_09837_),
    .A2(_09842_),
    .B1(_09844_),
    .C1(_09847_),
    .Y(_09853_));
 sky130_fd_sc_hd__o2bb2a_2 _20034_ (.A1_N(_09379_),
    .A2_N(_09405_),
    .B1(_09849_),
    .B2(_09851_),
    .X(_09854_));
 sky130_fd_sc_hd__a22o_2 _20035_ (.A1(_09379_),
    .A2(_09405_),
    .B1(_09850_),
    .B2(_09853_),
    .X(_09855_));
 sky130_fd_sc_hd__a21oi_2 _20036_ (.A1(_09845_),
    .A2(_09848_),
    .B1(_09406_),
    .Y(_09856_));
 sky130_fd_sc_hd__o31a_2 _20037_ (.A1(_09340_),
    .A2(_09845_),
    .A3(_09846_),
    .B1(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__nand4_4 _20038_ (.A(_09379_),
    .B(_09405_),
    .C(_09850_),
    .D(_09853_),
    .Y(_09858_));
 sky130_fd_sc_hd__nand2_1 _20039_ (.A(_09855_),
    .B(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__o221ai_4 _20040_ (.A1(_09784_),
    .A2(_09789_),
    .B1(_09854_),
    .B2(_09857_),
    .C1(_09793_),
    .Y(_09860_));
 sky130_fd_sc_hd__a21o_1 _20041_ (.A1(_09791_),
    .A2(_09793_),
    .B1(_09859_),
    .X(_09861_));
 sky130_fd_sc_hd__o2bb2ai_4 _20042_ (.A1_N(_09791_),
    .A2_N(_09793_),
    .B1(_09854_),
    .B2(_09857_),
    .Y(_09862_));
 sky130_fd_sc_hd__nand3_2 _20043_ (.A(_09793_),
    .B(_09855_),
    .C(_09858_),
    .Y(_09864_));
 sky130_fd_sc_hd__nand4_2 _20044_ (.A(_09791_),
    .B(_09793_),
    .C(_09855_),
    .D(_09858_),
    .Y(_09865_));
 sky130_fd_sc_hd__a22oi_4 _20045_ (.A1(_09362_),
    .A2(_09702_),
    .B1(_09862_),
    .B2(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__o211ai_4 _20046_ (.A1(_09361_),
    .A2(_09701_),
    .B1(_09860_),
    .C1(_09861_),
    .Y(_09867_));
 sky130_fd_sc_hd__o211a_1 _20047_ (.A1(_09790_),
    .A2(_09864_),
    .B1(_09703_),
    .C1(_09862_),
    .X(_09868_));
 sky130_fd_sc_hd__o2111ai_4 _20048_ (.A1(_09790_),
    .A2(_09864_),
    .B1(_09862_),
    .C1(_09362_),
    .D1(_09702_),
    .Y(_09869_));
 sky130_fd_sc_hd__a21oi_1 _20049_ (.A1(_09210_),
    .A2(_09211_),
    .B1(_09247_),
    .Y(_09870_));
 sky130_fd_sc_hd__a32o_1 _20050_ (.A1(_09242_),
    .A2(_09243_),
    .A3(_09244_),
    .B1(_09249_),
    .B2(_09212_),
    .X(_09871_));
 sky130_fd_sc_hd__o21ai_1 _20051_ (.A1(_09418_),
    .A2(_09411_),
    .B1(_09415_),
    .Y(_09872_));
 sky130_fd_sc_hd__a21oi_2 _20052_ (.A1(_09412_),
    .A2(_09417_),
    .B1(_09414_),
    .Y(_09873_));
 sky130_fd_sc_hd__o32a_2 _20053_ (.A1(_04896_),
    .A2(_03957_),
    .A3(_03951_),
    .B1(_04048_),
    .B2(_04898_),
    .X(_09875_));
 sky130_fd_sc_hd__nand3_2 _20054_ (.A(net229),
    .B(net228),
    .C(net279),
    .Y(_09876_));
 sky130_fd_sc_hd__or3b_1 _20055_ (.A(_04059_),
    .B(net42),
    .C_N(net41),
    .X(_09877_));
 sky130_fd_sc_hd__nand3_2 _20056_ (.A(net222),
    .B(net280),
    .C(net188),
    .Y(_09878_));
 sky130_fd_sc_hd__or3b_2 _20057_ (.A(net41),
    .B(_04069_),
    .C_N(net40),
    .X(_09879_));
 sky130_fd_sc_hd__a22oi_2 _20058_ (.A1(_09876_),
    .A2(_09877_),
    .B1(_09878_),
    .B2(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__a22o_1 _20059_ (.A1(_09876_),
    .A2(_09877_),
    .B1(_09878_),
    .B2(_09879_),
    .X(_09881_));
 sky130_fd_sc_hd__o2111a_1 _20060_ (.A1(_04059_),
    .A2(_04483_),
    .B1(_09876_),
    .C1(_09878_),
    .D1(_09879_),
    .X(_09882_));
 sky130_fd_sc_hd__o2111ai_2 _20061_ (.A1(_04059_),
    .A2(_04483_),
    .B1(_09876_),
    .C1(_09878_),
    .D1(_09879_),
    .Y(_09883_));
 sky130_fd_sc_hd__o21ai_2 _20062_ (.A1(_09880_),
    .A2(_09882_),
    .B1(_09875_),
    .Y(_09884_));
 sky130_fd_sc_hd__nand3b_2 _20063_ (.A_N(_09875_),
    .B(_09881_),
    .C(_09883_),
    .Y(_09886_));
 sky130_fd_sc_hd__nand3_1 _20064_ (.A(_09881_),
    .B(_09883_),
    .C(_09875_),
    .Y(_09887_));
 sky130_fd_sc_hd__o21bai_1 _20065_ (.A1(_09880_),
    .A2(_09882_),
    .B1_N(_09875_),
    .Y(_09888_));
 sky130_fd_sc_hd__o2111ai_4 _20066_ (.A1(_09183_),
    .A2(_09186_),
    .B1(_09191_),
    .C1(_09887_),
    .D1(_09888_),
    .Y(_09889_));
 sky130_fd_sc_hd__o211a_1 _20067_ (.A1(_09187_),
    .A2(_09190_),
    .B1(_09884_),
    .C1(_09886_),
    .X(_09890_));
 sky130_fd_sc_hd__o211ai_4 _20068_ (.A1(_09187_),
    .A2(_09190_),
    .B1(_09884_),
    .C1(_09886_),
    .Y(_09891_));
 sky130_fd_sc_hd__a41o_1 _20069_ (.A1(net307),
    .A2(net293),
    .A3(net288),
    .A4(_00635_),
    .B1(_05226_),
    .X(_09892_));
 sky130_fd_sc_hd__o32a_4 _20070_ (.A1(_04015_),
    .A2(_04124_),
    .A3(net46),
    .B1(_00614_),
    .B2(_09892_),
    .X(_09893_));
 sky130_fd_sc_hd__o2111ai_4 _20071_ (.A1(net253),
    .A2(_02442_),
    .B1(net45),
    .C1(_02421_),
    .D1(_04102_),
    .Y(_09894_));
 sky130_fd_sc_hd__or3_1 _20072_ (.A(net45),
    .B(_04102_),
    .C(_04026_),
    .X(_09895_));
 sky130_fd_sc_hd__a21oi_2 _20073_ (.A1(_09894_),
    .A2(_09895_),
    .B1(_09893_),
    .Y(_09897_));
 sky130_fd_sc_hd__o311a_1 _20074_ (.A1(_04026_),
    .A2(_04102_),
    .A3(net45),
    .B1(_09894_),
    .C1(_09893_),
    .X(_09898_));
 sky130_fd_sc_hd__o211ai_1 _20075_ (.A1(_04026_),
    .A2(_04989_),
    .B1(_09894_),
    .C1(_09893_),
    .Y(_09899_));
 sky130_fd_sc_hd__or3b_1 _20076_ (.A(_04004_),
    .B(net47),
    .C_N(net46),
    .X(_09900_));
 sky130_fd_sc_hd__o211ai_2 _20077_ (.A1(_11387_),
    .A2(_12988_),
    .B1(_05462_),
    .C1(net234),
    .Y(_09901_));
 sky130_fd_sc_hd__o21a_1 _20078_ (.A1(_04004_),
    .A2(_05465_),
    .B1(_09901_),
    .X(_09902_));
 sky130_fd_sc_hd__a32o_1 _20079_ (.A1(net234),
    .A2(net251),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net4),
    .X(_09903_));
 sky130_fd_sc_hd__nand3b_1 _20080_ (.A_N(_09897_),
    .B(_09899_),
    .C(_09902_),
    .Y(_09904_));
 sky130_fd_sc_hd__o21ai_1 _20081_ (.A1(_09897_),
    .A2(_09898_),
    .B1(_09903_),
    .Y(_09905_));
 sky130_fd_sc_hd__o211a_1 _20082_ (.A1(_09897_),
    .A2(_09898_),
    .B1(_09900_),
    .C1(_09901_),
    .X(_09906_));
 sky130_fd_sc_hd__a211oi_1 _20083_ (.A1(_09900_),
    .A2(_09901_),
    .B1(_09897_),
    .C1(_09898_),
    .Y(_09908_));
 sky130_fd_sc_hd__nand2_1 _20084_ (.A(_09904_),
    .B(_09905_),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_2 _20085_ (.A(_09889_),
    .B(_09909_),
    .Y(_09910_));
 sky130_fd_sc_hd__and3_1 _20086_ (.A(_09889_),
    .B(_09891_),
    .C(_09909_),
    .X(_09911_));
 sky130_fd_sc_hd__a21o_1 _20087_ (.A1(_09889_),
    .A2(_09891_),
    .B1(_09909_),
    .X(_09912_));
 sky130_fd_sc_hd__inv_2 _20088_ (.A(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__o21ai_2 _20089_ (.A1(_09890_),
    .A2(_09910_),
    .B1(_09912_),
    .Y(_09914_));
 sky130_fd_sc_hd__a21oi_1 _20090_ (.A1(_09223_),
    .A2(_09229_),
    .B1(_09224_),
    .Y(_09915_));
 sky130_fd_sc_hd__nand3_4 _20091_ (.A(net214),
    .B(net285),
    .C(net184),
    .Y(_09916_));
 sky130_fd_sc_hd__nor2_1 _20092_ (.A(_04091_),
    .B(_03737_),
    .Y(_09917_));
 sky130_fd_sc_hd__or3_2 _20093_ (.A(net39),
    .B(_04091_),
    .C(_04037_),
    .X(_09919_));
 sky130_fd_sc_hd__and3_1 _20094_ (.A(_04037_),
    .B(net13),
    .C(net37),
    .X(_09920_));
 sky130_fd_sc_hd__or3b_2 _20095_ (.A(net38),
    .B(_04113_),
    .C_N(net37),
    .X(_09921_));
 sky130_fd_sc_hd__o311a_1 _20096_ (.A1(net11),
    .A2(_04557_),
    .A3(net208),
    .B1(_02858_),
    .C1(net211),
    .X(_09922_));
 sky130_fd_sc_hd__o211ai_4 _20097_ (.A1(_04787_),
    .A2(net208),
    .B1(_02858_),
    .C1(net211),
    .Y(_09923_));
 sky130_fd_sc_hd__a22oi_4 _20098_ (.A1(_09916_),
    .A2(_09919_),
    .B1(_09921_),
    .B2(_09923_),
    .Y(_09924_));
 sky130_fd_sc_hd__o2bb2ai_4 _20099_ (.A1_N(_09916_),
    .A2_N(_09919_),
    .B1(_09920_),
    .B2(_09922_),
    .Y(_09925_));
 sky130_fd_sc_hd__o211ai_2 _20100_ (.A1(_04113_),
    .A2(_02891_),
    .B1(_09916_),
    .C1(_09923_),
    .Y(_09926_));
 sky130_fd_sc_hd__o2111a_1 _20101_ (.A1(_04091_),
    .A2(_03737_),
    .B1(_09916_),
    .C1(_09921_),
    .D1(_09923_),
    .X(_09927_));
 sky130_fd_sc_hd__o2111ai_1 _20102_ (.A1(_04091_),
    .A2(_03737_),
    .B1(_09916_),
    .C1(_09921_),
    .D1(_09923_),
    .Y(_09928_));
 sky130_fd_sc_hd__a32o_2 _20103_ (.A1(net218),
    .A2(net186),
    .A3(net281),
    .B1(_04217_),
    .B2(net10),
    .X(_09930_));
 sky130_fd_sc_hd__a21oi_1 _20104_ (.A1(_09925_),
    .A2(_09928_),
    .B1(_09930_),
    .Y(_09931_));
 sky130_fd_sc_hd__o21bai_2 _20105_ (.A1(_09924_),
    .A2(_09927_),
    .B1_N(_09930_),
    .Y(_09932_));
 sky130_fd_sc_hd__o211a_2 _20106_ (.A1(_09917_),
    .A2(_09926_),
    .B1(_09930_),
    .C1(_09925_),
    .X(_09933_));
 sky130_fd_sc_hd__o211ai_4 _20107_ (.A1(_09917_),
    .A2(_09926_),
    .B1(_09930_),
    .C1(_09925_),
    .Y(_09934_));
 sky130_fd_sc_hd__a22oi_2 _20108_ (.A1(_09393_),
    .A2(_09397_),
    .B1(_09932_),
    .B2(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__o2bb2ai_2 _20109_ (.A1_N(_09393_),
    .A2_N(_09397_),
    .B1(_09931_),
    .B2(_09933_),
    .Y(_09936_));
 sky130_fd_sc_hd__o21ai_2 _20110_ (.A1(_09394_),
    .A2(_09398_),
    .B1(_09932_),
    .Y(_09937_));
 sky130_fd_sc_hd__o211a_2 _20111_ (.A1(_09394_),
    .A2(_09398_),
    .B1(_09932_),
    .C1(_09934_),
    .X(_09938_));
 sky130_fd_sc_hd__o211ai_1 _20112_ (.A1(_09394_),
    .A2(_09398_),
    .B1(_09932_),
    .C1(_09934_),
    .Y(_09939_));
 sky130_fd_sc_hd__a21boi_1 _20113_ (.A1(_09936_),
    .A2(_09939_),
    .B1_N(_09915_),
    .Y(_09941_));
 sky130_fd_sc_hd__o21ai_2 _20114_ (.A1(_09935_),
    .A2(_09938_),
    .B1(_09915_),
    .Y(_09942_));
 sky130_fd_sc_hd__o21ai_1 _20115_ (.A1(_09224_),
    .A2(_09232_),
    .B1(_09936_),
    .Y(_09943_));
 sky130_fd_sc_hd__o221a_2 _20116_ (.A1(_09224_),
    .A2(_09232_),
    .B1(_09933_),
    .B2(_09937_),
    .C1(_09936_),
    .X(_09944_));
 sky130_fd_sc_hd__o221ai_4 _20117_ (.A1(_09224_),
    .A2(_09232_),
    .B1(_09933_),
    .B2(_09937_),
    .C1(_09936_),
    .Y(_09945_));
 sky130_fd_sc_hd__o22ai_4 _20118_ (.A1(_09232_),
    .A2(_09238_),
    .B1(_09039_),
    .B2(_09235_),
    .Y(_09946_));
 sky130_fd_sc_hd__o22a_1 _20119_ (.A1(_09232_),
    .A2(_09238_),
    .B1(_09039_),
    .B2(_09235_),
    .X(_09947_));
 sky130_fd_sc_hd__a21oi_4 _20120_ (.A1(_09942_),
    .A2(_09945_),
    .B1(_09946_),
    .Y(_09948_));
 sky130_fd_sc_hd__o21ai_1 _20121_ (.A1(_09941_),
    .A2(_09944_),
    .B1(_09947_),
    .Y(_09949_));
 sky130_fd_sc_hd__o211a_1 _20122_ (.A1(_09938_),
    .A2(_09943_),
    .B1(_09942_),
    .C1(_09946_),
    .X(_09950_));
 sky130_fd_sc_hd__o211ai_2 _20123_ (.A1(_09938_),
    .A2(_09943_),
    .B1(_09942_),
    .C1(_09946_),
    .Y(_09952_));
 sky130_fd_sc_hd__a31o_1 _20124_ (.A1(_09942_),
    .A2(_09946_),
    .A3(_09945_),
    .B1(_09914_),
    .X(_09953_));
 sky130_fd_sc_hd__o2111ai_2 _20125_ (.A1(_09890_),
    .A2(_09910_),
    .B1(_09912_),
    .C1(_09949_),
    .D1(_09952_),
    .Y(_09954_));
 sky130_fd_sc_hd__o22ai_4 _20126_ (.A1(_09911_),
    .A2(_09913_),
    .B1(_09948_),
    .B2(_09950_),
    .Y(_09955_));
 sky130_fd_sc_hd__o211a_1 _20127_ (.A1(_09941_),
    .A2(_09944_),
    .B1(_09947_),
    .C1(_09914_),
    .X(_09956_));
 sky130_fd_sc_hd__o32a_2 _20128_ (.A1(_09941_),
    .A2(_09944_),
    .A3(_09947_),
    .B1(_09913_),
    .B2(_09911_),
    .X(_09957_));
 sky130_fd_sc_hd__o21ai_2 _20129_ (.A1(_09914_),
    .A2(_09948_),
    .B1(_09952_),
    .Y(_09958_));
 sky130_fd_sc_hd__o21ai_1 _20130_ (.A1(_09948_),
    .A2(_09953_),
    .B1(_09955_),
    .Y(_09959_));
 sky130_fd_sc_hd__o221a_1 _20131_ (.A1(_09948_),
    .A2(_09953_),
    .B1(_09414_),
    .B2(_09421_),
    .C1(_09955_),
    .X(_09960_));
 sky130_fd_sc_hd__o221ai_4 _20132_ (.A1(_09948_),
    .A2(_09953_),
    .B1(_09414_),
    .B2(_09421_),
    .C1(_09955_),
    .Y(_09961_));
 sky130_fd_sc_hd__a21oi_2 _20133_ (.A1(_09954_),
    .A2(_09955_),
    .B1(_09872_),
    .Y(_09963_));
 sky130_fd_sc_hd__o221ai_1 _20134_ (.A1(_09914_),
    .A2(_09952_),
    .B1(_09956_),
    .B2(_09958_),
    .C1(_09873_),
    .Y(_09964_));
 sky130_fd_sc_hd__a2bb2oi_2 _20135_ (.A1_N(_09247_),
    .A2_N(_09253_),
    .B1(_09873_),
    .B2(_09959_),
    .Y(_09965_));
 sky130_fd_sc_hd__o21ai_2 _20136_ (.A1(_09873_),
    .A2(_09959_),
    .B1(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__a2bb2oi_1 _20137_ (.A1_N(_09245_),
    .A2_N(_09870_),
    .B1(_09961_),
    .B2(_09964_),
    .Y(_09967_));
 sky130_fd_sc_hd__o21ai_2 _20138_ (.A1(_09960_),
    .A2(_09963_),
    .B1(_09871_),
    .Y(_09968_));
 sky130_fd_sc_hd__a21oi_2 _20139_ (.A1(_09961_),
    .A2(_09965_),
    .B1(_09967_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand2_2 _20140_ (.A(_09966_),
    .B(_09968_),
    .Y(_09970_));
 sky130_fd_sc_hd__nand3_4 _20141_ (.A(_09867_),
    .B(_09869_),
    .C(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__o21ai_4 _20142_ (.A1(_09866_),
    .A2(_09868_),
    .B1(_09969_),
    .Y(_09972_));
 sky130_fd_sc_hd__o21ai_1 _20143_ (.A1(_09866_),
    .A2(_09868_),
    .B1(_09970_),
    .Y(_09974_));
 sky130_fd_sc_hd__nand4_1 _20144_ (.A(_09867_),
    .B(_09869_),
    .C(_09966_),
    .D(_09968_),
    .Y(_09975_));
 sky130_fd_sc_hd__a22oi_1 _20145_ (.A1(_09433_),
    .A2(_09438_),
    .B1(_09974_),
    .B2(_09975_),
    .Y(_09976_));
 sky130_fd_sc_hd__o2111ai_4 _20146_ (.A1(_09264_),
    .A2(_09432_),
    .B1(_09436_),
    .C1(_09971_),
    .D1(_09972_),
    .Y(_09977_));
 sky130_fd_sc_hd__a2bb2oi_4 _20147_ (.A1_N(_09434_),
    .A2_N(_09439_),
    .B1(_09971_),
    .B2(_09972_),
    .Y(_09978_));
 sky130_fd_sc_hd__nand3_1 _20148_ (.A(_09974_),
    .B(_09975_),
    .C(_09699_),
    .Y(_09979_));
 sky130_fd_sc_hd__o211ai_2 _20149_ (.A1(_09691_),
    .A2(_09695_),
    .B1(_09977_),
    .C1(_09979_),
    .Y(_09980_));
 sky130_fd_sc_hd__a21o_1 _20150_ (.A1(_09977_),
    .A2(_09979_),
    .B1(_09697_),
    .X(_09981_));
 sky130_fd_sc_hd__a31oi_2 _20151_ (.A1(_09700_),
    .A2(_09971_),
    .A3(_09972_),
    .B1(_09697_),
    .Y(_09982_));
 sky130_fd_sc_hd__nand2_1 _20152_ (.A(_09977_),
    .B(_09696_),
    .Y(_09983_));
 sky130_fd_sc_hd__o22ai_2 _20153_ (.A1(_09691_),
    .A2(_09695_),
    .B1(_09976_),
    .B2(_09978_),
    .Y(_09985_));
 sky130_fd_sc_hd__o21ai_1 _20154_ (.A1(_09978_),
    .A2(_09983_),
    .B1(_09985_),
    .Y(_09986_));
 sky130_fd_sc_hd__o211ai_4 _20155_ (.A1(_09978_),
    .A2(_09983_),
    .B1(_09590_),
    .C1(_09985_),
    .Y(_09987_));
 sky130_fd_sc_hd__o211a_1 _20156_ (.A1(_09447_),
    .A2(_09589_),
    .B1(_09980_),
    .C1(_09981_),
    .X(_09988_));
 sky130_fd_sc_hd__o211ai_4 _20157_ (.A1(_09447_),
    .A2(_09589_),
    .B1(_09980_),
    .C1(_09981_),
    .Y(_09989_));
 sky130_fd_sc_hd__o311a_1 _20158_ (.A1(_08761_),
    .A2(_08795_),
    .A3(_08799_),
    .B1(_08835_),
    .C1(_09546_),
    .X(_09990_));
 sky130_fd_sc_hd__a21oi_1 _20159_ (.A1(_08805_),
    .A2(_08835_),
    .B1(_09542_),
    .Y(_09991_));
 sky130_fd_sc_hd__o21ai_1 _20160_ (.A1(_09547_),
    .A2(_09991_),
    .B1(_09989_),
    .Y(_09992_));
 sky130_fd_sc_hd__o211ai_1 _20161_ (.A1(_09547_),
    .A2(_09991_),
    .B1(_09989_),
    .C1(_09987_),
    .Y(_09993_));
 sky130_fd_sc_hd__o2bb2ai_1 _20162_ (.A1_N(_09987_),
    .A2_N(_09989_),
    .B1(_09990_),
    .B2(_09542_),
    .Y(_09994_));
 sky130_fd_sc_hd__o2bb2ai_1 _20163_ (.A1_N(_09987_),
    .A2_N(_09989_),
    .B1(_09991_),
    .B2(_09547_),
    .Y(_09996_));
 sky130_fd_sc_hd__o2111ai_4 _20164_ (.A1(_09548_),
    .A2(_09542_),
    .B1(_09546_),
    .C1(_09987_),
    .D1(_09989_),
    .Y(_09997_));
 sky130_fd_sc_hd__a31oi_2 _20165_ (.A1(_09134_),
    .A2(_09554_),
    .A3(_09558_),
    .B1(_09563_),
    .Y(_09998_));
 sky130_fd_sc_hd__o22ai_1 _20166_ (.A1(_09557_),
    .A2(_09561_),
    .B1(_09564_),
    .B2(_09559_),
    .Y(_09999_));
 sky130_fd_sc_hd__o211ai_4 _20167_ (.A1(_09559_),
    .A2(_09998_),
    .B1(_09997_),
    .C1(_09996_),
    .Y(_10000_));
 sky130_fd_sc_hd__inv_2 _20168_ (.A(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__nand3_2 _20169_ (.A(_09993_),
    .B(_09994_),
    .C(_09999_),
    .Y(_10002_));
 sky130_fd_sc_hd__nor2_1 _20170_ (.A(_09499_),
    .B(_09531_),
    .Y(_10003_));
 sky130_fd_sc_hd__nor2_1 _20171_ (.A(_09498_),
    .B(_09530_),
    .Y(_10004_));
 sky130_fd_sc_hd__o21ai_1 _20172_ (.A1(_09531_),
    .A2(_09535_),
    .B1(_10000_),
    .Y(_10005_));
 sky130_fd_sc_hd__o211ai_1 _20173_ (.A1(_09531_),
    .A2(_09535_),
    .B1(_10000_),
    .C1(_10002_),
    .Y(_10007_));
 sky130_fd_sc_hd__inv_2 _20174_ (.A(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__o2bb2ai_1 _20175_ (.A1_N(_10000_),
    .A2_N(_10002_),
    .B1(_10003_),
    .B2(_09530_),
    .Y(_10009_));
 sky130_fd_sc_hd__o2bb2ai_1 _20176_ (.A1_N(_10000_),
    .A2_N(_10002_),
    .B1(_10004_),
    .B2(_09531_),
    .Y(_10010_));
 sky130_fd_sc_hd__o2111ai_1 _20177_ (.A1(_09533_),
    .A2(_09498_),
    .B1(_09532_),
    .C1(_10000_),
    .D1(_10002_),
    .Y(_10011_));
 sky130_fd_sc_hd__nand4_2 _20178_ (.A(_09572_),
    .B(_09579_),
    .C(_10010_),
    .D(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__o21ai_2 _20179_ (.A1(_09571_),
    .A2(_09577_),
    .B1(_10009_),
    .Y(_10013_));
 sky130_fd_sc_hd__o21ai_1 _20180_ (.A1(_10008_),
    .A2(_10013_),
    .B1(_10012_),
    .Y(_10014_));
 sky130_fd_sc_hd__a21o_1 _20181_ (.A1(_09160_),
    .A2(_09585_),
    .B1(_09583_),
    .X(_10015_));
 sky130_fd_sc_hd__nand4_1 _20182_ (.A(_09159_),
    .B(_09160_),
    .C(_09584_),
    .D(_09585_),
    .Y(_10016_));
 sky130_fd_sc_hd__o21ai_1 _20183_ (.A1(_10016_),
    .A2(_09170_),
    .B1(_10015_),
    .Y(_10018_));
 sky130_fd_sc_hd__xnor2_1 _20184_ (.A(_10014_),
    .B(_10018_),
    .Y(net92));
 sky130_fd_sc_hd__o211a_1 _20185_ (.A1(_09533_),
    .A2(_09498_),
    .B1(_09532_),
    .C1(_10002_),
    .X(_10019_));
 sky130_fd_sc_hd__nand2_1 _20186_ (.A(_10002_),
    .B(_10005_),
    .Y(_10020_));
 sky130_fd_sc_hd__nor2_1 _20187_ (.A(_09641_),
    .B(_09670_),
    .Y(_10021_));
 sky130_fd_sc_hd__a31o_1 _20188_ (.A1(_09664_),
    .A2(_09666_),
    .A3(_09669_),
    .B1(_09674_),
    .X(_10022_));
 sky130_fd_sc_hd__o211a_1 _20189_ (.A1(_09548_),
    .A2(_09542_),
    .B1(_09546_),
    .C1(_09987_),
    .X(_10023_));
 sky130_fd_sc_hd__o31ai_1 _20190_ (.A1(_09447_),
    .A2(_09589_),
    .A3(_09986_),
    .B1(_09992_),
    .Y(_10024_));
 sky130_fd_sc_hd__o21ai_2 _20191_ (.A1(_09683_),
    .A2(_09685_),
    .B1(_09694_),
    .Y(_10025_));
 sky130_fd_sc_hd__a21oi_1 _20192_ (.A1(_09977_),
    .A2(_09696_),
    .B1(_09978_),
    .Y(_10026_));
 sky130_fd_sc_hd__nand2_1 _20193_ (.A(_09601_),
    .B(_09603_),
    .Y(_10028_));
 sky130_fd_sc_hd__a32o_1 _20194_ (.A1(net255),
    .A2(_09698_),
    .A3(net273),
    .B1(_06326_),
    .B2(net2),
    .X(_10029_));
 sky130_fd_sc_hd__o211ai_4 _20195_ (.A1(net259),
    .A2(_11387_),
    .B1(net274),
    .C1(_11354_),
    .Y(_10030_));
 sky130_fd_sc_hd__or3b_2 _20196_ (.A(_03982_),
    .B(net49),
    .C_N(net48),
    .X(_10031_));
 sky130_fd_sc_hd__o211ai_4 _20197_ (.A1(_11387_),
    .A2(_12988_),
    .B1(net275),
    .C1(net234),
    .Y(_10032_));
 sky130_fd_sc_hd__or3b_2 _20198_ (.A(_04004_),
    .B(net48),
    .C_N(net47),
    .X(_10033_));
 sky130_fd_sc_hd__a22oi_2 _20199_ (.A1(_10030_),
    .A2(_10031_),
    .B1(_10032_),
    .B2(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__a22o_1 _20200_ (.A1(_10030_),
    .A2(_10031_),
    .B1(_10032_),
    .B2(_10033_),
    .X(_10035_));
 sky130_fd_sc_hd__and4_1 _20201_ (.A(_10030_),
    .B(_10031_),
    .C(_10032_),
    .D(_10033_),
    .X(_10036_));
 sky130_fd_sc_hd__nand4_1 _20202_ (.A(_10030_),
    .B(_10031_),
    .C(_10032_),
    .D(_10033_),
    .Y(_10037_));
 sky130_fd_sc_hd__o21bai_1 _20203_ (.A1(_10034_),
    .A2(_10036_),
    .B1_N(_10029_),
    .Y(_10039_));
 sky130_fd_sc_hd__nand3_1 _20204_ (.A(_10029_),
    .B(_10035_),
    .C(_10037_),
    .Y(_10040_));
 sky130_fd_sc_hd__o21ai_1 _20205_ (.A1(_10034_),
    .A2(_10036_),
    .B1(_10029_),
    .Y(_10041_));
 sky130_fd_sc_hd__nand3b_1 _20206_ (.A_N(_10029_),
    .B(_10035_),
    .C(_10037_),
    .Y(_10042_));
 sky130_fd_sc_hd__a31oi_1 _20207_ (.A1(_09893_),
    .A2(_09894_),
    .A3(_09895_),
    .B1(_09902_),
    .Y(_10043_));
 sky130_fd_sc_hd__a21oi_1 _20208_ (.A1(_09899_),
    .A2(_09903_),
    .B1(_09897_),
    .Y(_10044_));
 sky130_fd_sc_hd__nand3_2 _20209_ (.A(_10041_),
    .B(_10042_),
    .C(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__o211ai_2 _20210_ (.A1(_09897_),
    .A2(_10043_),
    .B1(_10040_),
    .C1(_10039_),
    .Y(_10046_));
 sky130_fd_sc_hd__a21o_1 _20211_ (.A1(_10045_),
    .A2(_10046_),
    .B1(_10028_),
    .X(_10047_));
 sky130_fd_sc_hd__nand3_1 _20212_ (.A(_10028_),
    .B(_10045_),
    .C(_10046_),
    .Y(_10048_));
 sky130_fd_sc_hd__nand4_1 _20213_ (.A(_09601_),
    .B(_09603_),
    .C(_10045_),
    .D(_10046_),
    .Y(_10050_));
 sky130_fd_sc_hd__a22o_1 _20214_ (.A1(_09601_),
    .A2(_09603_),
    .B1(_10045_),
    .B2(_10046_),
    .X(_10051_));
 sky130_fd_sc_hd__o21ai_1 _20215_ (.A1(_09906_),
    .A2(_09908_),
    .B1(_09891_),
    .Y(_10052_));
 sky130_fd_sc_hd__nand4_4 _20216_ (.A(_09889_),
    .B(_10047_),
    .C(_10048_),
    .D(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__nand4_4 _20217_ (.A(_09891_),
    .B(_09910_),
    .C(_10050_),
    .D(_10051_),
    .Y(_10054_));
 sky130_fd_sc_hd__o31a_1 _20218_ (.A1(_09602_),
    .A2(_09604_),
    .A3(_09607_),
    .B1(_09615_),
    .X(_10055_));
 sky130_fd_sc_hd__o2bb2ai_4 _20219_ (.A1_N(_10053_),
    .A2_N(_10054_),
    .B1(_10055_),
    .B2(_09608_),
    .Y(_10056_));
 sky130_fd_sc_hd__o211ai_4 _20220_ (.A1(_09611_),
    .A2(_09616_),
    .B1(_10053_),
    .C1(_10054_),
    .Y(_10057_));
 sky130_fd_sc_hd__a32o_1 _20221_ (.A1(_09618_),
    .A2(_09619_),
    .A3(_09624_),
    .B1(_09625_),
    .B2(_09629_),
    .X(_10058_));
 sky130_fd_sc_hd__a21oi_4 _20222_ (.A1(_10056_),
    .A2(_10057_),
    .B1(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__o211a_1 _20223_ (.A1(_09626_),
    .A2(_09633_),
    .B1(_10056_),
    .C1(_10057_),
    .X(_10061_));
 sky130_fd_sc_hd__o211ai_4 _20224_ (.A1(_09626_),
    .A2(_09633_),
    .B1(_10056_),
    .C1(_10057_),
    .Y(_10062_));
 sky130_fd_sc_hd__a32oi_4 _20225_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net28),
    .Y(_10063_));
 sky130_fd_sc_hd__a32o_1 _20226_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net28),
    .X(_10064_));
 sky130_fd_sc_hd__a21oi_1 _20227_ (.A1(_09653_),
    .A2(_09655_),
    .B1(_09650_),
    .Y(_10065_));
 sky130_fd_sc_hd__a21o_1 _20228_ (.A1(_09653_),
    .A2(_09655_),
    .B1(_09650_),
    .X(_10066_));
 sky130_fd_sc_hd__a32o_1 _20229_ (.A1(_06486_),
    .A2(net259),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net30),
    .X(_10067_));
 sky130_fd_sc_hd__or3_1 _20230_ (.A(net51),
    .B(_04190_),
    .C(_03949_),
    .X(_10068_));
 sky130_fd_sc_hd__o211ai_4 _20231_ (.A1(net259),
    .A2(_08656_),
    .B1(_06863_),
    .C1(_08700_),
    .Y(_10069_));
 sky130_fd_sc_hd__nor2_1 _20232_ (.A(_03938_),
    .B(_07226_),
    .Y(_10070_));
 sky130_fd_sc_hd__and3_1 _20233_ (.A(_07242_),
    .B(net257),
    .C(_07223_),
    .X(_10072_));
 sky130_fd_sc_hd__a31oi_2 _20234_ (.A1(_07242_),
    .A2(net257),
    .A3(_07223_),
    .B1(_10070_),
    .Y(_10073_));
 sky130_fd_sc_hd__a21oi_2 _20235_ (.A1(_10068_),
    .A2(_10069_),
    .B1(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__o2bb2ai_2 _20236_ (.A1_N(_10068_),
    .A2_N(_10069_),
    .B1(_10070_),
    .B2(_10072_),
    .Y(_10075_));
 sky130_fd_sc_hd__o211ai_2 _20237_ (.A1(_03949_),
    .A2(_06866_),
    .B1(_10069_),
    .C1(_10073_),
    .Y(_10076_));
 sky130_fd_sc_hd__a21oi_1 _20238_ (.A1(_10075_),
    .A2(_10076_),
    .B1(_10067_),
    .Y(_10077_));
 sky130_fd_sc_hd__a21o_1 _20239_ (.A1(_10075_),
    .A2(_10076_),
    .B1(_10067_),
    .X(_10078_));
 sky130_fd_sc_hd__nand2_1 _20240_ (.A(_10067_),
    .B(_10076_),
    .Y(_10079_));
 sky130_fd_sc_hd__and3_1 _20241_ (.A(_10067_),
    .B(_10075_),
    .C(_10076_),
    .X(_10080_));
 sky130_fd_sc_hd__o21a_1 _20242_ (.A1(_10077_),
    .A2(_10080_),
    .B1(_10065_),
    .X(_10081_));
 sky130_fd_sc_hd__o21ai_2 _20243_ (.A1(_10077_),
    .A2(_10080_),
    .B1(_10065_),
    .Y(_10083_));
 sky130_fd_sc_hd__o211ai_4 _20244_ (.A1(_10079_),
    .A2(_10074_),
    .B1(_10066_),
    .C1(_10078_),
    .Y(_10084_));
 sky130_fd_sc_hd__a22oi_4 _20245_ (.A1(_05874_),
    .A2(_07642_),
    .B1(_07643_),
    .B2(net29),
    .Y(_10085_));
 sky130_fd_sc_hd__a32o_1 _20246_ (.A1(_05841_),
    .A2(net265),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net29),
    .X(_10086_));
 sky130_fd_sc_hd__a21o_1 _20247_ (.A1(_10083_),
    .A2(_10084_),
    .B1(_10086_),
    .X(_10087_));
 sky130_fd_sc_hd__nand3_1 _20248_ (.A(_10083_),
    .B(_10084_),
    .C(_10086_),
    .Y(_10088_));
 sky130_fd_sc_hd__a21o_1 _20249_ (.A1(_10083_),
    .A2(_10084_),
    .B1(_10085_),
    .X(_10089_));
 sky130_fd_sc_hd__nand3_1 _20250_ (.A(_10083_),
    .B(_10084_),
    .C(_10085_),
    .Y(_10090_));
 sky130_fd_sc_hd__o21ai_1 _20251_ (.A1(_09642_),
    .A2(_09644_),
    .B1(_09660_),
    .Y(_10091_));
 sky130_fd_sc_hd__o31a_1 _20252_ (.A1(_09642_),
    .A2(_09644_),
    .A3(_09662_),
    .B1(_09660_),
    .X(_10092_));
 sky130_fd_sc_hd__and4_1 _20253_ (.A(_09663_),
    .B(_10089_),
    .C(_10090_),
    .D(_10091_),
    .X(_10094_));
 sky130_fd_sc_hd__o2111ai_2 _20254_ (.A1(_09645_),
    .A2(_09659_),
    .B1(_09663_),
    .C1(_10089_),
    .D1(_10090_),
    .Y(_10095_));
 sky130_fd_sc_hd__nand3_2 _20255_ (.A(_10087_),
    .B(_10088_),
    .C(_10092_),
    .Y(_10096_));
 sky130_fd_sc_hd__a21o_1 _20256_ (.A1(_10095_),
    .A2(_10096_),
    .B1(_10064_),
    .X(_10097_));
 sky130_fd_sc_hd__nand3_1 _20257_ (.A(_10064_),
    .B(_10095_),
    .C(_10096_),
    .Y(_10098_));
 sky130_fd_sc_hd__nand2_2 _20258_ (.A(_10097_),
    .B(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__nand3b_2 _20259_ (.A_N(_10059_),
    .B(_10062_),
    .C(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__o21bai_2 _20260_ (.A1(_10059_),
    .A2(_10061_),
    .B1_N(_10099_),
    .Y(_10101_));
 sky130_fd_sc_hd__o2111a_1 _20261_ (.A1(_09871_),
    .A2(_09963_),
    .B1(_10100_),
    .C1(_10101_),
    .D1(_09961_),
    .X(_10102_));
 sky130_fd_sc_hd__o2111ai_2 _20262_ (.A1(_09871_),
    .A2(_09963_),
    .B1(_10100_),
    .C1(_10101_),
    .D1(_09961_),
    .Y(_10103_));
 sky130_fd_sc_hd__a2bb2oi_2 _20263_ (.A1_N(_09960_),
    .A2_N(_09965_),
    .B1(_10100_),
    .B2(_10101_),
    .Y(_10105_));
 sky130_fd_sc_hd__a2bb2o_1 _20264_ (.A1_N(_09960_),
    .A2_N(_09965_),
    .B1(_10100_),
    .B2(_10101_),
    .X(_10106_));
 sky130_fd_sc_hd__o21ai_1 _20265_ (.A1(_09637_),
    .A2(_09675_),
    .B1(_09639_),
    .Y(_10107_));
 sky130_fd_sc_hd__o221a_1 _20266_ (.A1(_09637_),
    .A2(_09675_),
    .B1(_10102_),
    .B2(_10105_),
    .C1(_09639_),
    .X(_10108_));
 sky130_fd_sc_hd__o22ai_1 _20267_ (.A1(_09637_),
    .A2(_09679_),
    .B1(_10102_),
    .B2(_10105_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand2_1 _20268_ (.A(_10103_),
    .B(_10107_),
    .Y(_10110_));
 sky130_fd_sc_hd__and3_1 _20269_ (.A(_10103_),
    .B(_10106_),
    .C(_10107_),
    .X(_10111_));
 sky130_fd_sc_hd__o21a_1 _20270_ (.A1(_10102_),
    .A2(_10105_),
    .B1(_10107_),
    .X(_10112_));
 sky130_fd_sc_hd__o211a_1 _20271_ (.A1(_09637_),
    .A2(_09679_),
    .B1(_10103_),
    .C1(_10106_),
    .X(_10113_));
 sky130_fd_sc_hd__o21a_1 _20272_ (.A1(_10105_),
    .A2(_10110_),
    .B1(_10109_),
    .X(_10114_));
 sky130_fd_sc_hd__o21ai_1 _20273_ (.A1(_10105_),
    .A2(_10110_),
    .B1(_10109_),
    .Y(_10116_));
 sky130_fd_sc_hd__a32o_1 _20274_ (.A1(_09703_),
    .A2(_09862_),
    .A3(_09865_),
    .B1(_09966_),
    .B2(_09968_),
    .X(_10117_));
 sky130_fd_sc_hd__nand2_2 _20275_ (.A(_09867_),
    .B(_09969_),
    .Y(_10118_));
 sky130_fd_sc_hd__o22a_1 _20276_ (.A1(_09937_),
    .A2(_09933_),
    .B1(_09915_),
    .B2(_09935_),
    .X(_10119_));
 sky130_fd_sc_hd__a21o_1 _20277_ (.A1(_09928_),
    .A2(_09930_),
    .B1(_09924_),
    .X(_10120_));
 sky130_fd_sc_hd__a21oi_2 _20278_ (.A1(_09799_),
    .A2(_09802_),
    .B1(_09795_),
    .Y(_10121_));
 sky130_fd_sc_hd__o21a_1 _20279_ (.A1(_09799_),
    .A2(_09802_),
    .B1(_09795_),
    .X(_10122_));
 sky130_fd_sc_hd__o311a_1 _20280_ (.A1(net7),
    .A2(net248),
    .A3(_04787_),
    .B1(net281),
    .C1(net214),
    .X(_10123_));
 sky130_fd_sc_hd__nor2_1 _20281_ (.A(_04091_),
    .B(_04218_),
    .Y(_10124_));
 sky130_fd_sc_hd__a31o_1 _20282_ (.A1(net214),
    .A2(net281),
    .A3(net184),
    .B1(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__nand3_2 _20283_ (.A(net182),
    .B(net179),
    .C(_02858_),
    .Y(_10127_));
 sky130_fd_sc_hd__or3b_1 _20284_ (.A(net38),
    .B(_04135_),
    .C_N(net37),
    .X(_10128_));
 sky130_fd_sc_hd__nor2_1 _20285_ (.A(_04113_),
    .B(_03737_),
    .Y(_10129_));
 sky130_fd_sc_hd__o311a_1 _20286_ (.A1(net11),
    .A2(_04557_),
    .A3(net208),
    .B1(net285),
    .C1(net210),
    .X(_10130_));
 sky130_fd_sc_hd__a31oi_2 _20287_ (.A1(net210),
    .A2(net183),
    .A3(net285),
    .B1(_10129_),
    .Y(_10131_));
 sky130_fd_sc_hd__o211ai_4 _20288_ (.A1(_04135_),
    .A2(_02891_),
    .B1(_10127_),
    .C1(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__o2bb2a_2 _20289_ (.A1_N(_10127_),
    .A2_N(_10128_),
    .B1(_10129_),
    .B2(_10130_),
    .X(_10133_));
 sky130_fd_sc_hd__o2bb2ai_2 _20290_ (.A1_N(_10127_),
    .A2_N(_10128_),
    .B1(_10129_),
    .B2(_10130_),
    .Y(_10134_));
 sky130_fd_sc_hd__o211a_2 _20291_ (.A1(_10123_),
    .A2(_10124_),
    .B1(_10132_),
    .C1(_10134_),
    .X(_10135_));
 sky130_fd_sc_hd__o211ai_2 _20292_ (.A1(_10123_),
    .A2(_10124_),
    .B1(_10132_),
    .C1(_10134_),
    .Y(_10136_));
 sky130_fd_sc_hd__a21oi_2 _20293_ (.A1(_10132_),
    .A2(_10134_),
    .B1(_10125_),
    .Y(_10138_));
 sky130_fd_sc_hd__a21o_1 _20294_ (.A1(_10132_),
    .A2(_10134_),
    .B1(_10125_),
    .X(_10139_));
 sky130_fd_sc_hd__o211a_1 _20295_ (.A1(_09803_),
    .A2(_10122_),
    .B1(_10136_),
    .C1(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__o211ai_2 _20296_ (.A1(_09803_),
    .A2(_10122_),
    .B1(_10136_),
    .C1(_10139_),
    .Y(_10141_));
 sky130_fd_sc_hd__o22ai_4 _20297_ (.A1(_09805_),
    .A2(_10121_),
    .B1(_10135_),
    .B2(_10138_),
    .Y(_10142_));
 sky130_fd_sc_hd__a21o_1 _20298_ (.A1(_10141_),
    .A2(_10142_),
    .B1(_10120_),
    .X(_10143_));
 sky130_fd_sc_hd__o21ai_4 _20299_ (.A1(_09924_),
    .A2(_09933_),
    .B1(_10142_),
    .Y(_10144_));
 sky130_fd_sc_hd__nand4_1 _20300_ (.A(_09925_),
    .B(_09934_),
    .C(_10141_),
    .D(_10142_),
    .Y(_10145_));
 sky130_fd_sc_hd__a22o_1 _20301_ (.A1(_09925_),
    .A2(_09934_),
    .B1(_10141_),
    .B2(_10142_),
    .X(_10146_));
 sky130_fd_sc_hd__nand3_2 _20302_ (.A(_10146_),
    .B(_10119_),
    .C(_10145_),
    .Y(_10147_));
 sky130_fd_sc_hd__o221ai_4 _20303_ (.A1(_10140_),
    .A2(_10144_),
    .B1(_09938_),
    .B2(_09944_),
    .C1(_10143_),
    .Y(_10149_));
 sky130_fd_sc_hd__nand2_1 _20304_ (.A(_10147_),
    .B(_10149_),
    .Y(_10150_));
 sky130_fd_sc_hd__a32o_1 _20305_ (.A1(_00625_),
    .A2(net250),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net5),
    .X(_10151_));
 sky130_fd_sc_hd__nand2_1 _20306_ (.A(net248),
    .B(net276),
    .Y(_10152_));
 sky130_fd_sc_hd__o32a_1 _20307_ (.A1(_04026_),
    .A2(_04124_),
    .A3(net46),
    .B1(_02410_),
    .B2(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__o22ai_1 _20308_ (.A1(_04026_),
    .A2(_05229_),
    .B1(_02410_),
    .B2(_10152_),
    .Y(_10154_));
 sky130_fd_sc_hd__a311o_1 _20309_ (.A1(_06519_),
    .A2(net286),
    .A3(net283),
    .B1(_04986_),
    .C1(_03951_),
    .X(_10155_));
 sky130_fd_sc_hd__or3_1 _20310_ (.A(net45),
    .B(_04102_),
    .C(_04048_),
    .X(_10156_));
 sky130_fd_sc_hd__o32a_1 _20311_ (.A1(_04986_),
    .A2(_03957_),
    .A3(_03951_),
    .B1(_04048_),
    .B2(_04989_),
    .X(_10157_));
 sky130_fd_sc_hd__o31ai_1 _20312_ (.A1(_04986_),
    .A2(_03957_),
    .A3(_03951_),
    .B1(_10156_),
    .Y(_10158_));
 sky130_fd_sc_hd__a21oi_1 _20313_ (.A1(_10155_),
    .A2(_10156_),
    .B1(_10153_),
    .Y(_10160_));
 sky130_fd_sc_hd__a21o_1 _20314_ (.A1(_10155_),
    .A2(_10156_),
    .B1(_10153_),
    .X(_10161_));
 sky130_fd_sc_hd__o311a_1 _20315_ (.A1(_04048_),
    .A2(_04102_),
    .A3(net45),
    .B1(_10153_),
    .C1(_10155_),
    .X(_10162_));
 sky130_fd_sc_hd__a221o_1 _20316_ (.A1(_03959_),
    .A2(net242),
    .B1(_04988_),
    .B2(net7),
    .C1(_10154_),
    .X(_10163_));
 sky130_fd_sc_hd__o21bai_2 _20317_ (.A1(_10160_),
    .A2(_10162_),
    .B1_N(_10151_),
    .Y(_10164_));
 sky130_fd_sc_hd__nand3_2 _20318_ (.A(_10151_),
    .B(_10161_),
    .C(_10163_),
    .Y(_10165_));
 sky130_fd_sc_hd__nand2_1 _20319_ (.A(_10164_),
    .B(_10165_),
    .Y(_10166_));
 sky130_fd_sc_hd__o21ai_1 _20320_ (.A1(_09875_),
    .A2(_09882_),
    .B1(_09881_),
    .Y(_10167_));
 sky130_fd_sc_hd__o21a_1 _20321_ (.A1(_09875_),
    .A2(_09882_),
    .B1(_09881_),
    .X(_10168_));
 sky130_fd_sc_hd__o22a_1 _20322_ (.A1(_04133_),
    .A2(_04896_),
    .B1(_04898_),
    .B2(_04059_),
    .X(_10169_));
 sky130_fd_sc_hd__a32o_1 _20323_ (.A1(net229),
    .A2(net228),
    .A3(net243),
    .B1(_04897_),
    .B2(net8),
    .X(_10171_));
 sky130_fd_sc_hd__nor2_1 _20324_ (.A(_04069_),
    .B(_04483_),
    .Y(_10172_));
 sky130_fd_sc_hd__o311a_1 _20325_ (.A1(net7),
    .A2(net248),
    .A3(_04407_),
    .B1(net279),
    .C1(net222),
    .X(_10173_));
 sky130_fd_sc_hd__a31oi_2 _20326_ (.A1(net188),
    .A2(net222),
    .A3(net279),
    .B1(_10172_),
    .Y(_10174_));
 sky130_fd_sc_hd__nor2_1 _20327_ (.A(_04080_),
    .B(_04270_),
    .Y(_10175_));
 sky130_fd_sc_hd__a31o_1 _20328_ (.A1(net218),
    .A2(net186),
    .A3(net280),
    .B1(_10175_),
    .X(_10176_));
 sky130_fd_sc_hd__o221a_2 _20329_ (.A1(_04080_),
    .A2(_04270_),
    .B1(_04562_),
    .B2(_04268_),
    .C1(_10174_),
    .X(_10177_));
 sky130_fd_sc_hd__o221ai_4 _20330_ (.A1(_04080_),
    .A2(_04270_),
    .B1(_04562_),
    .B2(_04268_),
    .C1(_10174_),
    .Y(_10178_));
 sky130_fd_sc_hd__o21ai_4 _20331_ (.A1(_10172_),
    .A2(_10173_),
    .B1(_10176_),
    .Y(_10179_));
 sky130_fd_sc_hd__o221a_1 _20332_ (.A1(_04133_),
    .A2(_04896_),
    .B1(_04898_),
    .B2(_04059_),
    .C1(_10179_),
    .X(_10180_));
 sky130_fd_sc_hd__o21ai_2 _20333_ (.A1(_10169_),
    .A2(_10177_),
    .B1(_10179_),
    .Y(_10182_));
 sky130_fd_sc_hd__a21o_1 _20334_ (.A1(_10178_),
    .A2(_10179_),
    .B1(_10169_),
    .X(_10183_));
 sky130_fd_sc_hd__nand3_2 _20335_ (.A(_10178_),
    .B(_10179_),
    .C(_10169_),
    .Y(_10184_));
 sky130_fd_sc_hd__a21o_1 _20336_ (.A1(_10178_),
    .A2(_10179_),
    .B1(_10171_),
    .X(_10185_));
 sky130_fd_sc_hd__nand3_1 _20337_ (.A(_10171_),
    .B(_10178_),
    .C(_10179_),
    .Y(_10186_));
 sky130_fd_sc_hd__a21o_2 _20338_ (.A1(_10185_),
    .A2(_10186_),
    .B1(_10167_),
    .X(_10187_));
 sky130_fd_sc_hd__a21oi_2 _20339_ (.A1(_10183_),
    .A2(_10184_),
    .B1(_10168_),
    .Y(_10188_));
 sky130_fd_sc_hd__nand3_1 _20340_ (.A(_10185_),
    .B(_10186_),
    .C(_10167_),
    .Y(_10189_));
 sky130_fd_sc_hd__nor2_1 _20341_ (.A(_10166_),
    .B(_10188_),
    .Y(_10190_));
 sky130_fd_sc_hd__and4_1 _20342_ (.A(_10164_),
    .B(_10165_),
    .C(_10187_),
    .D(_10189_),
    .X(_10191_));
 sky130_fd_sc_hd__a22oi_2 _20343_ (.A1(_10164_),
    .A2(_10165_),
    .B1(_10187_),
    .B2(_10189_),
    .Y(_10193_));
 sky130_fd_sc_hd__a21oi_1 _20344_ (.A1(_10187_),
    .A2(_10190_),
    .B1(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__inv_2 _20345_ (.A(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__o2bb2ai_2 _20346_ (.A1_N(_10147_),
    .A2_N(_10149_),
    .B1(_10191_),
    .B2(_10193_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand3_2 _20347_ (.A(_10147_),
    .B(_10149_),
    .C(_10194_),
    .Y(_10197_));
 sky130_fd_sc_hd__o21ai_1 _20348_ (.A1(_09406_),
    .A2(_09849_),
    .B1(_09853_),
    .Y(_10198_));
 sky130_fd_sc_hd__a21oi_2 _20349_ (.A1(_10196_),
    .A2(_10197_),
    .B1(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__o211a_1 _20350_ (.A1(_09851_),
    .A2(_09856_),
    .B1(_10196_),
    .C1(_10197_),
    .X(_10200_));
 sky130_fd_sc_hd__o211ai_4 _20351_ (.A1(_09851_),
    .A2(_09856_),
    .B1(_10196_),
    .C1(_10197_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand3b_4 _20352_ (.A_N(_10199_),
    .B(_10201_),
    .C(_09958_),
    .Y(_10202_));
 sky130_fd_sc_hd__o22ai_4 _20353_ (.A1(_09948_),
    .A2(_09957_),
    .B1(_10199_),
    .B2(_10200_),
    .Y(_10204_));
 sky130_fd_sc_hd__nand2_1 _20354_ (.A(_10202_),
    .B(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__a32oi_4 _20355_ (.A1(_09704_),
    .A2(_09783_),
    .A3(_09785_),
    .B1(_09855_),
    .B2(_09858_),
    .Y(_10206_));
 sky130_fd_sc_hd__o22ai_4 _20356_ (.A1(_09784_),
    .A2(_09789_),
    .B1(_09792_),
    .B2(_09859_),
    .Y(_10207_));
 sky130_fd_sc_hd__o22a_1 _20357_ (.A1(_09784_),
    .A2(_09789_),
    .B1(_09792_),
    .B2(_09859_),
    .X(_10208_));
 sky130_fd_sc_hd__a311oi_4 _20358_ (.A1(_09284_),
    .A2(_09721_),
    .A3(_09723_),
    .B1(_09330_),
    .C1(_09335_),
    .Y(_10209_));
 sky130_fd_sc_hd__o21ai_1 _20359_ (.A1(_09330_),
    .A2(_09335_),
    .B1(_09725_),
    .Y(_10210_));
 sky130_fd_sc_hd__o21ai_1 _20360_ (.A1(_09719_),
    .A2(_09726_),
    .B1(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__o2111ai_4 _20361_ (.A1(_05927_),
    .A2(_06220_),
    .B1(net35),
    .C1(net201),
    .D1(_03971_),
    .Y(_10212_));
 sky130_fd_sc_hd__or3_2 _20362_ (.A(net35),
    .B(_04168_),
    .C(_03971_),
    .X(_10213_));
 sky130_fd_sc_hd__o211ai_4 _20363_ (.A1(net231),
    .A2(_05927_),
    .B1(_12330_),
    .C1(_05933_),
    .Y(_10215_));
 sky130_fd_sc_hd__or3_1 _20364_ (.A(net36),
    .B(_04157_),
    .C(_03993_),
    .X(_10216_));
 sky130_fd_sc_hd__a22oi_4 _20365_ (.A1(_10212_),
    .A2(_10213_),
    .B1(_10215_),
    .B2(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__a22o_1 _20366_ (.A1(_10212_),
    .A2(_10213_),
    .B1(_10215_),
    .B2(_10216_),
    .X(_10218_));
 sky130_fd_sc_hd__o2111ai_4 _20367_ (.A1(_04157_),
    .A2(_12363_),
    .B1(_10212_),
    .C1(_10213_),
    .D1(_10215_),
    .Y(_10219_));
 sky130_fd_sc_hd__o32a_1 _20368_ (.A1(_01304_),
    .A2(_05548_),
    .A3(net206),
    .B1(_01326_),
    .B2(_04146_),
    .X(_10220_));
 sky130_fd_sc_hd__a32o_1 _20369_ (.A1(net178),
    .A2(net177),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net15),
    .X(_10221_));
 sky130_fd_sc_hd__a21oi_2 _20370_ (.A1(_10218_),
    .A2(_10219_),
    .B1(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__nor2_1 _20371_ (.A(_10217_),
    .B(_10220_),
    .Y(_10223_));
 sky130_fd_sc_hd__and3_2 _20372_ (.A(_10218_),
    .B(_10219_),
    .C(_10221_),
    .X(_10224_));
 sky130_fd_sc_hd__a21oi_2 _20373_ (.A1(_10219_),
    .A2(_10223_),
    .B1(_10222_),
    .Y(_10226_));
 sky130_fd_sc_hd__and3_1 _20374_ (.A(_03971_),
    .B(net18),
    .C(net64),
    .X(_10227_));
 sky130_fd_sc_hd__o311a_1 _20375_ (.A1(net246),
    .A2(_05928_),
    .A3(_06451_),
    .B1(net289),
    .C1(net199),
    .X(_10228_));
 sky130_fd_sc_hd__o22a_1 _20376_ (.A1(_04179_),
    .A2(_10346_),
    .B1(_06454_),
    .B2(_10324_),
    .X(_10229_));
 sky130_fd_sc_hd__a31o_1 _20377_ (.A1(net199),
    .A2(net172),
    .A3(net289),
    .B1(_10227_),
    .X(_10230_));
 sky130_fd_sc_hd__nand3_2 _20378_ (.A(net195),
    .B(net171),
    .C(net291),
    .Y(_10231_));
 sky130_fd_sc_hd__or3b_1 _20379_ (.A(net64),
    .B(_04201_),
    .C_N(net63),
    .X(_10232_));
 sky130_fd_sc_hd__a32oi_4 _20380_ (.A1(net195),
    .A2(net171),
    .A3(net291),
    .B1(_08272_),
    .B2(net19),
    .Y(_10233_));
 sky130_fd_sc_hd__nor2_2 _20381_ (.A(_04212_),
    .B(_07691_),
    .Y(_10234_));
 sky130_fd_sc_hd__a221oi_2 _20382_ (.A1(net203),
    .A2(_07073_),
    .B1(net171),
    .B2(net20),
    .C1(_07669_),
    .Y(_10235_));
 sky130_fd_sc_hd__o211ai_2 _20383_ (.A1(net175),
    .A2(_07074_),
    .B1(_07658_),
    .C1(_07072_),
    .Y(_10237_));
 sky130_fd_sc_hd__o211ai_4 _20384_ (.A1(_04201_),
    .A2(_08283_),
    .B1(_10231_),
    .C1(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__o221ai_4 _20385_ (.A1(_04212_),
    .A2(_07691_),
    .B1(_07079_),
    .B2(_07669_),
    .C1(_10233_),
    .Y(_10239_));
 sky130_fd_sc_hd__o2bb2ai_4 _20386_ (.A1_N(_10231_),
    .A2_N(_10232_),
    .B1(_10234_),
    .B2(_10235_),
    .Y(_10240_));
 sky130_fd_sc_hd__o21ai_2 _20387_ (.A1(_10234_),
    .A2(_10238_),
    .B1(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__o221a_4 _20388_ (.A1(_10227_),
    .A2(_10228_),
    .B1(_10234_),
    .B2(_10238_),
    .C1(_10240_),
    .X(_10242_));
 sky130_fd_sc_hd__o221ai_4 _20389_ (.A1(_10227_),
    .A2(_10228_),
    .B1(_10234_),
    .B2(_10238_),
    .C1(_10240_),
    .Y(_10243_));
 sky130_fd_sc_hd__a21oi_2 _20390_ (.A1(_10239_),
    .A2(_10240_),
    .B1(_10230_),
    .Y(_10244_));
 sky130_fd_sc_hd__a21o_1 _20391_ (.A1(_10239_),
    .A2(_10240_),
    .B1(_10230_),
    .X(_10245_));
 sky130_fd_sc_hd__o2bb2ai_2 _20392_ (.A1_N(_10229_),
    .A2_N(_10241_),
    .B1(_09827_),
    .B2(_09832_),
    .Y(_10246_));
 sky130_fd_sc_hd__o211ai_1 _20393_ (.A1(_09827_),
    .A2(_09832_),
    .B1(_10243_),
    .C1(_10245_),
    .Y(_10248_));
 sky130_fd_sc_hd__o221a_1 _20394_ (.A1(_09814_),
    .A2(_09826_),
    .B1(_10242_),
    .B2(_10244_),
    .C1(_09828_),
    .X(_10249_));
 sky130_fd_sc_hd__o22ai_4 _20395_ (.A1(_09826_),
    .A2(_09831_),
    .B1(_10242_),
    .B2(_10244_),
    .Y(_10250_));
 sky130_fd_sc_hd__o21ai_1 _20396_ (.A1(_10242_),
    .A2(_10246_),
    .B1(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__o211a_1 _20397_ (.A1(_10242_),
    .A2(_10246_),
    .B1(_10226_),
    .C1(_10250_),
    .X(_10252_));
 sky130_fd_sc_hd__o211ai_4 _20398_ (.A1(_10242_),
    .A2(_10246_),
    .B1(_10226_),
    .C1(_10250_),
    .Y(_10253_));
 sky130_fd_sc_hd__a21oi_2 _20399_ (.A1(_10248_),
    .A2(_10250_),
    .B1(_10226_),
    .Y(_10254_));
 sky130_fd_sc_hd__o21ai_2 _20400_ (.A1(_10222_),
    .A2(_10224_),
    .B1(_10251_),
    .Y(_10255_));
 sky130_fd_sc_hd__a21oi_2 _20401_ (.A1(_09727_),
    .A2(_10210_),
    .B1(_10254_),
    .Y(_10256_));
 sky130_fd_sc_hd__nand3_2 _20402_ (.A(_10211_),
    .B(_10253_),
    .C(_10255_),
    .Y(_10257_));
 sky130_fd_sc_hd__a2bb2oi_2 _20403_ (.A1_N(_09724_),
    .A2_N(_10209_),
    .B1(_10253_),
    .B2(_10255_),
    .Y(_10259_));
 sky130_fd_sc_hd__o22ai_4 _20404_ (.A1(_09724_),
    .A2(_10209_),
    .B1(_10252_),
    .B2(_10254_),
    .Y(_10260_));
 sky130_fd_sc_hd__o31a_1 _20405_ (.A1(_09807_),
    .A2(_09809_),
    .A3(_09839_),
    .B1(_09838_),
    .X(_10261_));
 sky130_fd_sc_hd__a21o_2 _20406_ (.A1(_09811_),
    .A2(_09840_),
    .B1(_09837_),
    .X(_10262_));
 sky130_fd_sc_hd__a21oi_2 _20407_ (.A1(_10257_),
    .A2(_10260_),
    .B1(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__a21o_2 _20408_ (.A1(_10257_),
    .A2(_10260_),
    .B1(_10262_),
    .X(_10264_));
 sky130_fd_sc_hd__a31o_1 _20409_ (.A1(_10211_),
    .A2(_10253_),
    .A3(_10255_),
    .B1(_10261_),
    .X(_10265_));
 sky130_fd_sc_hd__and3_2 _20410_ (.A(_10257_),
    .B(_10260_),
    .C(_10262_),
    .X(_10266_));
 sky130_fd_sc_hd__nand3_2 _20411_ (.A(_10257_),
    .B(_10260_),
    .C(_10262_),
    .Y(_10267_));
 sky130_fd_sc_hd__o211ai_4 _20412_ (.A1(_09741_),
    .A2(_09747_),
    .B1(_09767_),
    .C1(_09768_),
    .Y(_10268_));
 sky130_fd_sc_hd__a31oi_1 _20413_ (.A1(_09743_),
    .A2(_09744_),
    .A3(_09745_),
    .B1(_09769_),
    .Y(_10270_));
 sky130_fd_sc_hd__a31o_1 _20414_ (.A1(_09746_),
    .A2(_09770_),
    .A3(_09771_),
    .B1(_09748_),
    .X(_10271_));
 sky130_fd_sc_hd__a21oi_2 _20415_ (.A1(_10270_),
    .A2(_09771_),
    .B1(_09748_),
    .Y(_10272_));
 sky130_fd_sc_hd__a32o_2 _20416_ (.A1(_04998_),
    .A2(net300),
    .A3(_08657_),
    .B1(_08659_),
    .B2(net27),
    .X(_10273_));
 sky130_fd_sc_hd__a31oi_4 _20417_ (.A1(net162),
    .A2(net33),
    .A3(net319),
    .B1(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__a31o_1 _20418_ (.A1(net162),
    .A2(net33),
    .A3(net319),
    .B1(_10273_),
    .X(_10275_));
 sky130_fd_sc_hd__and3_1 _20419_ (.A(_10273_),
    .B(net33),
    .C(net319),
    .X(_10276_));
 sky130_fd_sc_hd__nand3_1 _20420_ (.A(_10273_),
    .B(net33),
    .C(net319),
    .Y(_10277_));
 sky130_fd_sc_hd__o21ai_2 _20421_ (.A1(_10274_),
    .A2(_10276_),
    .B1(net148),
    .Y(_10278_));
 sky130_fd_sc_hd__o22ai_1 _20422_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_10274_),
    .B2(_10276_),
    .Y(_10279_));
 sky130_fd_sc_hd__nand3_1 _20423_ (.A(_10275_),
    .B(_10277_),
    .C(net148),
    .Y(_10281_));
 sky130_fd_sc_hd__o21ai_1 _20424_ (.A1(net147),
    .A2(_10274_),
    .B1(_10278_),
    .Y(_10282_));
 sky130_fd_sc_hd__o211ai_1 _20425_ (.A1(net319),
    .A2(_04331_),
    .B1(_09298_),
    .C1(_09739_),
    .Y(_10283_));
 sky130_fd_sc_hd__o21ai_1 _20426_ (.A1(net148),
    .A2(_09737_),
    .B1(_09739_),
    .Y(_10284_));
 sky130_fd_sc_hd__o21ai_2 _20427_ (.A1(_09736_),
    .A2(_08877_),
    .B1(_10283_),
    .Y(_10285_));
 sky130_fd_sc_hd__nand3_2 _20428_ (.A(_10279_),
    .B(_10281_),
    .C(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__o221a_1 _20429_ (.A1(_09738_),
    .A2(_09741_),
    .B1(_10274_),
    .B2(net148),
    .C1(_10278_),
    .X(_10287_));
 sky130_fd_sc_hd__o211ai_4 _20430_ (.A1(net148),
    .A2(_10274_),
    .B1(_10284_),
    .C1(_10278_),
    .Y(_10288_));
 sky130_fd_sc_hd__a21oi_2 _20431_ (.A1(net151),
    .A2(net158),
    .B1(_04900_),
    .Y(_10289_));
 sky130_fd_sc_hd__and3b_2 _20432_ (.A_N(net59),
    .B(net25),
    .C(net58),
    .X(_10290_));
 sky130_fd_sc_hd__or3b_2 _20433_ (.A(net59),
    .B(net319),
    .C_N(net58),
    .X(_10292_));
 sky130_fd_sc_hd__a22oi_4 _20434_ (.A1(net25),
    .A2(_04911_),
    .B1(_08670_),
    .B2(_04889_),
    .Y(_10293_));
 sky130_fd_sc_hd__o211ai_1 _20435_ (.A1(net169),
    .A2(net268),
    .B1(net319),
    .C1(_04627_),
    .Y(_10294_));
 sky130_fd_sc_hd__a31oi_4 _20436_ (.A1(net319),
    .A2(net163),
    .A3(_04627_),
    .B1(_09758_),
    .Y(_10295_));
 sky130_fd_sc_hd__a31o_4 _20437_ (.A1(_04277_),
    .A2(net163),
    .A3(_04627_),
    .B1(_09758_),
    .X(_10296_));
 sky130_fd_sc_hd__o311a_4 _20438_ (.A1(net25),
    .A2(_04638_),
    .A3(_08207_),
    .B1(_09759_),
    .C1(_09754_),
    .X(_10297_));
 sky130_fd_sc_hd__o211a_1 _20439_ (.A1(_04900_),
    .A2(_08669_),
    .B1(_10292_),
    .C1(_10297_),
    .X(_10298_));
 sky130_fd_sc_hd__nand2_1 _20440_ (.A(_10293_),
    .B(_10297_),
    .Y(_10299_));
 sky130_fd_sc_hd__o22a_2 _20441_ (.A1(_09755_),
    .A2(_10296_),
    .B1(_10290_),
    .B2(_10289_),
    .X(_10300_));
 sky130_fd_sc_hd__o22ai_4 _20442_ (.A1(_09755_),
    .A2(_10296_),
    .B1(_10290_),
    .B2(_10289_),
    .Y(_10301_));
 sky130_fd_sc_hd__a22oi_2 _20443_ (.A1(_10286_),
    .A2(_10288_),
    .B1(_10299_),
    .B2(_10301_),
    .Y(_10303_));
 sky130_fd_sc_hd__o2bb2ai_2 _20444_ (.A1_N(_10286_),
    .A2_N(_10288_),
    .B1(_10298_),
    .B2(_10300_),
    .Y(_10304_));
 sky130_fd_sc_hd__nand3_4 _20445_ (.A(_10286_),
    .B(_10299_),
    .C(_10301_),
    .Y(_10305_));
 sky130_fd_sc_hd__and4_1 _20446_ (.A(_10286_),
    .B(_10288_),
    .C(_10299_),
    .D(_10301_),
    .X(_10306_));
 sky130_fd_sc_hd__o21ai_2 _20447_ (.A1(_10287_),
    .A2(_10305_),
    .B1(_10304_),
    .Y(_10307_));
 sky130_fd_sc_hd__inv_2 _20448_ (.A(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__o2111ai_4 _20449_ (.A1(_10287_),
    .A2(_10305_),
    .B1(_10304_),
    .C1(_09746_),
    .D1(_10268_),
    .Y(_10309_));
 sky130_fd_sc_hd__o2bb2ai_4 _20450_ (.A1_N(_09746_),
    .A2_N(_10268_),
    .B1(_10303_),
    .B2(_10306_),
    .Y(_10310_));
 sky130_fd_sc_hd__a21oi_2 _20451_ (.A1(_09707_),
    .A2(_09718_),
    .B1(_09716_),
    .Y(_10311_));
 sky130_fd_sc_hd__a21o_1 _20452_ (.A1(_09707_),
    .A2(_09718_),
    .B1(_09716_),
    .X(_10312_));
 sky130_fd_sc_hd__nand2_1 _20453_ (.A(_09766_),
    .B(_09770_),
    .Y(_10314_));
 sky130_fd_sc_hd__o21a_1 _20454_ (.A1(_09761_),
    .A2(_09762_),
    .B1(_09766_),
    .X(_10315_));
 sky130_fd_sc_hd__o211ai_2 _20455_ (.A1(net168),
    .A2(_07765_),
    .B1(_05688_),
    .C1(_07771_),
    .Y(_10316_));
 sky130_fd_sc_hd__nor2_1 _20456_ (.A(_04245_),
    .B(_05720_),
    .Y(_10317_));
 sky130_fd_sc_hd__or3b_1 _20457_ (.A(net61),
    .B(_04245_),
    .C_N(net60),
    .X(_10318_));
 sky130_fd_sc_hd__a31oi_4 _20458_ (.A1(_07771_),
    .A2(_05688_),
    .A3(_07769_),
    .B1(_10317_),
    .Y(_10319_));
 sky130_fd_sc_hd__o211ai_2 _20459_ (.A1(net168),
    .A2(_08206_),
    .B1(_05227_),
    .C1(_08204_),
    .Y(_10320_));
 sky130_fd_sc_hd__or3b_2 _20460_ (.A(net60),
    .B(_04256_),
    .C_N(net59),
    .X(_10321_));
 sky130_fd_sc_hd__a22oi_4 _20461_ (.A1(_10316_),
    .A2(_10318_),
    .B1(_10320_),
    .B2(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__o311a_4 _20462_ (.A1(_05238_),
    .A2(_08203_),
    .A3(net154),
    .B1(_10321_),
    .C1(_10319_),
    .X(_10323_));
 sky130_fd_sc_hd__o221ai_4 _20463_ (.A1(_04256_),
    .A2(_05260_),
    .B1(_08209_),
    .B2(_05238_),
    .C1(_10319_),
    .Y(_10325_));
 sky130_fd_sc_hd__o32a_2 _20464_ (.A1(_06837_),
    .A2(_07498_),
    .A3(_07502_),
    .B1(_06859_),
    .B2(_04223_),
    .X(_10326_));
 sky130_fd_sc_hd__a32o_2 _20465_ (.A1(_07499_),
    .A2(net167),
    .A3(_06826_),
    .B1(_06848_),
    .B2(net21),
    .X(_10327_));
 sky130_fd_sc_hd__nor3_1 _20466_ (.A(_10322_),
    .B(_10327_),
    .C(_10323_),
    .Y(_10328_));
 sky130_fd_sc_hd__nand3b_4 _20467_ (.A_N(_10322_),
    .B(_10325_),
    .C(_10326_),
    .Y(_10329_));
 sky130_fd_sc_hd__o21a_1 _20468_ (.A1(_10322_),
    .A2(_10323_),
    .B1(_10327_),
    .X(_10330_));
 sky130_fd_sc_hd__o21ai_4 _20469_ (.A1(_10322_),
    .A2(_10323_),
    .B1(_10327_),
    .Y(_10331_));
 sky130_fd_sc_hd__o21ai_2 _20470_ (.A1(_10322_),
    .A2(_10323_),
    .B1(_10326_),
    .Y(_10332_));
 sky130_fd_sc_hd__nand3b_1 _20471_ (.A_N(_10322_),
    .B(_10325_),
    .C(_10327_),
    .Y(_10333_));
 sky130_fd_sc_hd__o2111ai_4 _20472_ (.A1(_09761_),
    .A2(_09762_),
    .B1(_09766_),
    .C1(_10329_),
    .D1(_10331_),
    .Y(_10334_));
 sky130_fd_sc_hd__a2bb2oi_1 _20473_ (.A1_N(_09765_),
    .A2_N(_09769_),
    .B1(_10329_),
    .B2(_10331_),
    .Y(_10336_));
 sky130_fd_sc_hd__o211ai_4 _20474_ (.A1(_09765_),
    .A2(_09769_),
    .B1(_10332_),
    .C1(_10333_),
    .Y(_10337_));
 sky130_fd_sc_hd__o211a_1 _20475_ (.A1(_09716_),
    .A2(_09722_),
    .B1(_10334_),
    .C1(_10337_),
    .X(_10338_));
 sky130_fd_sc_hd__o211ai_2 _20476_ (.A1(_09716_),
    .A2(_09722_),
    .B1(_10334_),
    .C1(_10337_),
    .Y(_10339_));
 sky130_fd_sc_hd__a21oi_1 _20477_ (.A1(_10334_),
    .A2(_10337_),
    .B1(_10312_),
    .Y(_10340_));
 sky130_fd_sc_hd__a21o_1 _20478_ (.A1(_10334_),
    .A2(_10337_),
    .B1(_10312_),
    .X(_10341_));
 sky130_fd_sc_hd__and3_1 _20479_ (.A(_10334_),
    .B(_10337_),
    .C(_10311_),
    .X(_10342_));
 sky130_fd_sc_hd__nand4_2 _20480_ (.A(_09717_),
    .B(_09723_),
    .C(_10334_),
    .D(_10337_),
    .Y(_10343_));
 sky130_fd_sc_hd__a21oi_1 _20481_ (.A1(_10334_),
    .A2(_10337_),
    .B1(_10311_),
    .Y(_10344_));
 sky130_fd_sc_hd__a22o_1 _20482_ (.A1(_09717_),
    .A2(_09723_),
    .B1(_10334_),
    .B2(_10337_),
    .X(_10345_));
 sky130_fd_sc_hd__nand4_2 _20483_ (.A(_10309_),
    .B(_10310_),
    .C(_10343_),
    .D(_10345_),
    .Y(_10347_));
 sky130_fd_sc_hd__o2bb2ai_2 _20484_ (.A1_N(_10309_),
    .A2_N(_10310_),
    .B1(_10342_),
    .B2(_10344_),
    .Y(_10348_));
 sky130_fd_sc_hd__o2bb2ai_1 _20485_ (.A1_N(_10309_),
    .A2_N(_10310_),
    .B1(_10338_),
    .B2(_10340_),
    .Y(_10349_));
 sky130_fd_sc_hd__nand4_2 _20486_ (.A(_10309_),
    .B(_10310_),
    .C(_10339_),
    .D(_10341_),
    .Y(_10350_));
 sky130_fd_sc_hd__nand2_2 _20487_ (.A(_10347_),
    .B(_10348_),
    .Y(_10351_));
 sky130_fd_sc_hd__o21ai_2 _20488_ (.A1(_09729_),
    .A2(_09732_),
    .B1(_09782_),
    .Y(_10352_));
 sky130_fd_sc_hd__a31o_2 _20489_ (.A1(_09730_),
    .A2(_09733_),
    .A3(_09780_),
    .B1(_09781_),
    .X(_10353_));
 sky130_fd_sc_hd__o2111ai_4 _20490_ (.A1(_09779_),
    .A2(_09735_),
    .B1(_10347_),
    .C1(_09782_),
    .D1(_10348_),
    .Y(_10354_));
 sky130_fd_sc_hd__inv_2 _20491_ (.A(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__nand4_4 _20492_ (.A(_09780_),
    .B(_10349_),
    .C(_10350_),
    .D(_10352_),
    .Y(_10356_));
 sky130_fd_sc_hd__nand2_1 _20493_ (.A(_10354_),
    .B(_10356_),
    .Y(_10358_));
 sky130_fd_sc_hd__nand4_4 _20494_ (.A(_10264_),
    .B(_10267_),
    .C(_10354_),
    .D(_10356_),
    .Y(_10359_));
 sky130_fd_sc_hd__a22o_2 _20495_ (.A1(_10264_),
    .A2(_10267_),
    .B1(_10354_),
    .B2(_10356_),
    .X(_10360_));
 sky130_fd_sc_hd__o211ai_4 _20496_ (.A1(_10263_),
    .A2(_10266_),
    .B1(_10354_),
    .C1(_10356_),
    .Y(_10361_));
 sky130_fd_sc_hd__o211ai_4 _20497_ (.A1(_10265_),
    .A2(_10259_),
    .B1(_10264_),
    .C1(_10358_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand3_2 _20498_ (.A(_10207_),
    .B(_10359_),
    .C(_10360_),
    .Y(_10363_));
 sky130_fd_sc_hd__and3_1 _20499_ (.A(_10208_),
    .B(_10361_),
    .C(_10362_),
    .X(_10364_));
 sky130_fd_sc_hd__o211ai_4 _20500_ (.A1(_09792_),
    .A2(_10206_),
    .B1(_10361_),
    .C1(_10362_),
    .Y(_10365_));
 sky130_fd_sc_hd__a21o_2 _20501_ (.A1(_10363_),
    .A2(_10365_),
    .B1(_10205_),
    .X(_10366_));
 sky130_fd_sc_hd__nand3_4 _20502_ (.A(_10205_),
    .B(_10363_),
    .C(_10365_),
    .Y(_10367_));
 sky130_fd_sc_hd__nand4_2 _20503_ (.A(_10202_),
    .B(_10204_),
    .C(_10363_),
    .D(_10365_),
    .Y(_10369_));
 sky130_fd_sc_hd__a22o_1 _20504_ (.A1(_10202_),
    .A2(_10204_),
    .B1(_10363_),
    .B2(_10365_),
    .X(_10370_));
 sky130_fd_sc_hd__a22oi_4 _20505_ (.A1(_09869_),
    .A2(_10118_),
    .B1(_10366_),
    .B2(_10367_),
    .Y(_10371_));
 sky130_fd_sc_hd__nand4_2 _20506_ (.A(_09867_),
    .B(_10117_),
    .C(_10369_),
    .D(_10370_),
    .Y(_10372_));
 sky130_fd_sc_hd__a22oi_2 _20507_ (.A1(_09867_),
    .A2(_10117_),
    .B1(_10369_),
    .B2(_10370_),
    .Y(_10373_));
 sky130_fd_sc_hd__o2111ai_4 _20508_ (.A1(_09970_),
    .A2(_09866_),
    .B1(_09869_),
    .C1(_10366_),
    .D1(_10367_),
    .Y(_10374_));
 sky130_fd_sc_hd__a41oi_4 _20509_ (.A1(_09869_),
    .A2(_10118_),
    .A3(_10366_),
    .A4(_10367_),
    .B1(_10116_),
    .Y(_10375_));
 sky130_fd_sc_hd__o211ai_2 _20510_ (.A1(_10112_),
    .A2(_10113_),
    .B1(_10372_),
    .C1(_10374_),
    .Y(_10376_));
 sky130_fd_sc_hd__o22ai_2 _20511_ (.A1(_10108_),
    .A2(_10111_),
    .B1(_10371_),
    .B2(_10373_),
    .Y(_10377_));
 sky130_fd_sc_hd__o211ai_2 _20512_ (.A1(_10108_),
    .A2(_10111_),
    .B1(_10372_),
    .C1(_10374_),
    .Y(_10378_));
 sky130_fd_sc_hd__o22ai_2 _20513_ (.A1(_10112_),
    .A2(_10113_),
    .B1(_10371_),
    .B2(_10373_),
    .Y(_10380_));
 sky130_fd_sc_hd__o211ai_4 _20514_ (.A1(_09978_),
    .A2(_09982_),
    .B1(_10376_),
    .C1(_10377_),
    .Y(_10381_));
 sky130_fd_sc_hd__nand3_2 _20515_ (.A(_10380_),
    .B(_10026_),
    .C(_10378_),
    .Y(_10382_));
 sky130_fd_sc_hd__a32oi_2 _20516_ (.A1(_10380_),
    .A2(_10026_),
    .A3(_10378_),
    .B1(_09694_),
    .B2(_09689_),
    .Y(_10383_));
 sky130_fd_sc_hd__o211a_1 _20517_ (.A1(_09688_),
    .A2(_09695_),
    .B1(_10381_),
    .C1(_10382_),
    .X(_10384_));
 sky130_fd_sc_hd__nand3_2 _20518_ (.A(_10025_),
    .B(_10381_),
    .C(_10382_),
    .Y(_10385_));
 sky130_fd_sc_hd__a21oi_2 _20519_ (.A1(_10381_),
    .A2(_10382_),
    .B1(_10025_),
    .Y(_10386_));
 sky130_fd_sc_hd__a21o_1 _20520_ (.A1(_10381_),
    .A2(_10382_),
    .B1(_10025_),
    .X(_10387_));
 sky130_fd_sc_hd__a221oi_2 _20521_ (.A1(_10383_),
    .A2(_10381_),
    .B1(_09992_),
    .B2(_09987_),
    .C1(_10386_),
    .Y(_10388_));
 sky130_fd_sc_hd__nand3_2 _20522_ (.A(_10024_),
    .B(_10385_),
    .C(_10387_),
    .Y(_10389_));
 sky130_fd_sc_hd__o22a_1 _20523_ (.A1(_09988_),
    .A2(_10023_),
    .B1(_10384_),
    .B2(_10386_),
    .X(_10391_));
 sky130_fd_sc_hd__o22ai_4 _20524_ (.A1(_09988_),
    .A2(_10023_),
    .B1(_10384_),
    .B2(_10386_),
    .Y(_10392_));
 sky130_fd_sc_hd__o211a_1 _20525_ (.A1(_09670_),
    .A2(_09674_),
    .B1(_10389_),
    .C1(_10392_),
    .X(_10393_));
 sky130_fd_sc_hd__o211ai_2 _20526_ (.A1(_09670_),
    .A2(_09674_),
    .B1(_10389_),
    .C1(_10392_),
    .Y(_10394_));
 sky130_fd_sc_hd__a21oi_1 _20527_ (.A1(_10389_),
    .A2(_10392_),
    .B1(_10022_),
    .Y(_10395_));
 sky130_fd_sc_hd__o22ai_1 _20528_ (.A1(_09671_),
    .A2(_10021_),
    .B1(_10388_),
    .B2(_10391_),
    .Y(_10396_));
 sky130_fd_sc_hd__nand3_2 _20529_ (.A(_10396_),
    .B(_10020_),
    .C(_10394_),
    .Y(_10397_));
 sky130_fd_sc_hd__o22a_1 _20530_ (.A1(_10001_),
    .A2(_10019_),
    .B1(_10393_),
    .B2(_10395_),
    .X(_10398_));
 sky130_fd_sc_hd__o22ai_2 _20531_ (.A1(_10001_),
    .A2(_10019_),
    .B1(_10393_),
    .B2(_10395_),
    .Y(_10399_));
 sky130_fd_sc_hd__nand2_1 _20532_ (.A(_10397_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__o2bb2a_1 _20533_ (.A1_N(_10012_),
    .A2_N(_10018_),
    .B1(_10013_),
    .B2(_10008_),
    .X(_10402_));
 sky130_fd_sc_hd__xor2_1 _20534_ (.A(_10400_),
    .B(_10402_),
    .X(net93));
 sky130_fd_sc_hd__a21o_1 _20535_ (.A1(_10392_),
    .A2(_10022_),
    .B1(_10388_),
    .X(_10403_));
 sky130_fd_sc_hd__and2_1 _20536_ (.A(_10096_),
    .B(_10063_),
    .X(_10404_));
 sky130_fd_sc_hd__a41o_1 _20537_ (.A1(_09663_),
    .A2(_10089_),
    .A3(_10090_),
    .A4(_10091_),
    .B1(_10063_),
    .X(_10405_));
 sky130_fd_sc_hd__a32o_1 _20538_ (.A1(_10087_),
    .A2(_10088_),
    .A3(_10092_),
    .B1(_10095_),
    .B2(_10064_),
    .X(_10406_));
 sky130_fd_sc_hd__a21boi_1 _20539_ (.A1(_10025_),
    .A2(_10382_),
    .B1_N(_10381_),
    .Y(_10407_));
 sky130_fd_sc_hd__nand2_1 _20540_ (.A(_10381_),
    .B(_10385_),
    .Y(_10408_));
 sky130_fd_sc_hd__o31a_2 _20541_ (.A1(_09637_),
    .A2(_09679_),
    .A3(_10102_),
    .B1(_10106_),
    .X(_10409_));
 sky130_fd_sc_hd__inv_2 _20542_ (.A(_10409_),
    .Y(_10410_));
 sky130_fd_sc_hd__a32oi_4 _20543_ (.A1(_10207_),
    .A2(_10359_),
    .A3(_10360_),
    .B1(_10204_),
    .B2(_10202_),
    .Y(_10412_));
 sky130_fd_sc_hd__a32o_1 _20544_ (.A1(_10207_),
    .A2(_10359_),
    .A3(_10360_),
    .B1(_10204_),
    .B2(_10202_),
    .X(_10413_));
 sky130_fd_sc_hd__a32o_1 _20545_ (.A1(_10208_),
    .A2(_10361_),
    .A3(_10362_),
    .B1(_10363_),
    .B2(_10205_),
    .X(_10414_));
 sky130_fd_sc_hd__a22oi_4 _20546_ (.A1(_10256_),
    .A2(_10253_),
    .B1(_10262_),
    .B2(_10260_),
    .Y(_10415_));
 sky130_fd_sc_hd__o2bb2ai_2 _20547_ (.A1_N(_10256_),
    .A2_N(_10253_),
    .B1(_10261_),
    .B2(_10259_),
    .Y(_10416_));
 sky130_fd_sc_hd__a21oi_4 _20548_ (.A1(_10125_),
    .A2(_10132_),
    .B1(_10133_),
    .Y(_10417_));
 sky130_fd_sc_hd__a21oi_2 _20549_ (.A1(_10219_),
    .A2(_10221_),
    .B1(_10217_),
    .Y(_10418_));
 sky130_fd_sc_hd__a21o_1 _20550_ (.A1(_10219_),
    .A2(_10221_),
    .B1(_10217_),
    .X(_10419_));
 sky130_fd_sc_hd__o22a_1 _20551_ (.A1(_04113_),
    .A2(_04218_),
    .B1(_05077_),
    .B2(_04216_),
    .X(_10420_));
 sky130_fd_sc_hd__a32o_1 _20552_ (.A1(net210),
    .A2(net183),
    .A3(net281),
    .B1(_04217_),
    .B2(net13),
    .X(_10421_));
 sky130_fd_sc_hd__nand3_4 _20553_ (.A(net182),
    .B(net179),
    .C(net285),
    .Y(_10423_));
 sky130_fd_sc_hd__or3_4 _20554_ (.A(net39),
    .B(_04135_),
    .C(_04037_),
    .X(_10424_));
 sky130_fd_sc_hd__o211ai_4 _20555_ (.A1(net184),
    .A2(_05551_),
    .B1(_02858_),
    .C1(net178),
    .Y(_10425_));
 sky130_fd_sc_hd__or3b_2 _20556_ (.A(net38),
    .B(_04146_),
    .C_N(net37),
    .X(_10426_));
 sky130_fd_sc_hd__a22oi_4 _20557_ (.A1(_10423_),
    .A2(_10424_),
    .B1(_10425_),
    .B2(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__a22o_2 _20558_ (.A1(_10423_),
    .A2(_10424_),
    .B1(_10425_),
    .B2(_10426_),
    .X(_10428_));
 sky130_fd_sc_hd__o2111a_2 _20559_ (.A1(_04146_),
    .A2(_02891_),
    .B1(_10423_),
    .C1(_10424_),
    .D1(_10425_),
    .X(_10429_));
 sky130_fd_sc_hd__o2111ai_4 _20560_ (.A1(_04146_),
    .A2(_02891_),
    .B1(_10423_),
    .C1(_10424_),
    .D1(_10425_),
    .Y(_10430_));
 sky130_fd_sc_hd__o21ai_4 _20561_ (.A1(_10427_),
    .A2(_10429_),
    .B1(_10420_),
    .Y(_10431_));
 sky130_fd_sc_hd__nand2_2 _20562_ (.A(_10421_),
    .B(_10428_),
    .Y(_10432_));
 sky130_fd_sc_hd__and3_1 _20563_ (.A(_10421_),
    .B(_10428_),
    .C(_10430_),
    .X(_10434_));
 sky130_fd_sc_hd__nand3_2 _20564_ (.A(_10421_),
    .B(_10428_),
    .C(_10430_),
    .Y(_10435_));
 sky130_fd_sc_hd__o21ai_1 _20565_ (.A1(_10429_),
    .A2(_10432_),
    .B1(_10431_),
    .Y(_10436_));
 sky130_fd_sc_hd__a21oi_4 _20566_ (.A1(_10431_),
    .A2(_10435_),
    .B1(_10419_),
    .Y(_10437_));
 sky130_fd_sc_hd__o211a_4 _20567_ (.A1(_10429_),
    .A2(_10432_),
    .B1(_10431_),
    .C1(_10419_),
    .X(_10438_));
 sky130_fd_sc_hd__o221ai_4 _20568_ (.A1(_10429_),
    .A2(_10432_),
    .B1(_10217_),
    .B2(_10224_),
    .C1(_10431_),
    .Y(_10439_));
 sky130_fd_sc_hd__a21oi_2 _20569_ (.A1(_10436_),
    .A2(_10418_),
    .B1(_10417_),
    .Y(_10440_));
 sky130_fd_sc_hd__o2bb2ai_2 _20570_ (.A1_N(_10418_),
    .A2_N(_10436_),
    .B1(_10133_),
    .B2(_10135_),
    .Y(_10441_));
 sky130_fd_sc_hd__o21ai_2 _20571_ (.A1(_10437_),
    .A2(_10438_),
    .B1(_10417_),
    .Y(_10442_));
 sky130_fd_sc_hd__nand3b_1 _20572_ (.A_N(_10437_),
    .B(_10439_),
    .C(_10417_),
    .Y(_10443_));
 sky130_fd_sc_hd__o22ai_2 _20573_ (.A1(_10133_),
    .A2(_10135_),
    .B1(_10437_),
    .B2(_10438_),
    .Y(_10445_));
 sky130_fd_sc_hd__o41ai_4 _20574_ (.A1(_09805_),
    .A2(_10121_),
    .A3(_10135_),
    .A4(_10138_),
    .B1(_10144_),
    .Y(_10446_));
 sky130_fd_sc_hd__a21oi_1 _20575_ (.A1(_10120_),
    .A2(_10142_),
    .B1(_10140_),
    .Y(_10447_));
 sky130_fd_sc_hd__nand3_2 _20576_ (.A(_10443_),
    .B(_10445_),
    .C(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__inv_2 _20577_ (.A(_10448_),
    .Y(_10449_));
 sky130_fd_sc_hd__o211a_1 _20578_ (.A1(_10438_),
    .A2(_10441_),
    .B1(_10446_),
    .C1(_10442_),
    .X(_10450_));
 sky130_fd_sc_hd__o211ai_4 _20579_ (.A1(_10438_),
    .A2(_10441_),
    .B1(_10446_),
    .C1(_10442_),
    .Y(_10451_));
 sky130_fd_sc_hd__and3_1 _20580_ (.A(_04102_),
    .B(net42),
    .C(net9),
    .X(_10452_));
 sky130_fd_sc_hd__o311a_1 _20581_ (.A1(net7),
    .A2(net248),
    .A3(_04407_),
    .B1(net243),
    .C1(net222),
    .X(_10453_));
 sky130_fd_sc_hd__a31o_1 _20582_ (.A1(net188),
    .A2(net222),
    .A3(net243),
    .B1(_10452_),
    .X(_10454_));
 sky130_fd_sc_hd__nor2_1 _20583_ (.A(_04091_),
    .B(_04270_),
    .Y(_10456_));
 sky130_fd_sc_hd__o311a_1 _20584_ (.A1(net7),
    .A2(net248),
    .A3(_04787_),
    .B1(net280),
    .C1(net214),
    .X(_10457_));
 sky130_fd_sc_hd__a31oi_2 _20585_ (.A1(net214),
    .A2(net280),
    .A3(net184),
    .B1(_10456_),
    .Y(_10458_));
 sky130_fd_sc_hd__o211ai_2 _20586_ (.A1(net231),
    .A2(_04557_),
    .B1(net279),
    .C1(net218),
    .Y(_10459_));
 sky130_fd_sc_hd__or3b_1 _20587_ (.A(net42),
    .B(_04080_),
    .C_N(net41),
    .X(_10460_));
 sky130_fd_sc_hd__o31ai_2 _20588_ (.A1(net216),
    .A2(_04481_),
    .A3(_04554_),
    .B1(_10460_),
    .Y(_10461_));
 sky130_fd_sc_hd__a21oi_1 _20589_ (.A1(_10459_),
    .A2(_10460_),
    .B1(_10458_),
    .Y(_10462_));
 sky130_fd_sc_hd__o21ai_4 _20590_ (.A1(_10456_),
    .A2(_10457_),
    .B1(_10461_),
    .Y(_10463_));
 sky130_fd_sc_hd__o211ai_4 _20591_ (.A1(_04080_),
    .A2(_04483_),
    .B1(_10459_),
    .C1(_10458_),
    .Y(_10464_));
 sky130_fd_sc_hd__a21oi_2 _20592_ (.A1(_10463_),
    .A2(_10464_),
    .B1(_10454_),
    .Y(_10465_));
 sky130_fd_sc_hd__a211o_2 _20593_ (.A1(_10463_),
    .A2(_10464_),
    .B1(_10452_),
    .C1(_10453_),
    .X(_10467_));
 sky130_fd_sc_hd__o211a_1 _20594_ (.A1(_10452_),
    .A2(_10453_),
    .B1(_10463_),
    .C1(_10464_),
    .X(_10468_));
 sky130_fd_sc_hd__o211ai_4 _20595_ (.A1(_10452_),
    .A2(_10453_),
    .B1(_10463_),
    .C1(_10464_),
    .Y(_10469_));
 sky130_fd_sc_hd__o22ai_4 _20596_ (.A1(_10177_),
    .A2(_10180_),
    .B1(_10465_),
    .B2(_10468_),
    .Y(_10470_));
 sky130_fd_sc_hd__nand3_4 _20597_ (.A(_10467_),
    .B(_10469_),
    .C(_10182_),
    .Y(_10471_));
 sky130_fd_sc_hd__a32o_1 _20598_ (.A1(_02421_),
    .A2(net248),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net6),
    .X(_10472_));
 sky130_fd_sc_hd__and3_1 _20599_ (.A(_04124_),
    .B(net43),
    .C(net8),
    .X(_10473_));
 sky130_fd_sc_hd__a31oi_4 _20600_ (.A1(net229),
    .A2(net228),
    .A3(net242),
    .B1(_10473_),
    .Y(_10474_));
 sky130_fd_sc_hd__a31o_1 _20601_ (.A1(net229),
    .A2(net228),
    .A3(net242),
    .B1(_10473_),
    .X(_10475_));
 sky130_fd_sc_hd__nor2_1 _20602_ (.A(_04048_),
    .B(_05229_),
    .Y(_10476_));
 sky130_fd_sc_hd__o32a_1 _20603_ (.A1(_05226_),
    .A2(_03957_),
    .A3(_03951_),
    .B1(_04048_),
    .B2(_05229_),
    .X(_10478_));
 sky130_fd_sc_hd__a31o_1 _20604_ (.A1(_03952_),
    .A2(net231),
    .A3(net276),
    .B1(_10476_),
    .X(_10479_));
 sky130_fd_sc_hd__nand2_1 _20605_ (.A(_10475_),
    .B(_10479_),
    .Y(_10480_));
 sky130_fd_sc_hd__o221a_1 _20606_ (.A1(_03961_),
    .A2(_05226_),
    .B1(_05229_),
    .B2(_04048_),
    .C1(_10474_),
    .X(_10481_));
 sky130_fd_sc_hd__nand2_1 _20607_ (.A(_10474_),
    .B(_10478_),
    .Y(_10482_));
 sky130_fd_sc_hd__o221a_1 _20608_ (.A1(_02475_),
    .A2(_05463_),
    .B1(_05465_),
    .B2(_04026_),
    .C1(_10480_),
    .X(_10483_));
 sky130_fd_sc_hd__o21ai_1 _20609_ (.A1(_10475_),
    .A2(_10479_),
    .B1(_10472_),
    .Y(_10484_));
 sky130_fd_sc_hd__o21ai_4 _20610_ (.A1(_10474_),
    .A2(_10478_),
    .B1(_10484_),
    .Y(_10485_));
 sky130_fd_sc_hd__a21oi_1 _20611_ (.A1(_10480_),
    .A2(_10482_),
    .B1(_10472_),
    .Y(_10486_));
 sky130_fd_sc_hd__a21oi_4 _20612_ (.A1(_10480_),
    .A2(_10485_),
    .B1(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__a21oi_2 _20613_ (.A1(_10470_),
    .A2(_10471_),
    .B1(_10487_),
    .Y(_10489_));
 sky130_fd_sc_hd__and2_1 _20614_ (.A(_10470_),
    .B(_10487_),
    .X(_10490_));
 sky130_fd_sc_hd__nand2_2 _20615_ (.A(_10470_),
    .B(_10487_),
    .Y(_10491_));
 sky130_fd_sc_hd__and3_1 _20616_ (.A(_10470_),
    .B(_10471_),
    .C(_10487_),
    .X(_10492_));
 sky130_fd_sc_hd__a21oi_1 _20617_ (.A1(_10490_),
    .A2(_10471_),
    .B1(_10489_),
    .Y(_10493_));
 sky130_fd_sc_hd__a21o_1 _20618_ (.A1(_10490_),
    .A2(_10471_),
    .B1(_10489_),
    .X(_10494_));
 sky130_fd_sc_hd__nand2_1 _20619_ (.A(_10493_),
    .B(_10448_),
    .Y(_10495_));
 sky130_fd_sc_hd__o2bb2ai_1 _20620_ (.A1_N(_10448_),
    .A2_N(_10451_),
    .B1(_10489_),
    .B2(_10492_),
    .Y(_10496_));
 sky130_fd_sc_hd__o211ai_2 _20621_ (.A1(_10489_),
    .A2(_10492_),
    .B1(_10448_),
    .C1(_10451_),
    .Y(_10497_));
 sky130_fd_sc_hd__a21o_1 _20622_ (.A1(_10448_),
    .A2(_10451_),
    .B1(_10494_),
    .X(_10498_));
 sky130_fd_sc_hd__nand3_4 _20623_ (.A(_10498_),
    .B(_10415_),
    .C(_10497_),
    .Y(_10500_));
 sky130_fd_sc_hd__o211ai_4 _20624_ (.A1(_10450_),
    .A2(_10495_),
    .B1(_10496_),
    .C1(_10416_),
    .Y(_10501_));
 sky130_fd_sc_hd__o31a_1 _20625_ (.A1(_10191_),
    .A2(_10193_),
    .A3(_10150_),
    .B1(_10149_),
    .X(_10502_));
 sky130_fd_sc_hd__o21ai_2 _20626_ (.A1(_10150_),
    .A2(_10195_),
    .B1(_10149_),
    .Y(_10503_));
 sky130_fd_sc_hd__a21o_1 _20627_ (.A1(_10500_),
    .A2(_10501_),
    .B1(_10503_),
    .X(_10504_));
 sky130_fd_sc_hd__nand3_1 _20628_ (.A(_10500_),
    .B(_10501_),
    .C(_10503_),
    .Y(_10505_));
 sky130_fd_sc_hd__a21oi_1 _20629_ (.A1(_10500_),
    .A2(_10501_),
    .B1(_10502_),
    .Y(_10506_));
 sky130_fd_sc_hd__a22o_1 _20630_ (.A1(_10149_),
    .A2(_10197_),
    .B1(_10500_),
    .B2(_10501_),
    .X(_10507_));
 sky130_fd_sc_hd__o2111a_1 _20631_ (.A1(_10195_),
    .A2(_10150_),
    .B1(_10149_),
    .C1(_10501_),
    .D1(_10500_),
    .X(_10508_));
 sky130_fd_sc_hd__o2111ai_1 _20632_ (.A1(_10195_),
    .A2(_10150_),
    .B1(_10149_),
    .C1(_10501_),
    .D1(_10500_),
    .Y(_10509_));
 sky130_fd_sc_hd__nand2_1 _20633_ (.A(_10507_),
    .B(_10509_),
    .Y(_10511_));
 sky130_fd_sc_hd__nand2_2 _20634_ (.A(_10504_),
    .B(_10505_),
    .Y(_10512_));
 sky130_fd_sc_hd__a22oi_2 _20635_ (.A1(_10351_),
    .A2(_10353_),
    .B1(_10264_),
    .B2(_10267_),
    .Y(_10513_));
 sky130_fd_sc_hd__o2bb2ai_4 _20636_ (.A1_N(_10351_),
    .A2_N(_10353_),
    .B1(_10263_),
    .B2(_10266_),
    .Y(_10514_));
 sky130_fd_sc_hd__o211ai_2 _20637_ (.A1(_10272_),
    .A2(_10307_),
    .B1(_10343_),
    .C1(_10345_),
    .Y(_10515_));
 sky130_fd_sc_hd__nand3_1 _20638_ (.A(_10310_),
    .B(_10339_),
    .C(_10341_),
    .Y(_10516_));
 sky130_fd_sc_hd__o21ai_1 _20639_ (.A1(_10272_),
    .A2(_10307_),
    .B1(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__o21ai_4 _20640_ (.A1(_10271_),
    .A2(_10308_),
    .B1(_10515_),
    .Y(_10518_));
 sky130_fd_sc_hd__o21ai_1 _20641_ (.A1(net147),
    .A2(_10274_),
    .B1(_10277_),
    .Y(_10519_));
 sky130_fd_sc_hd__a31o_1 _20642_ (.A1(_08882_),
    .A2(_09298_),
    .A3(_10277_),
    .B1(_10274_),
    .X(_10520_));
 sky130_fd_sc_hd__o22a_1 _20643_ (.A1(_05457_),
    .A2(_08658_),
    .B1(_08660_),
    .B2(_03725_),
    .X(_10522_));
 sky130_fd_sc_hd__a32o_2 _20644_ (.A1(_05414_),
    .A2(_05446_),
    .A3(_08657_),
    .B1(_08659_),
    .B2(net28),
    .X(_10523_));
 sky130_fd_sc_hd__a31oi_2 _20645_ (.A1(net162),
    .A2(net33),
    .A3(net319),
    .B1(_10523_),
    .Y(_10524_));
 sky130_fd_sc_hd__a31o_1 _20646_ (.A1(net162),
    .A2(net33),
    .A3(net319),
    .B1(_10523_),
    .X(_10525_));
 sky130_fd_sc_hd__and3_2 _20647_ (.A(_10523_),
    .B(net33),
    .C(net319),
    .X(_10526_));
 sky130_fd_sc_hd__nand3_2 _20648_ (.A(_10523_),
    .B(net33),
    .C(net319),
    .Y(_10527_));
 sky130_fd_sc_hd__o21ai_1 _20649_ (.A1(_10524_),
    .A2(_10526_),
    .B1(net147),
    .Y(_10528_));
 sky130_fd_sc_hd__a21oi_2 _20650_ (.A1(_08878_),
    .A2(_10522_),
    .B1(net147),
    .Y(_10529_));
 sky130_fd_sc_hd__a22o_2 _20651_ (.A1(_08882_),
    .A2(_09298_),
    .B1(_10522_),
    .B2(_08878_),
    .X(_10530_));
 sky130_fd_sc_hd__o22ai_2 _20652_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_10524_),
    .B2(_10526_),
    .Y(_10531_));
 sky130_fd_sc_hd__nand3_1 _20653_ (.A(_10525_),
    .B(_10527_),
    .C(net148),
    .Y(_10533_));
 sky130_fd_sc_hd__nand3_4 _20654_ (.A(_10528_),
    .B(_10530_),
    .C(_10519_),
    .Y(_10534_));
 sky130_fd_sc_hd__nand3_2 _20655_ (.A(_10520_),
    .B(_10531_),
    .C(_10533_),
    .Y(_10535_));
 sky130_fd_sc_hd__nand2_1 _20656_ (.A(_10534_),
    .B(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__nor2_1 _20657_ (.A(net25),
    .B(_04900_),
    .Y(_10537_));
 sky130_fd_sc_hd__a21oi_4 _20658_ (.A1(net162),
    .A2(_10537_),
    .B1(_10290_),
    .Y(_10538_));
 sky130_fd_sc_hd__a31o_2 _20659_ (.A1(_04277_),
    .A2(net162),
    .A3(_04889_),
    .B1(_10290_),
    .X(_10539_));
 sky130_fd_sc_hd__o2111a_4 _20660_ (.A1(_04900_),
    .A2(net151),
    .B1(_09754_),
    .C1(_10292_),
    .D1(_10295_),
    .X(_10540_));
 sky130_fd_sc_hd__o2111ai_4 _20661_ (.A1(_04900_),
    .A2(net151),
    .B1(_09754_),
    .C1(_10292_),
    .D1(_10295_),
    .Y(_10541_));
 sky130_fd_sc_hd__a21oi_4 _20662_ (.A1(_09754_),
    .A2(_10295_),
    .B1(_10538_),
    .Y(_10542_));
 sky130_fd_sc_hd__a31o_4 _20663_ (.A1(_09754_),
    .A2(_09759_),
    .A3(_10294_),
    .B1(_10538_),
    .X(_10544_));
 sky130_fd_sc_hd__nor2_8 _20664_ (.A(net140),
    .B(net136),
    .Y(_10545_));
 sky130_fd_sc_hd__nand2_8 _20665_ (.A(net139),
    .B(_10544_),
    .Y(_10546_));
 sky130_fd_sc_hd__o2bb2ai_2 _20666_ (.A1_N(_10534_),
    .A2_N(_10535_),
    .B1(_10540_),
    .B2(net137),
    .Y(_10547_));
 sky130_fd_sc_hd__nand3_2 _20667_ (.A(_10535_),
    .B(_10541_),
    .C(net134),
    .Y(_10548_));
 sky130_fd_sc_hd__nand4_4 _20668_ (.A(_10534_),
    .B(_10535_),
    .C(_10541_),
    .D(net134),
    .Y(_10549_));
 sky130_fd_sc_hd__nand2_2 _20669_ (.A(_10547_),
    .B(_10549_),
    .Y(_10550_));
 sky130_fd_sc_hd__o21a_2 _20670_ (.A1(_10282_),
    .A2(_10285_),
    .B1(_10305_),
    .X(_10551_));
 sky130_fd_sc_hd__o21ai_2 _20671_ (.A1(_10282_),
    .A2(_10285_),
    .B1(_10305_),
    .Y(_10552_));
 sky130_fd_sc_hd__a21oi_1 _20672_ (.A1(_10547_),
    .A2(_10549_),
    .B1(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__a21o_1 _20673_ (.A1(_10547_),
    .A2(_10549_),
    .B1(_10552_),
    .X(_10555_));
 sky130_fd_sc_hd__a22oi_4 _20674_ (.A1(_10288_),
    .A2(_10305_),
    .B1(_10536_),
    .B2(_10546_),
    .Y(_10556_));
 sky130_fd_sc_hd__nand3_1 _20675_ (.A(_10547_),
    .B(_10549_),
    .C(_10552_),
    .Y(_10557_));
 sky130_fd_sc_hd__a21oi_1 _20676_ (.A1(_10556_),
    .A2(_10549_),
    .B1(_10553_),
    .Y(_10558_));
 sky130_fd_sc_hd__nand2_1 _20677_ (.A(_10555_),
    .B(_10557_),
    .Y(_10559_));
 sky130_fd_sc_hd__o311a_1 _20678_ (.A1(_03958_),
    .A2(_05927_),
    .A3(_07767_),
    .B1(_07771_),
    .C1(_06826_),
    .X(_10560_));
 sky130_fd_sc_hd__and3_1 _20679_ (.A(_03927_),
    .B(net22),
    .C(net61),
    .X(_10561_));
 sky130_fd_sc_hd__a31o_1 _20680_ (.A1(_07771_),
    .A2(_06826_),
    .A3(net165),
    .B1(_10561_),
    .X(_10562_));
 sky130_fd_sc_hd__o211ai_4 _20681_ (.A1(_07076_),
    .A2(_08206_),
    .B1(_05688_),
    .C1(_08204_),
    .Y(_10563_));
 sky130_fd_sc_hd__or3b_1 _20682_ (.A(net61),
    .B(_04256_),
    .C_N(net60),
    .X(_10564_));
 sky130_fd_sc_hd__nor2_8 _20683_ (.A(net319),
    .B(_05260_),
    .Y(_10566_));
 sky130_fd_sc_hd__or3b_1 _20684_ (.A(net60),
    .B(_04277_),
    .C_N(net59),
    .X(_10567_));
 sky130_fd_sc_hd__a21oi_2 _20685_ (.A1(net151),
    .A2(net158),
    .B1(_05238_),
    .Y(_10568_));
 sky130_fd_sc_hd__o21ai_1 _20686_ (.A1(_08664_),
    .A2(_08666_),
    .B1(_05227_),
    .Y(_10569_));
 sky130_fd_sc_hd__o2111ai_4 _20687_ (.A1(_04256_),
    .A2(_05720_),
    .B1(_10563_),
    .C1(_10567_),
    .D1(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__o2bb2a_2 _20688_ (.A1_N(_10563_),
    .A2_N(_10564_),
    .B1(_10566_),
    .B2(_10568_),
    .X(_10571_));
 sky130_fd_sc_hd__o2bb2ai_4 _20689_ (.A1_N(_10563_),
    .A2_N(_10564_),
    .B1(_10566_),
    .B2(_10568_),
    .Y(_10572_));
 sky130_fd_sc_hd__a21oi_2 _20690_ (.A1(_10570_),
    .A2(_10572_),
    .B1(_10562_),
    .Y(_10573_));
 sky130_fd_sc_hd__a21o_1 _20691_ (.A1(_10570_),
    .A2(_10572_),
    .B1(_10562_),
    .X(_10574_));
 sky130_fd_sc_hd__o211a_2 _20692_ (.A1(_10560_),
    .A2(_10561_),
    .B1(_10570_),
    .C1(_10572_),
    .X(_10575_));
 sky130_fd_sc_hd__o211ai_4 _20693_ (.A1(_10560_),
    .A2(_10561_),
    .B1(_10570_),
    .C1(_10572_),
    .Y(_10577_));
 sky130_fd_sc_hd__o22a_1 _20694_ (.A1(_10293_),
    .A2(_10297_),
    .B1(_10573_),
    .B2(_10575_),
    .X(_10578_));
 sky130_fd_sc_hd__o22ai_4 _20695_ (.A1(_10293_),
    .A2(_10297_),
    .B1(_10573_),
    .B2(_10575_),
    .Y(_10579_));
 sky130_fd_sc_hd__nand3_4 _20696_ (.A(_10574_),
    .B(_10577_),
    .C(_10300_),
    .Y(_10580_));
 sky130_fd_sc_hd__nor2_1 _20697_ (.A(_10327_),
    .B(_10322_),
    .Y(_10581_));
 sky130_fd_sc_hd__nor2_1 _20698_ (.A(_10323_),
    .B(_10326_),
    .Y(_10582_));
 sky130_fd_sc_hd__a21o_1 _20699_ (.A1(_10325_),
    .A2(_10327_),
    .B1(_10322_),
    .X(_10583_));
 sky130_fd_sc_hd__o2bb2ai_1 _20700_ (.A1_N(_10579_),
    .A2_N(_10580_),
    .B1(_10582_),
    .B2(_10322_),
    .Y(_10584_));
 sky130_fd_sc_hd__o211ai_2 _20701_ (.A1(_10323_),
    .A2(_10581_),
    .B1(_10580_),
    .C1(_10579_),
    .Y(_10585_));
 sky130_fd_sc_hd__o2bb2ai_4 _20702_ (.A1_N(_10579_),
    .A2_N(_10580_),
    .B1(_10581_),
    .B2(_10323_),
    .Y(_10586_));
 sky130_fd_sc_hd__o211ai_2 _20703_ (.A1(_10322_),
    .A2(_10582_),
    .B1(_10580_),
    .C1(_10579_),
    .Y(_10588_));
 sky130_fd_sc_hd__nand3_2 _20704_ (.A(_10558_),
    .B(_10584_),
    .C(_10585_),
    .Y(_10589_));
 sky130_fd_sc_hd__nand3_2 _20705_ (.A(_10559_),
    .B(_10586_),
    .C(_10588_),
    .Y(_10590_));
 sky130_fd_sc_hd__nand3_1 _20706_ (.A(_10559_),
    .B(_10584_),
    .C(_10585_),
    .Y(_10591_));
 sky130_fd_sc_hd__nand4_2 _20707_ (.A(_10555_),
    .B(_10557_),
    .C(_10586_),
    .D(_10588_),
    .Y(_10592_));
 sky130_fd_sc_hd__nand3_4 _20708_ (.A(_10518_),
    .B(_10589_),
    .C(_10590_),
    .Y(_10593_));
 sky130_fd_sc_hd__a21oi_4 _20709_ (.A1(_10589_),
    .A2(_10590_),
    .B1(_10518_),
    .Y(_10594_));
 sky130_fd_sc_hd__nand3_4 _20710_ (.A(_10517_),
    .B(_10591_),
    .C(_10592_),
    .Y(_10595_));
 sky130_fd_sc_hd__o32a_2 _20711_ (.A1(_01304_),
    .A2(net203),
    .A3(_05932_),
    .B1(_01326_),
    .B2(_04157_),
    .X(_10596_));
 sky130_fd_sc_hd__a32o_1 _20712_ (.A1(_05933_),
    .A2(_01293_),
    .A3(net174),
    .B1(_01315_),
    .B2(net16),
    .X(_10597_));
 sky130_fd_sc_hd__nor2_1 _20713_ (.A(_04168_),
    .B(_12363_),
    .Y(_10599_));
 sky130_fd_sc_hd__a31oi_4 _20714_ (.A1(net201),
    .A2(net173),
    .A3(_12330_),
    .B1(_10599_),
    .Y(_10600_));
 sky130_fd_sc_hd__o211ai_4 _20715_ (.A1(net174),
    .A2(_06451_),
    .B1(net252),
    .C1(net198),
    .Y(_10601_));
 sky130_fd_sc_hd__or3_1 _20716_ (.A(net35),
    .B(_04179_),
    .C(_03971_),
    .X(_10602_));
 sky130_fd_sc_hd__a21oi_4 _20717_ (.A1(_10601_),
    .A2(_10602_),
    .B1(_10600_),
    .Y(_10603_));
 sky130_fd_sc_hd__o221a_1 _20718_ (.A1(_04179_),
    .A2(_11804_),
    .B1(_06454_),
    .B2(_11782_),
    .C1(_10600_),
    .X(_10604_));
 sky130_fd_sc_hd__o211ai_2 _20719_ (.A1(_04179_),
    .A2(_11804_),
    .B1(_10601_),
    .C1(_10600_),
    .Y(_10605_));
 sky130_fd_sc_hd__o21a_1 _20720_ (.A1(_10603_),
    .A2(_10604_),
    .B1(_10596_),
    .X(_10606_));
 sky130_fd_sc_hd__o21ai_1 _20721_ (.A1(_10603_),
    .A2(_10604_),
    .B1(_10596_),
    .Y(_10607_));
 sky130_fd_sc_hd__nor3b_4 _20722_ (.A(_10596_),
    .B(_10603_),
    .C_N(_10605_),
    .Y(_10608_));
 sky130_fd_sc_hd__or3_1 _20723_ (.A(_10596_),
    .B(_10603_),
    .C(_10604_),
    .X(_10610_));
 sky130_fd_sc_hd__nor2_1 _20724_ (.A(_10606_),
    .B(_10608_),
    .Y(_10611_));
 sky130_fd_sc_hd__a21bo_1 _20725_ (.A1(_10230_),
    .A2(_10239_),
    .B1_N(_10240_),
    .X(_10612_));
 sky130_fd_sc_hd__a32oi_4 _20726_ (.A1(net194),
    .A2(net171),
    .A3(net289),
    .B1(_10335_),
    .B2(net19),
    .Y(_10613_));
 sky130_fd_sc_hd__a32o_1 _20727_ (.A1(net194),
    .A2(net171),
    .A3(net289),
    .B1(_10335_),
    .B2(net19),
    .X(_10614_));
 sky130_fd_sc_hd__nor2_2 _20728_ (.A(_04212_),
    .B(_08283_),
    .Y(_10615_));
 sky130_fd_sc_hd__or3b_1 _20729_ (.A(net64),
    .B(_04212_),
    .C_N(net63),
    .X(_10616_));
 sky130_fd_sc_hd__a221oi_2 _20730_ (.A1(net203),
    .A2(_07073_),
    .B1(net171),
    .B2(net20),
    .C1(_08261_),
    .Y(_10617_));
 sky130_fd_sc_hd__o221ai_4 _20731_ (.A1(net175),
    .A2(_07074_),
    .B1(_04212_),
    .B2(net189),
    .C1(net291),
    .Y(_10618_));
 sky130_fd_sc_hd__a31oi_4 _20732_ (.A1(_07072_),
    .A2(net168),
    .A3(net291),
    .B1(_10615_),
    .Y(_10619_));
 sky130_fd_sc_hd__a31oi_2 _20733_ (.A1(_03957_),
    .A2(_05926_),
    .A3(_07500_),
    .B1(_07669_),
    .Y(_10621_));
 sky130_fd_sc_hd__a22oi_4 _20734_ (.A1(net21),
    .A2(_07680_),
    .B1(_10621_),
    .B2(_07499_),
    .Y(_10622_));
 sky130_fd_sc_hd__o2bb2ai_1 _20735_ (.A1_N(_07499_),
    .A2_N(_10621_),
    .B1(_04223_),
    .B2(_07691_),
    .Y(_10623_));
 sky130_fd_sc_hd__a21oi_2 _20736_ (.A1(_10616_),
    .A2(_10618_),
    .B1(_10622_),
    .Y(_10624_));
 sky130_fd_sc_hd__o21ai_4 _20737_ (.A1(_10615_),
    .A2(_10617_),
    .B1(_10623_),
    .Y(_10625_));
 sky130_fd_sc_hd__nand3_2 _20738_ (.A(_10622_),
    .B(_10618_),
    .C(_10616_),
    .Y(_10626_));
 sky130_fd_sc_hd__a21oi_4 _20739_ (.A1(_10619_),
    .A2(_10622_),
    .B1(_10613_),
    .Y(_10627_));
 sky130_fd_sc_hd__and3_1 _20740_ (.A(_10614_),
    .B(_10625_),
    .C(_10626_),
    .X(_10628_));
 sky130_fd_sc_hd__o21ai_2 _20741_ (.A1(_10619_),
    .A2(_10622_),
    .B1(_10627_),
    .Y(_10629_));
 sky130_fd_sc_hd__a21oi_2 _20742_ (.A1(_10625_),
    .A2(_10626_),
    .B1(_10614_),
    .Y(_10630_));
 sky130_fd_sc_hd__a21o_1 _20743_ (.A1(_10625_),
    .A2(_10626_),
    .B1(_10614_),
    .X(_10632_));
 sky130_fd_sc_hd__a221oi_4 _20744_ (.A1(_10627_),
    .A2(_10625_),
    .B1(_10243_),
    .B2(_10240_),
    .C1(_10630_),
    .Y(_10633_));
 sky130_fd_sc_hd__nand3_2 _20745_ (.A(_10612_),
    .B(_10629_),
    .C(_10632_),
    .Y(_10634_));
 sky130_fd_sc_hd__a21oi_4 _20746_ (.A1(_10629_),
    .A2(_10632_),
    .B1(_10612_),
    .Y(_10635_));
 sky130_fd_sc_hd__o221ai_4 _20747_ (.A1(_10241_),
    .A2(_10229_),
    .B1(_10630_),
    .B2(_10628_),
    .C1(_10240_),
    .Y(_10636_));
 sky130_fd_sc_hd__o22ai_2 _20748_ (.A1(_10606_),
    .A2(_10608_),
    .B1(_10633_),
    .B2(_10635_),
    .Y(_10637_));
 sky130_fd_sc_hd__and3_2 _20749_ (.A(_10607_),
    .B(_10610_),
    .C(_10636_),
    .X(_10638_));
 sky130_fd_sc_hd__nand3_1 _20750_ (.A(_10636_),
    .B(_10611_),
    .C(_10634_),
    .Y(_10639_));
 sky130_fd_sc_hd__o21ai_2 _20751_ (.A1(_10633_),
    .A2(_10635_),
    .B1(_10611_),
    .Y(_10640_));
 sky130_fd_sc_hd__o211ai_2 _20752_ (.A1(_10606_),
    .A2(_10608_),
    .B1(_10634_),
    .C1(_10636_),
    .Y(_10641_));
 sky130_fd_sc_hd__a32oi_4 _20753_ (.A1(_10315_),
    .A2(_10329_),
    .A3(_10331_),
    .B1(_10337_),
    .B2(_10311_),
    .Y(_10643_));
 sky130_fd_sc_hd__o32ai_4 _20754_ (.A1(_10314_),
    .A2(_10328_),
    .A3(_10330_),
    .B1(_10312_),
    .B2(_10336_),
    .Y(_10644_));
 sky130_fd_sc_hd__nand3_4 _20755_ (.A(_10640_),
    .B(_10641_),
    .C(_10644_),
    .Y(_10645_));
 sky130_fd_sc_hd__nand3_4 _20756_ (.A(_10637_),
    .B(_10643_),
    .C(_10639_),
    .Y(_10646_));
 sky130_fd_sc_hd__o32a_1 _20757_ (.A1(_10242_),
    .A2(_10244_),
    .A3(_09834_),
    .B1(_10222_),
    .B2(_10224_),
    .X(_10647_));
 sky130_fd_sc_hd__a2bb2o_1 _20758_ (.A1_N(_10242_),
    .A2_N(_10246_),
    .B1(_10226_),
    .B2(_10250_),
    .X(_10648_));
 sky130_fd_sc_hd__o31a_1 _20759_ (.A1(_09834_),
    .A2(_10242_),
    .A3(_10244_),
    .B1(_10253_),
    .X(_10649_));
 sky130_fd_sc_hd__a31oi_1 _20760_ (.A1(_10640_),
    .A2(_10641_),
    .A3(_10644_),
    .B1(_10649_),
    .Y(_10650_));
 sky130_fd_sc_hd__and3_1 _20761_ (.A(_10645_),
    .B(_10646_),
    .C(_10648_),
    .X(_10651_));
 sky130_fd_sc_hd__nand2_1 _20762_ (.A(_10650_),
    .B(_10646_),
    .Y(_10652_));
 sky130_fd_sc_hd__a21oi_2 _20763_ (.A1(_10645_),
    .A2(_10646_),
    .B1(_10648_),
    .Y(_10654_));
 sky130_fd_sc_hd__a21o_1 _20764_ (.A1(_10645_),
    .A2(_10646_),
    .B1(_10648_),
    .X(_10655_));
 sky130_fd_sc_hd__o211a_1 _20765_ (.A1(_10249_),
    .A2(_10647_),
    .B1(_10646_),
    .C1(_10645_),
    .X(_10656_));
 sky130_fd_sc_hd__a21oi_2 _20766_ (.A1(_10645_),
    .A2(_10646_),
    .B1(_10649_),
    .Y(_10657_));
 sky130_fd_sc_hd__a21oi_1 _20767_ (.A1(_10646_),
    .A2(_10650_),
    .B1(_10654_),
    .Y(_10658_));
 sky130_fd_sc_hd__o211a_1 _20768_ (.A1(_10656_),
    .A2(_10657_),
    .B1(_10593_),
    .C1(_10595_),
    .X(_10659_));
 sky130_fd_sc_hd__o211ai_4 _20769_ (.A1(_10656_),
    .A2(_10657_),
    .B1(_10593_),
    .C1(_10595_),
    .Y(_10660_));
 sky130_fd_sc_hd__a21oi_1 _20770_ (.A1(_10593_),
    .A2(_10595_),
    .B1(_10658_),
    .Y(_10661_));
 sky130_fd_sc_hd__o2bb2ai_4 _20771_ (.A1_N(_10593_),
    .A2_N(_10595_),
    .B1(_10651_),
    .B2(_10654_),
    .Y(_10662_));
 sky130_fd_sc_hd__a22oi_4 _20772_ (.A1(_10354_),
    .A2(_10514_),
    .B1(_10660_),
    .B2(_10662_),
    .Y(_10663_));
 sky130_fd_sc_hd__o22ai_4 _20773_ (.A1(_10355_),
    .A2(_10513_),
    .B1(_10659_),
    .B2(_10661_),
    .Y(_10665_));
 sky130_fd_sc_hd__o2111a_2 _20774_ (.A1(_10351_),
    .A2(_10353_),
    .B1(_10514_),
    .C1(_10660_),
    .D1(_10662_),
    .X(_10666_));
 sky130_fd_sc_hd__o2111ai_4 _20775_ (.A1(_10351_),
    .A2(_10353_),
    .B1(_10514_),
    .C1(_10660_),
    .D1(_10662_),
    .Y(_10667_));
 sky130_fd_sc_hd__o21ai_2 _20776_ (.A1(_10506_),
    .A2(_10508_),
    .B1(_10667_),
    .Y(_10668_));
 sky130_fd_sc_hd__o211a_1 _20777_ (.A1(_10506_),
    .A2(_10508_),
    .B1(_10665_),
    .C1(_10667_),
    .X(_10669_));
 sky130_fd_sc_hd__o211ai_1 _20778_ (.A1(_10506_),
    .A2(_10508_),
    .B1(_10665_),
    .C1(_10667_),
    .Y(_10670_));
 sky130_fd_sc_hd__a21oi_1 _20779_ (.A1(_10665_),
    .A2(_10667_),
    .B1(_10511_),
    .Y(_10671_));
 sky130_fd_sc_hd__o2bb2ai_2 _20780_ (.A1_N(_10504_),
    .A2_N(_10505_),
    .B1(_10663_),
    .B2(_10666_),
    .Y(_10672_));
 sky130_fd_sc_hd__o21ai_1 _20781_ (.A1(_10663_),
    .A2(_10668_),
    .B1(_10672_),
    .Y(_10673_));
 sky130_fd_sc_hd__o2111ai_4 _20782_ (.A1(_10668_),
    .A2(_10663_),
    .B1(_10413_),
    .C1(_10365_),
    .D1(_10672_),
    .Y(_10674_));
 sky130_fd_sc_hd__a22oi_2 _20783_ (.A1(_10365_),
    .A2(_10413_),
    .B1(_10670_),
    .B2(_10672_),
    .Y(_10676_));
 sky130_fd_sc_hd__o22ai_4 _20784_ (.A1(_10364_),
    .A2(_10412_),
    .B1(_10669_),
    .B2(_10671_),
    .Y(_10677_));
 sky130_fd_sc_hd__o31ai_2 _20785_ (.A1(_09948_),
    .A2(_09957_),
    .A3(_10199_),
    .B1(_10201_),
    .Y(_10678_));
 sky130_fd_sc_hd__nand2_2 _20786_ (.A(_10053_),
    .B(_10057_),
    .Y(_10679_));
 sky130_fd_sc_hd__and3_1 _20787_ (.A(_04190_),
    .B(net49),
    .C(net3),
    .X(_10680_));
 sky130_fd_sc_hd__o311a_1 _20788_ (.A1(_04747_),
    .A2(net264),
    .A3(_11387_),
    .B1(net273),
    .C1(_11354_),
    .X(_10681_));
 sky130_fd_sc_hd__a31o_1 _20789_ (.A1(_11354_),
    .A2(net253),
    .A3(net273),
    .B1(_10680_),
    .X(_10682_));
 sky130_fd_sc_hd__or3b_1 _20790_ (.A(_04015_),
    .B(net48),
    .C_N(net47),
    .X(_10683_));
 sky130_fd_sc_hd__o211ai_4 _20791_ (.A1(net253),
    .A2(_00646_),
    .B1(net275),
    .C1(_00625_),
    .Y(_10684_));
 sky130_fd_sc_hd__nor2_1 _20792_ (.A(_04004_),
    .B(_06030_),
    .Y(_10685_));
 sky130_fd_sc_hd__o311a_1 _20793_ (.A1(net3),
    .A2(_09665_),
    .A3(_12988_),
    .B1(net274),
    .C1(net234),
    .X(_10687_));
 sky130_fd_sc_hd__a31oi_2 _20794_ (.A1(net234),
    .A2(net251),
    .A3(net274),
    .B1(_10685_),
    .Y(_10688_));
 sky130_fd_sc_hd__o211ai_4 _20795_ (.A1(_04015_),
    .A2(_05766_),
    .B1(_10684_),
    .C1(_10688_),
    .Y(_10689_));
 sky130_fd_sc_hd__o2bb2a_1 _20796_ (.A1_N(_10683_),
    .A2_N(_10684_),
    .B1(_10685_),
    .B2(_10687_),
    .X(_10690_));
 sky130_fd_sc_hd__o2bb2ai_2 _20797_ (.A1_N(_10683_),
    .A2_N(_10684_),
    .B1(_10685_),
    .B2(_10687_),
    .Y(_10691_));
 sky130_fd_sc_hd__a21oi_2 _20798_ (.A1(_10689_),
    .A2(_10691_),
    .B1(_10682_),
    .Y(_10692_));
 sky130_fd_sc_hd__and3_1 _20799_ (.A(_10682_),
    .B(_10689_),
    .C(_10691_),
    .X(_10693_));
 sky130_fd_sc_hd__o211ai_2 _20800_ (.A1(_10680_),
    .A2(_10681_),
    .B1(_10689_),
    .C1(_10691_),
    .Y(_10694_));
 sky130_fd_sc_hd__o21ai_1 _20801_ (.A1(_10154_),
    .A2(_10158_),
    .B1(_10151_),
    .Y(_10695_));
 sky130_fd_sc_hd__o21ai_2 _20802_ (.A1(_10153_),
    .A2(_10157_),
    .B1(_10695_),
    .Y(_10696_));
 sky130_fd_sc_hd__o21bai_4 _20803_ (.A1(_10692_),
    .A2(_10693_),
    .B1_N(_10696_),
    .Y(_10698_));
 sky130_fd_sc_hd__nand3b_4 _20804_ (.A_N(_10692_),
    .B(_10694_),
    .C(_10696_),
    .Y(_10699_));
 sky130_fd_sc_hd__inv_2 _20805_ (.A(_10699_),
    .Y(_10700_));
 sky130_fd_sc_hd__nor2_1 _20806_ (.A(_10029_),
    .B(_10034_),
    .Y(_10701_));
 sky130_fd_sc_hd__a41o_1 _20807_ (.A1(_10030_),
    .A2(_10031_),
    .A3(_10032_),
    .A4(_10033_),
    .B1(_10701_),
    .X(_10702_));
 sky130_fd_sc_hd__o2bb2ai_4 _20808_ (.A1_N(_10698_),
    .A2_N(_10699_),
    .B1(_10701_),
    .B2(_10036_),
    .Y(_10703_));
 sky130_fd_sc_hd__and3b_2 _20809_ (.A_N(_10702_),
    .B(_10699_),
    .C(_10698_),
    .X(_10704_));
 sky130_fd_sc_hd__nand3b_4 _20810_ (.A_N(_10702_),
    .B(_10699_),
    .C(_10698_),
    .Y(_10705_));
 sky130_fd_sc_hd__a32o_1 _20811_ (.A1(_10185_),
    .A2(_10186_),
    .A3(_10167_),
    .B1(_10165_),
    .B2(_10164_),
    .X(_10706_));
 sky130_fd_sc_hd__a31oi_4 _20812_ (.A1(_10168_),
    .A2(_10183_),
    .A3(_10184_),
    .B1(_10166_),
    .Y(_10707_));
 sky130_fd_sc_hd__a22oi_4 _20813_ (.A1(_10703_),
    .A2(_10705_),
    .B1(_10706_),
    .B2(_10187_),
    .Y(_10709_));
 sky130_fd_sc_hd__a22o_1 _20814_ (.A1(_10703_),
    .A2(_10705_),
    .B1(_10706_),
    .B2(_10187_),
    .X(_10710_));
 sky130_fd_sc_hd__o21ai_2 _20815_ (.A1(_10188_),
    .A2(_10707_),
    .B1(_10703_),
    .Y(_10711_));
 sky130_fd_sc_hd__o211a_1 _20816_ (.A1(_10188_),
    .A2(_10707_),
    .B1(_10705_),
    .C1(_10703_),
    .X(_10712_));
 sky130_fd_sc_hd__o211ai_2 _20817_ (.A1(_10188_),
    .A2(_10707_),
    .B1(_10705_),
    .C1(_10703_),
    .Y(_10713_));
 sky130_fd_sc_hd__a21bo_1 _20818_ (.A1(_10028_),
    .A2(_10045_),
    .B1_N(_10046_),
    .X(_10714_));
 sky130_fd_sc_hd__inv_2 _20819_ (.A(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__o21ai_4 _20820_ (.A1(_10709_),
    .A2(_10712_),
    .B1(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__o211ai_4 _20821_ (.A1(_10704_),
    .A2(_10711_),
    .B1(_10714_),
    .C1(_10710_),
    .Y(_10717_));
 sky130_fd_sc_hd__a21oi_4 _20822_ (.A1(_10716_),
    .A2(_10717_),
    .B1(_10679_),
    .Y(_10718_));
 sky130_fd_sc_hd__and3_1 _20823_ (.A(_10679_),
    .B(_10716_),
    .C(_10717_),
    .X(_10720_));
 sky130_fd_sc_hd__nand3_4 _20824_ (.A(_10679_),
    .B(_10716_),
    .C(_10717_),
    .Y(_10721_));
 sky130_fd_sc_hd__o2bb2a_1 _20825_ (.A1_N(_05874_),
    .A2_N(_08005_),
    .B1(_08007_),
    .B2(_03835_),
    .X(_10722_));
 sky130_fd_sc_hd__a32o_2 _20826_ (.A1(_05841_),
    .A2(net265),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net29),
    .X(_10723_));
 sky130_fd_sc_hd__and3b_1 _20827_ (.A_N(net54),
    .B(net53),
    .C(net30),
    .X(_10724_));
 sky130_fd_sc_hd__o311a_1 _20828_ (.A1(net26),
    .A2(_04452_),
    .A3(net264),
    .B1(_07642_),
    .C1(_06486_),
    .X(_10725_));
 sky130_fd_sc_hd__a31o_1 _20829_ (.A1(_06486_),
    .A2(net259),
    .A3(_07642_),
    .B1(_10724_),
    .X(_10726_));
 sky130_fd_sc_hd__a21o_1 _20830_ (.A1(_10067_),
    .A2(_10076_),
    .B1(_10074_),
    .X(_10727_));
 sky130_fd_sc_hd__a32oi_4 _20831_ (.A1(_07242_),
    .A2(net257),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net31),
    .Y(_10728_));
 sky130_fd_sc_hd__a32o_1 _20832_ (.A1(_07242_),
    .A2(net257),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net31),
    .X(_10729_));
 sky130_fd_sc_hd__or3_2 _20833_ (.A(net51),
    .B(_04190_),
    .C(_03960_),
    .X(_10731_));
 sky130_fd_sc_hd__o211ai_4 _20834_ (.A1(net259),
    .A2(_09665_),
    .B1(_06863_),
    .C1(_09698_),
    .Y(_10732_));
 sky130_fd_sc_hd__or3b_2 _20835_ (.A(_03949_),
    .B(net52),
    .C_N(net51),
    .X(_10733_));
 sky130_fd_sc_hd__o211ai_4 _20836_ (.A1(net259),
    .A2(_08656_),
    .B1(net269),
    .C1(_08700_),
    .Y(_10734_));
 sky130_fd_sc_hd__o2111a_1 _20837_ (.A1(_03960_),
    .A2(_06866_),
    .B1(_10732_),
    .C1(_10733_),
    .D1(_10734_),
    .X(_10735_));
 sky130_fd_sc_hd__o2111ai_1 _20838_ (.A1(_03960_),
    .A2(_06866_),
    .B1(_10732_),
    .C1(_10733_),
    .D1(_10734_),
    .Y(_10736_));
 sky130_fd_sc_hd__a22oi_4 _20839_ (.A1(_10731_),
    .A2(_10732_),
    .B1(_10733_),
    .B2(_10734_),
    .Y(_10737_));
 sky130_fd_sc_hd__a22o_1 _20840_ (.A1(_10731_),
    .A2(_10732_),
    .B1(_10733_),
    .B2(_10734_),
    .X(_10738_));
 sky130_fd_sc_hd__a41o_1 _20841_ (.A1(_10731_),
    .A2(_10732_),
    .A3(_10733_),
    .A4(_10734_),
    .B1(_10728_),
    .X(_10739_));
 sky130_fd_sc_hd__o21ai_1 _20842_ (.A1(_10728_),
    .A2(_10735_),
    .B1(_10738_),
    .Y(_10740_));
 sky130_fd_sc_hd__nand3_1 _20843_ (.A(_10738_),
    .B(_10728_),
    .C(_10736_),
    .Y(_10742_));
 sky130_fd_sc_hd__o21ai_1 _20844_ (.A1(_10735_),
    .A2(_10737_),
    .B1(_10729_),
    .Y(_10743_));
 sky130_fd_sc_hd__o21ai_1 _20845_ (.A1(_10735_),
    .A2(_10737_),
    .B1(_10728_),
    .Y(_10744_));
 sky130_fd_sc_hd__nand4_2 _20846_ (.A(_10075_),
    .B(_10079_),
    .C(_10742_),
    .D(_10743_),
    .Y(_10745_));
 sky130_fd_sc_hd__o211ai_4 _20847_ (.A1(_10739_),
    .A2(_10737_),
    .B1(_10727_),
    .C1(_10744_),
    .Y(_10746_));
 sky130_fd_sc_hd__a21oi_2 _20848_ (.A1(_10745_),
    .A2(_10746_),
    .B1(_10726_),
    .Y(_10747_));
 sky130_fd_sc_hd__and3_1 _20849_ (.A(_10726_),
    .B(_10745_),
    .C(_10746_),
    .X(_10748_));
 sky130_fd_sc_hd__o211ai_1 _20850_ (.A1(_10724_),
    .A2(_10725_),
    .B1(_10745_),
    .C1(_10746_),
    .Y(_10749_));
 sky130_fd_sc_hd__o21ai_1 _20851_ (.A1(_10081_),
    .A2(_10085_),
    .B1(_10084_),
    .Y(_10750_));
 sky130_fd_sc_hd__o21a_1 _20852_ (.A1(_10081_),
    .A2(_10085_),
    .B1(_10084_),
    .X(_10751_));
 sky130_fd_sc_hd__nor3_1 _20853_ (.A(_10747_),
    .B(_10748_),
    .C(_10751_),
    .Y(_10753_));
 sky130_fd_sc_hd__nand3b_1 _20854_ (.A_N(_10747_),
    .B(_10749_),
    .C(_10750_),
    .Y(_10754_));
 sky130_fd_sc_hd__o221a_1 _20855_ (.A1(_10081_),
    .A2(_10085_),
    .B1(_10747_),
    .B2(_10748_),
    .C1(_10084_),
    .X(_10755_));
 sky130_fd_sc_hd__o21ai_1 _20856_ (.A1(_10747_),
    .A2(_10748_),
    .B1(_10751_),
    .Y(_10756_));
 sky130_fd_sc_hd__nand2_2 _20857_ (.A(_10754_),
    .B(_10756_),
    .Y(_10757_));
 sky130_fd_sc_hd__xor2_1 _20858_ (.A(_10722_),
    .B(_10757_),
    .X(_10758_));
 sky130_fd_sc_hd__xor2_4 _20859_ (.A(_10723_),
    .B(_10757_),
    .X(_10759_));
 sky130_fd_sc_hd__o21ai_1 _20860_ (.A1(_10718_),
    .A2(_10720_),
    .B1(_10759_),
    .Y(_10760_));
 sky130_fd_sc_hd__nor2_1 _20861_ (.A(_10718_),
    .B(_10759_),
    .Y(_10761_));
 sky130_fd_sc_hd__nand3b_1 _20862_ (.A_N(_10718_),
    .B(_10758_),
    .C(_10721_),
    .Y(_10762_));
 sky130_fd_sc_hd__nand3b_1 _20863_ (.A_N(_10718_),
    .B(_10721_),
    .C(_10759_),
    .Y(_10764_));
 sky130_fd_sc_hd__o21ai_2 _20864_ (.A1(_10718_),
    .A2(_10720_),
    .B1(_10758_),
    .Y(_10765_));
 sky130_fd_sc_hd__and4_1 _20865_ (.A(_10201_),
    .B(_10202_),
    .C(_10764_),
    .D(_10765_),
    .X(_10766_));
 sky130_fd_sc_hd__nand4_4 _20866_ (.A(_10201_),
    .B(_10202_),
    .C(_10764_),
    .D(_10765_),
    .Y(_10767_));
 sky130_fd_sc_hd__nand3_2 _20867_ (.A(_10678_),
    .B(_10760_),
    .C(_10762_),
    .Y(_10768_));
 sky130_fd_sc_hd__inv_2 _20868_ (.A(_10768_),
    .Y(_10769_));
 sky130_fd_sc_hd__o21ai_4 _20869_ (.A1(_10059_),
    .A2(_10099_),
    .B1(_10062_),
    .Y(_10770_));
 sky130_fd_sc_hd__inv_2 _20870_ (.A(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__a21oi_1 _20871_ (.A1(_10767_),
    .A2(_10768_),
    .B1(_10771_),
    .Y(_10772_));
 sky130_fd_sc_hd__and3_1 _20872_ (.A(_10767_),
    .B(_10768_),
    .C(_10771_),
    .X(_10773_));
 sky130_fd_sc_hd__a21oi_1 _20873_ (.A1(_10767_),
    .A2(_10768_),
    .B1(_10770_),
    .Y(_10775_));
 sky130_fd_sc_hd__a21o_1 _20874_ (.A1(_10767_),
    .A2(_10768_),
    .B1(_10770_),
    .X(_10776_));
 sky130_fd_sc_hd__nor2_1 _20875_ (.A(_10766_),
    .B(_10771_),
    .Y(_10777_));
 sky130_fd_sc_hd__nand2_1 _20876_ (.A(_10767_),
    .B(_10770_),
    .Y(_10778_));
 sky130_fd_sc_hd__and3_1 _20877_ (.A(_10767_),
    .B(_10768_),
    .C(_10770_),
    .X(_10779_));
 sky130_fd_sc_hd__o21ai_2 _20878_ (.A1(_10778_),
    .A2(_10769_),
    .B1(_10776_),
    .Y(_10780_));
 sky130_fd_sc_hd__o2bb2ai_2 _20879_ (.A1_N(_10414_),
    .A2_N(_10673_),
    .B1(_10772_),
    .B2(_10773_),
    .Y(_10781_));
 sky130_fd_sc_hd__o2111ai_4 _20880_ (.A1(_10769_),
    .A2(_10778_),
    .B1(_10776_),
    .C1(_10674_),
    .D1(_10677_),
    .Y(_10782_));
 sky130_fd_sc_hd__o2bb2ai_1 _20881_ (.A1_N(_10674_),
    .A2_N(_10677_),
    .B1(_10775_),
    .B2(_10779_),
    .Y(_10783_));
 sky130_fd_sc_hd__nand3_2 _20882_ (.A(_10780_),
    .B(_10677_),
    .C(_10674_),
    .Y(_10784_));
 sky130_fd_sc_hd__o2bb2ai_2 _20883_ (.A1_N(_10674_),
    .A2_N(_10677_),
    .B1(_10772_),
    .B2(_10773_),
    .Y(_10786_));
 sky130_fd_sc_hd__o21ai_2 _20884_ (.A1(_10114_),
    .A2(_10371_),
    .B1(_10374_),
    .Y(_10787_));
 sky130_fd_sc_hd__nand3_4 _20885_ (.A(_10784_),
    .B(_10786_),
    .C(_10787_),
    .Y(_10788_));
 sky130_fd_sc_hd__o211ai_4 _20886_ (.A1(_10371_),
    .A2(_10375_),
    .B1(_10782_),
    .C1(_10783_),
    .Y(_10789_));
 sky130_fd_sc_hd__a22o_1 _20887_ (.A1(_10106_),
    .A2(_10110_),
    .B1(_10788_),
    .B2(_10789_),
    .X(_10790_));
 sky130_fd_sc_hd__nand4_2 _20888_ (.A(_10106_),
    .B(_10110_),
    .C(_10788_),
    .D(_10789_),
    .Y(_10791_));
 sky130_fd_sc_hd__a21o_1 _20889_ (.A1(_10788_),
    .A2(_10789_),
    .B1(_10410_),
    .X(_10792_));
 sky130_fd_sc_hd__a31o_1 _20890_ (.A1(_10787_),
    .A2(_10786_),
    .A3(_10784_),
    .B1(_10409_),
    .X(_10793_));
 sky130_fd_sc_hd__nand3_1 _20891_ (.A(_10410_),
    .B(_10788_),
    .C(_10789_),
    .Y(_10794_));
 sky130_fd_sc_hd__a22oi_4 _20892_ (.A1(_10381_),
    .A2(_10385_),
    .B1(_10790_),
    .B2(_10791_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand3_1 _20893_ (.A(_10408_),
    .B(_10792_),
    .C(_10794_),
    .Y(_10797_));
 sky130_fd_sc_hd__a21oi_1 _20894_ (.A1(_10792_),
    .A2(_10794_),
    .B1(_10408_),
    .Y(_10798_));
 sky130_fd_sc_hd__nand3_1 _20895_ (.A(_10790_),
    .B(_10791_),
    .C(_10407_),
    .Y(_10799_));
 sky130_fd_sc_hd__o22ai_2 _20896_ (.A1(_10094_),
    .A2(_10404_),
    .B1(_10795_),
    .B2(_10798_),
    .Y(_10800_));
 sky130_fd_sc_hd__nand2_1 _20897_ (.A(_10799_),
    .B(_10406_),
    .Y(_10801_));
 sky130_fd_sc_hd__o2bb2ai_1 _20898_ (.A1_N(_10096_),
    .A2_N(_10405_),
    .B1(_10795_),
    .B2(_10798_),
    .Y(_10802_));
 sky130_fd_sc_hd__o2111ai_1 _20899_ (.A1(_10063_),
    .A2(_10094_),
    .B1(_10096_),
    .C1(_10797_),
    .D1(_10799_),
    .Y(_10803_));
 sky130_fd_sc_hd__nand4_1 _20900_ (.A(_10389_),
    .B(_10394_),
    .C(_10802_),
    .D(_10803_),
    .Y(_10804_));
 sky130_fd_sc_hd__o211ai_4 _20901_ (.A1(_10795_),
    .A2(_10801_),
    .B1(_10800_),
    .C1(_10403_),
    .Y(_10805_));
 sky130_fd_sc_hd__nand2_1 _20902_ (.A(_10804_),
    .B(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__o2111ai_4 _20903_ (.A1(_10013_),
    .A2(_10008_),
    .B1(_10012_),
    .C1(_10397_),
    .D1(_10399_),
    .Y(_10808_));
 sky130_fd_sc_hd__o21a_1 _20904_ (.A1(_10008_),
    .A2(_10013_),
    .B1(_10397_),
    .X(_10809_));
 sky130_fd_sc_hd__o22ai_4 _20905_ (.A1(_10398_),
    .A2(_10809_),
    .B1(_10808_),
    .B2(_10015_),
    .Y(_10810_));
 sky130_fd_sc_hd__nor2_1 _20906_ (.A(_10016_),
    .B(_10808_),
    .Y(_10811_));
 sky130_fd_sc_hd__a21oi_2 _20907_ (.A1(_09171_),
    .A2(_10811_),
    .B1(_10810_),
    .Y(_10812_));
 sky130_fd_sc_hd__xor2_1 _20908_ (.A(_10806_),
    .B(_10812_),
    .X(net94));
 sky130_fd_sc_hd__o21ai_1 _20909_ (.A1(_10406_),
    .A2(_10795_),
    .B1(_10799_),
    .Y(_10813_));
 sky130_fd_sc_hd__a32o_1 _20910_ (.A1(_10408_),
    .A2(_10792_),
    .A3(_10794_),
    .B1(_10799_),
    .B2(_10406_),
    .X(_10814_));
 sky130_fd_sc_hd__o31a_1 _20911_ (.A1(_10747_),
    .A2(_10748_),
    .A3(_10751_),
    .B1(_10722_),
    .X(_10815_));
 sky130_fd_sc_hd__nor2_1 _20912_ (.A(_10722_),
    .B(_10755_),
    .Y(_10816_));
 sky130_fd_sc_hd__a21o_1 _20913_ (.A1(_10723_),
    .A2(_10756_),
    .B1(_10753_),
    .X(_10818_));
 sky130_fd_sc_hd__inv_2 _20914_ (.A(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__nand2_2 _20915_ (.A(_10789_),
    .B(_10409_),
    .Y(_10820_));
 sky130_fd_sc_hd__o32a_1 _20916_ (.A1(_10364_),
    .A2(_10412_),
    .A3(_10673_),
    .B1(_10676_),
    .B2(_10780_),
    .X(_10821_));
 sky130_fd_sc_hd__o21ai_2 _20917_ (.A1(_10676_),
    .A2(_10780_),
    .B1(_10674_),
    .Y(_10822_));
 sky130_fd_sc_hd__nand2_1 _20918_ (.A(_10502_),
    .B(_10501_),
    .Y(_10823_));
 sky130_fd_sc_hd__a21boi_2 _20919_ (.A1(_10500_),
    .A2(_10503_),
    .B1_N(_10501_),
    .Y(_10824_));
 sky130_fd_sc_hd__o2bb2a_2 _20920_ (.A1_N(_06541_),
    .A2_N(_08005_),
    .B1(_08007_),
    .B2(_03916_),
    .X(_10825_));
 sky130_fd_sc_hd__a32o_2 _20921_ (.A1(_07242_),
    .A2(net257),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net31),
    .X(_10826_));
 sky130_fd_sc_hd__o311a_1 _20922_ (.A1(_04747_),
    .A2(net264),
    .A3(_08656_),
    .B1(_07305_),
    .C1(_08700_),
    .X(_10827_));
 sky130_fd_sc_hd__and3_1 _20923_ (.A(_04234_),
    .B(net52),
    .C(net32),
    .X(_10829_));
 sky130_fd_sc_hd__a31o_1 _20924_ (.A1(net256),
    .A2(_08700_),
    .A3(_07305_),
    .B1(_10829_),
    .X(_10830_));
 sky130_fd_sc_hd__a31oi_4 _20925_ (.A1(net310),
    .A2(net294),
    .A3(net290),
    .B1(_07224_),
    .Y(_10831_));
 sky130_fd_sc_hd__a22oi_2 _20926_ (.A1(net2),
    .A2(_07225_),
    .B1(_09698_),
    .B2(_10831_),
    .Y(_10832_));
 sky130_fd_sc_hd__a22o_1 _20927_ (.A1(net2),
    .A2(_07225_),
    .B1(_09698_),
    .B2(_10831_),
    .X(_10833_));
 sky130_fd_sc_hd__nor2_1 _20928_ (.A(_03982_),
    .B(_06866_),
    .Y(_10834_));
 sky130_fd_sc_hd__or3_1 _20929_ (.A(net51),
    .B(_04190_),
    .C(_03982_),
    .X(_10835_));
 sky130_fd_sc_hd__a211oi_1 _20930_ (.A1(net255),
    .A2(net3),
    .B1(_06864_),
    .C1(_11420_),
    .Y(_10836_));
 sky130_fd_sc_hd__o211ai_2 _20931_ (.A1(net259),
    .A2(_11387_),
    .B1(_06863_),
    .C1(_11354_),
    .Y(_10837_));
 sky130_fd_sc_hd__o211ai_2 _20932_ (.A1(_03982_),
    .A2(_06866_),
    .B1(_10837_),
    .C1(_10832_),
    .Y(_10838_));
 sky130_fd_sc_hd__a21oi_1 _20933_ (.A1(_10835_),
    .A2(_10837_),
    .B1(_10832_),
    .Y(_10839_));
 sky130_fd_sc_hd__o21ai_1 _20934_ (.A1(_10834_),
    .A2(_10836_),
    .B1(_10833_),
    .Y(_10840_));
 sky130_fd_sc_hd__o211a_2 _20935_ (.A1(_10827_),
    .A2(_10829_),
    .B1(_10838_),
    .C1(_10840_),
    .X(_10841_));
 sky130_fd_sc_hd__a21oi_1 _20936_ (.A1(_10838_),
    .A2(_10840_),
    .B1(_10830_),
    .Y(_10842_));
 sky130_fd_sc_hd__a21o_1 _20937_ (.A1(_10838_),
    .A2(_10840_),
    .B1(_10830_),
    .X(_10843_));
 sky130_fd_sc_hd__nand2_1 _20938_ (.A(_10843_),
    .B(_10740_),
    .Y(_10844_));
 sky130_fd_sc_hd__nand3b_1 _20939_ (.A_N(_10841_),
    .B(_10843_),
    .C(_10740_),
    .Y(_10845_));
 sky130_fd_sc_hd__o21bai_4 _20940_ (.A1(_10841_),
    .A2(_10842_),
    .B1_N(_10740_),
    .Y(_10846_));
 sky130_fd_sc_hd__a21o_1 _20941_ (.A1(_10845_),
    .A2(_10846_),
    .B1(_10826_),
    .X(_10847_));
 sky130_fd_sc_hd__o211ai_2 _20942_ (.A1(_10841_),
    .A2(_10844_),
    .B1(_10846_),
    .C1(_10826_),
    .Y(_10848_));
 sky130_fd_sc_hd__nand3b_1 _20943_ (.A_N(_10826_),
    .B(_10845_),
    .C(_10846_),
    .Y(_10850_));
 sky130_fd_sc_hd__a21bo_1 _20944_ (.A1(_10845_),
    .A2(_10846_),
    .B1_N(_10826_),
    .X(_10851_));
 sky130_fd_sc_hd__o21ai_2 _20945_ (.A1(_10724_),
    .A2(_10725_),
    .B1(_10745_),
    .Y(_10852_));
 sky130_fd_sc_hd__nand2_1 _20946_ (.A(_10746_),
    .B(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__nand4_4 _20947_ (.A(_10746_),
    .B(_10850_),
    .C(_10851_),
    .D(_10852_),
    .Y(_10854_));
 sky130_fd_sc_hd__nand3_4 _20948_ (.A(_10853_),
    .B(_10848_),
    .C(_10847_),
    .Y(_10855_));
 sky130_fd_sc_hd__nand2_2 _20949_ (.A(_10854_),
    .B(_10855_),
    .Y(_10856_));
 sky130_fd_sc_hd__and3_1 _20950_ (.A(_10854_),
    .B(_10855_),
    .C(_10825_),
    .X(_10857_));
 sky130_fd_sc_hd__a21oi_1 _20951_ (.A1(_10854_),
    .A2(_10855_),
    .B1(_10825_),
    .Y(_10858_));
 sky130_fd_sc_hd__nand2_2 _20952_ (.A(_10856_),
    .B(_10825_),
    .Y(_10859_));
 sky130_fd_sc_hd__nand3b_4 _20953_ (.A_N(_10825_),
    .B(_10854_),
    .C(_10855_),
    .Y(_10861_));
 sky130_fd_sc_hd__nand2_2 _20954_ (.A(_10859_),
    .B(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__o22a_1 _20955_ (.A1(_10704_),
    .A2(_10711_),
    .B1(_10715_),
    .B2(_10709_),
    .X(_10863_));
 sky130_fd_sc_hd__o21ai_2 _20956_ (.A1(_10715_),
    .A2(_10709_),
    .B1(_10713_),
    .Y(_10864_));
 sky130_fd_sc_hd__nand2_1 _20957_ (.A(_10699_),
    .B(_10705_),
    .Y(_10865_));
 sky130_fd_sc_hd__nor2_1 _20958_ (.A(_04015_),
    .B(_06030_),
    .Y(_10866_));
 sky130_fd_sc_hd__a31oi_2 _20959_ (.A1(_00625_),
    .A2(net250),
    .A3(net274),
    .B1(_10866_),
    .Y(_10867_));
 sky130_fd_sc_hd__a31o_1 _20960_ (.A1(_00625_),
    .A2(net250),
    .A3(net274),
    .B1(_10866_),
    .X(_10868_));
 sky130_fd_sc_hd__nor2_1 _20961_ (.A(_04026_),
    .B(_05766_),
    .Y(_10869_));
 sky130_fd_sc_hd__o311a_1 _20962_ (.A1(net259),
    .A2(_11387_),
    .A3(_02442_),
    .B1(net275),
    .C1(_02421_),
    .X(_10870_));
 sky130_fd_sc_hd__o221ai_4 _20963_ (.A1(_02475_),
    .A2(_05763_),
    .B1(_05766_),
    .B2(_04026_),
    .C1(_10867_),
    .Y(_10872_));
 sky130_fd_sc_hd__o21a_2 _20964_ (.A1(_10869_),
    .A2(_10870_),
    .B1(_10868_),
    .X(_10873_));
 sky130_fd_sc_hd__o21ai_1 _20965_ (.A1(_10869_),
    .A2(_10870_),
    .B1(_10868_),
    .Y(_10874_));
 sky130_fd_sc_hd__a32o_2 _20966_ (.A1(net234),
    .A2(net251),
    .A3(net273),
    .B1(_06326_),
    .B2(net4),
    .X(_10875_));
 sky130_fd_sc_hd__a21oi_1 _20967_ (.A1(_10872_),
    .A2(_10874_),
    .B1(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__a21o_1 _20968_ (.A1(_10872_),
    .A2(_10874_),
    .B1(_10875_),
    .X(_10877_));
 sky130_fd_sc_hd__nand2_1 _20969_ (.A(_10872_),
    .B(_10875_),
    .Y(_10878_));
 sky130_fd_sc_hd__and3_2 _20970_ (.A(_10872_),
    .B(_10874_),
    .C(_10875_),
    .X(_10879_));
 sky130_fd_sc_hd__o22ai_4 _20971_ (.A1(_10481_),
    .A2(_10483_),
    .B1(_10876_),
    .B2(_10879_),
    .Y(_10880_));
 sky130_fd_sc_hd__o211ai_4 _20972_ (.A1(_10873_),
    .A2(_10878_),
    .B1(_10485_),
    .C1(_10877_),
    .Y(_10881_));
 sky130_fd_sc_hd__inv_2 _20973_ (.A(_10881_),
    .Y(_10883_));
 sky130_fd_sc_hd__o21a_1 _20974_ (.A1(_10680_),
    .A2(_10681_),
    .B1(_10689_),
    .X(_10884_));
 sky130_fd_sc_hd__a21oi_1 _20975_ (.A1(_10682_),
    .A2(_10689_),
    .B1(_10690_),
    .Y(_10885_));
 sky130_fd_sc_hd__inv_2 _20976_ (.A(_10885_),
    .Y(_10886_));
 sky130_fd_sc_hd__a21oi_4 _20977_ (.A1(_10880_),
    .A2(_10881_),
    .B1(_10886_),
    .Y(_10887_));
 sky130_fd_sc_hd__a21o_1 _20978_ (.A1(_10880_),
    .A2(_10881_),
    .B1(_10886_),
    .X(_10888_));
 sky130_fd_sc_hd__o21ai_1 _20979_ (.A1(_10690_),
    .A2(_10884_),
    .B1(_10880_),
    .Y(_10889_));
 sky130_fd_sc_hd__o211a_2 _20980_ (.A1(_10690_),
    .A2(_10884_),
    .B1(_10881_),
    .C1(_10880_),
    .X(_10890_));
 sky130_fd_sc_hd__a32oi_4 _20981_ (.A1(_10182_),
    .A2(_10467_),
    .A3(_10469_),
    .B1(_10470_),
    .B2(_10487_),
    .Y(_10891_));
 sky130_fd_sc_hd__o41ai_2 _20982_ (.A1(_10177_),
    .A2(_10180_),
    .A3(_10465_),
    .A4(_10468_),
    .B1(_10491_),
    .Y(_10892_));
 sky130_fd_sc_hd__o21a_1 _20983_ (.A1(_10887_),
    .A2(_10890_),
    .B1(_10891_),
    .X(_10894_));
 sky130_fd_sc_hd__o21ai_4 _20984_ (.A1(_10887_),
    .A2(_10890_),
    .B1(_10891_),
    .Y(_10895_));
 sky130_fd_sc_hd__a32o_1 _20985_ (.A1(_10880_),
    .A2(_10881_),
    .A3(_10886_),
    .B1(_10491_),
    .B2(_10471_),
    .X(_10896_));
 sky130_fd_sc_hd__a211oi_4 _20986_ (.A1(_10471_),
    .A2(_10491_),
    .B1(_10887_),
    .C1(_10890_),
    .Y(_10897_));
 sky130_fd_sc_hd__o211ai_4 _20987_ (.A1(_10889_),
    .A2(_10883_),
    .B1(_10888_),
    .C1(_10892_),
    .Y(_10898_));
 sky130_fd_sc_hd__o22ai_4 _20988_ (.A1(_10700_),
    .A2(_10704_),
    .B1(_10894_),
    .B2(_10897_),
    .Y(_10899_));
 sky130_fd_sc_hd__nand4_4 _20989_ (.A(_10699_),
    .B(_10705_),
    .C(_10895_),
    .D(_10898_),
    .Y(_10900_));
 sky130_fd_sc_hd__a21oi_1 _20990_ (.A1(_10895_),
    .A2(_10898_),
    .B1(_10865_),
    .Y(_10901_));
 sky130_fd_sc_hd__o21bai_2 _20991_ (.A1(_10894_),
    .A2(_10897_),
    .B1_N(_10865_),
    .Y(_10902_));
 sky130_fd_sc_hd__o211ai_4 _20992_ (.A1(_10700_),
    .A2(_10704_),
    .B1(_10895_),
    .C1(_10898_),
    .Y(_10903_));
 sky130_fd_sc_hd__nand2_1 _20993_ (.A(_10864_),
    .B(_10903_),
    .Y(_10905_));
 sky130_fd_sc_hd__a22oi_2 _20994_ (.A1(_10713_),
    .A2(_10717_),
    .B1(_10899_),
    .B2(_10900_),
    .Y(_10906_));
 sky130_fd_sc_hd__nand3_2 _20995_ (.A(_10864_),
    .B(_10902_),
    .C(_10903_),
    .Y(_10907_));
 sky130_fd_sc_hd__a21oi_2 _20996_ (.A1(_10902_),
    .A2(_10903_),
    .B1(_10864_),
    .Y(_10908_));
 sky130_fd_sc_hd__nand3_2 _20997_ (.A(_10899_),
    .B(_10900_),
    .C(_10863_),
    .Y(_10909_));
 sky130_fd_sc_hd__a31oi_2 _20998_ (.A1(_10863_),
    .A2(_10899_),
    .A3(_10900_),
    .B1(_10862_),
    .Y(_10910_));
 sky130_fd_sc_hd__o221a_1 _20999_ (.A1(_10857_),
    .A2(_10858_),
    .B1(_10901_),
    .B2(_10905_),
    .C1(_10909_),
    .X(_10911_));
 sky130_fd_sc_hd__o21ai_2 _21000_ (.A1(_10901_),
    .A2(_10905_),
    .B1(_10910_),
    .Y(_10912_));
 sky130_fd_sc_hd__a22oi_4 _21001_ (.A1(_10859_),
    .A2(_10861_),
    .B1(_10907_),
    .B2(_10909_),
    .Y(_10913_));
 sky130_fd_sc_hd__o2bb2ai_2 _21002_ (.A1_N(_10859_),
    .A2_N(_10861_),
    .B1(_10906_),
    .B2(_10908_),
    .Y(_10914_));
 sky130_fd_sc_hd__and4_1 _21003_ (.A(_10500_),
    .B(_10823_),
    .C(_10912_),
    .D(_10914_),
    .X(_10916_));
 sky130_fd_sc_hd__nand4_4 _21004_ (.A(_10500_),
    .B(_10823_),
    .C(_10912_),
    .D(_10914_),
    .Y(_10917_));
 sky130_fd_sc_hd__o21ai_4 _21005_ (.A1(_10911_),
    .A2(_10913_),
    .B1(_10824_),
    .Y(_10918_));
 sky130_fd_sc_hd__inv_2 _21006_ (.A(_10918_),
    .Y(_10919_));
 sky130_fd_sc_hd__o21ai_2 _21007_ (.A1(_10718_),
    .A2(_10759_),
    .B1(_10721_),
    .Y(_10920_));
 sky130_fd_sc_hd__inv_2 _21008_ (.A(_10920_),
    .Y(_10921_));
 sky130_fd_sc_hd__a21oi_2 _21009_ (.A1(_10917_),
    .A2(_10918_),
    .B1(_10920_),
    .Y(_10922_));
 sky130_fd_sc_hd__a21o_1 _21010_ (.A1(_10917_),
    .A2(_10918_),
    .B1(_10920_),
    .X(_10923_));
 sky130_fd_sc_hd__o21a_1 _21011_ (.A1(_10720_),
    .A2(_10761_),
    .B1(_10918_),
    .X(_10924_));
 sky130_fd_sc_hd__o311a_1 _21012_ (.A1(_10911_),
    .A2(_10913_),
    .A3(_10824_),
    .B1(_10920_),
    .C1(_10918_),
    .X(_10925_));
 sky130_fd_sc_hd__nand2_1 _21013_ (.A(_10924_),
    .B(_10917_),
    .Y(_10927_));
 sky130_fd_sc_hd__o2111a_1 _21014_ (.A1(_10759_),
    .A2(_10718_),
    .B1(_10721_),
    .C1(_10917_),
    .D1(_10918_),
    .X(_10928_));
 sky130_fd_sc_hd__o2111ai_4 _21015_ (.A1(_10759_),
    .A2(_10718_),
    .B1(_10721_),
    .C1(_10917_),
    .D1(_10918_),
    .Y(_10929_));
 sky130_fd_sc_hd__a21oi_1 _21016_ (.A1(_10917_),
    .A2(_10918_),
    .B1(_10921_),
    .Y(_10930_));
 sky130_fd_sc_hd__a21o_1 _21017_ (.A1(_10917_),
    .A2(_10918_),
    .B1(_10921_),
    .X(_10931_));
 sky130_fd_sc_hd__o21a_1 _21018_ (.A1(_10656_),
    .A2(_10657_),
    .B1(_10593_),
    .X(_10932_));
 sky130_fd_sc_hd__a31oi_2 _21019_ (.A1(_10593_),
    .A2(_10652_),
    .A3(_10655_),
    .B1(_10594_),
    .Y(_10933_));
 sky130_fd_sc_hd__a21oi_2 _21020_ (.A1(_10614_),
    .A2(_10626_),
    .B1(_10624_),
    .Y(_10934_));
 sky130_fd_sc_hd__and3_2 _21021_ (.A(_03971_),
    .B(net20),
    .C(net64),
    .X(_10935_));
 sky130_fd_sc_hd__o311a_1 _21022_ (.A1(net246),
    .A2(_05928_),
    .A3(_07074_),
    .B1(net289),
    .C1(_07072_),
    .X(_10936_));
 sky130_fd_sc_hd__a21oi_2 _21023_ (.A1(net289),
    .A2(_07077_),
    .B1(_10935_),
    .Y(_10938_));
 sky130_fd_sc_hd__a31o_1 _21024_ (.A1(_07072_),
    .A2(net168),
    .A3(net289),
    .B1(_10935_),
    .X(_10939_));
 sky130_fd_sc_hd__nor2_1 _21025_ (.A(_04223_),
    .B(_08283_),
    .Y(_10940_));
 sky130_fd_sc_hd__a31oi_4 _21026_ (.A1(_07499_),
    .A2(net167),
    .A3(net291),
    .B1(_10940_),
    .Y(_10941_));
 sky130_fd_sc_hd__o2111ai_4 _21027_ (.A1(net168),
    .A2(_07765_),
    .B1(net63),
    .C1(_07771_),
    .D1(_03927_),
    .Y(_10942_));
 sky130_fd_sc_hd__nor2_1 _21028_ (.A(_04245_),
    .B(_07691_),
    .Y(_10943_));
 sky130_fd_sc_hd__or3_1 _21029_ (.A(net63),
    .B(_04245_),
    .C(_03927_),
    .X(_10944_));
 sky130_fd_sc_hd__a31oi_4 _21030_ (.A1(_07771_),
    .A2(_07658_),
    .A3(net165),
    .B1(_10943_),
    .Y(_10945_));
 sky130_fd_sc_hd__a21oi_1 _21031_ (.A1(_10942_),
    .A2(_10944_),
    .B1(_10941_),
    .Y(_10946_));
 sky130_fd_sc_hd__a21o_2 _21032_ (.A1(_10942_),
    .A2(_10944_),
    .B1(_10941_),
    .X(_10947_));
 sky130_fd_sc_hd__o311a_1 _21033_ (.A1(_03927_),
    .A2(net63),
    .A3(_04245_),
    .B1(_10942_),
    .C1(_10941_),
    .X(_10949_));
 sky130_fd_sc_hd__nand2_2 _21034_ (.A(_10941_),
    .B(_10945_),
    .Y(_10950_));
 sky130_fd_sc_hd__and3_1 _21035_ (.A(_10939_),
    .B(_10947_),
    .C(_10950_),
    .X(_10951_));
 sky130_fd_sc_hd__o211ai_4 _21036_ (.A1(_10935_),
    .A2(_10936_),
    .B1(_10947_),
    .C1(_10950_),
    .Y(_10952_));
 sky130_fd_sc_hd__a21oi_1 _21037_ (.A1(_10947_),
    .A2(_10950_),
    .B1(_10939_),
    .Y(_10953_));
 sky130_fd_sc_hd__o21ai_2 _21038_ (.A1(_10946_),
    .A2(_10949_),
    .B1(_10938_),
    .Y(_10954_));
 sky130_fd_sc_hd__o2bb2ai_2 _21039_ (.A1_N(_10941_),
    .A2_N(_10945_),
    .B1(_10935_),
    .B2(_10936_),
    .Y(_10955_));
 sky130_fd_sc_hd__a21oi_2 _21040_ (.A1(_10939_),
    .A2(_10950_),
    .B1(_10946_),
    .Y(_10956_));
 sky130_fd_sc_hd__o21ai_4 _21041_ (.A1(_10941_),
    .A2(_10945_),
    .B1(_10955_),
    .Y(_10957_));
 sky130_fd_sc_hd__o2111ai_1 _21042_ (.A1(_04245_),
    .A2(_07691_),
    .B1(_10942_),
    .C1(_10941_),
    .D1(_10938_),
    .Y(_10958_));
 sky130_fd_sc_hd__o211ai_2 _21043_ (.A1(_10941_),
    .A2(_10945_),
    .B1(_10955_),
    .C1(_10958_),
    .Y(_10960_));
 sky130_fd_sc_hd__o211a_2 _21044_ (.A1(_10938_),
    .A2(_10947_),
    .B1(_10934_),
    .C1(_10960_),
    .X(_10961_));
 sky130_fd_sc_hd__o211ai_4 _21045_ (.A1(_10938_),
    .A2(_10947_),
    .B1(_10934_),
    .C1(_10960_),
    .Y(_10962_));
 sky130_fd_sc_hd__o211a_4 _21046_ (.A1(_10624_),
    .A2(_10627_),
    .B1(_10952_),
    .C1(_10954_),
    .X(_10963_));
 sky130_fd_sc_hd__o211ai_4 _21047_ (.A1(_10624_),
    .A2(_10627_),
    .B1(_10952_),
    .C1(_10954_),
    .Y(_10964_));
 sky130_fd_sc_hd__nor2_1 _21048_ (.A(_04179_),
    .B(_12363_),
    .Y(_10965_));
 sky130_fd_sc_hd__a31oi_2 _21049_ (.A1(net198),
    .A2(net172),
    .A3(_12330_),
    .B1(_10965_),
    .Y(_10966_));
 sky130_fd_sc_hd__or3_1 _21050_ (.A(net35),
    .B(_04201_),
    .C(_03971_),
    .X(_10967_));
 sky130_fd_sc_hd__o211ai_2 _21051_ (.A1(net174),
    .A2(_06759_),
    .B1(net252),
    .C1(net193),
    .Y(_10968_));
 sky130_fd_sc_hd__o311a_1 _21052_ (.A1(_03971_),
    .A2(net35),
    .A3(_04201_),
    .B1(_10968_),
    .C1(_10966_),
    .X(_10969_));
 sky130_fd_sc_hd__o211ai_2 _21053_ (.A1(_04201_),
    .A2(_11804_),
    .B1(_10968_),
    .C1(_10966_),
    .Y(_10971_));
 sky130_fd_sc_hd__o22a_1 _21054_ (.A1(_04168_),
    .A2(_01326_),
    .B1(_06222_),
    .B2(_01304_),
    .X(_10972_));
 sky130_fd_sc_hd__a32o_1 _21055_ (.A1(net201),
    .A2(net173),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net17),
    .X(_10973_));
 sky130_fd_sc_hd__nand2_1 _21056_ (.A(_10969_),
    .B(_10972_),
    .Y(_10974_));
 sky130_fd_sc_hd__a21oi_1 _21057_ (.A1(_10967_),
    .A2(_10968_),
    .B1(_10966_),
    .Y(_10975_));
 sky130_fd_sc_hd__a21o_1 _21058_ (.A1(_10967_),
    .A2(_10968_),
    .B1(_10966_),
    .X(_10976_));
 sky130_fd_sc_hd__nor2_1 _21059_ (.A(_10973_),
    .B(_10975_),
    .Y(_10977_));
 sky130_fd_sc_hd__a21o_1 _21060_ (.A1(_10971_),
    .A2(_10973_),
    .B1(_10975_),
    .X(_10978_));
 sky130_fd_sc_hd__a21oi_1 _21061_ (.A1(_10971_),
    .A2(_10973_),
    .B1(_10975_),
    .Y(_10979_));
 sky130_fd_sc_hd__and3_1 _21062_ (.A(_10971_),
    .B(_10973_),
    .C(_10976_),
    .X(_10980_));
 sky130_fd_sc_hd__a21oi_2 _21063_ (.A1(_10971_),
    .A2(_10976_),
    .B1(_10973_),
    .Y(_10982_));
 sky130_fd_sc_hd__o2bb2ai_2 _21064_ (.A1_N(_10974_),
    .A2_N(_10979_),
    .B1(_10976_),
    .B2(_10972_),
    .Y(_10983_));
 sky130_fd_sc_hd__o22a_2 _21065_ (.A1(_10961_),
    .A2(_10963_),
    .B1(_10980_),
    .B2(_10982_),
    .X(_10984_));
 sky130_fd_sc_hd__o2bb2ai_4 _21066_ (.A1_N(_10962_),
    .A2_N(_10964_),
    .B1(_10980_),
    .B2(_10982_),
    .Y(_10985_));
 sky130_fd_sc_hd__nand2_4 _21067_ (.A(_10962_),
    .B(_10983_),
    .Y(_10986_));
 sky130_fd_sc_hd__inv_2 _21068_ (.A(_10986_),
    .Y(_10987_));
 sky130_fd_sc_hd__nand3_2 _21069_ (.A(_10962_),
    .B(_10964_),
    .C(_10983_),
    .Y(_10988_));
 sky130_fd_sc_hd__a31oi_2 _21070_ (.A1(_10574_),
    .A2(_10577_),
    .A3(_10300_),
    .B1(_10583_),
    .Y(_10989_));
 sky130_fd_sc_hd__a31o_2 _21071_ (.A1(_10574_),
    .A2(_10577_),
    .A3(_10300_),
    .B1(_10583_),
    .X(_10990_));
 sky130_fd_sc_hd__a22oi_4 _21072_ (.A1(_10985_),
    .A2(_10988_),
    .B1(_10990_),
    .B2(_10579_),
    .Y(_10991_));
 sky130_fd_sc_hd__o2bb2ai_4 _21073_ (.A1_N(_10985_),
    .A2_N(_10988_),
    .B1(_10989_),
    .B2(_10578_),
    .Y(_10993_));
 sky130_fd_sc_hd__o211ai_4 _21074_ (.A1(_10986_),
    .A2(_10963_),
    .B1(_10579_),
    .C1(_10990_),
    .Y(_10994_));
 sky130_fd_sc_hd__o2111a_1 _21075_ (.A1(_10986_),
    .A2(_10963_),
    .B1(_10579_),
    .C1(_10985_),
    .D1(_10990_),
    .X(_10995_));
 sky130_fd_sc_hd__o2111ai_4 _21076_ (.A1(_10986_),
    .A2(_10963_),
    .B1(_10579_),
    .C1(_10985_),
    .D1(_10990_),
    .Y(_10996_));
 sky130_fd_sc_hd__o21a_1 _21077_ (.A1(_10606_),
    .A2(_10608_),
    .B1(_10634_),
    .X(_10997_));
 sky130_fd_sc_hd__a31o_1 _21078_ (.A1(_10607_),
    .A2(_10610_),
    .A3(_10636_),
    .B1(_10633_),
    .X(_10998_));
 sky130_fd_sc_hd__o31a_1 _21079_ (.A1(_10606_),
    .A2(_10608_),
    .A3(_10635_),
    .B1(_10634_),
    .X(_10999_));
 sky130_fd_sc_hd__o22ai_4 _21080_ (.A1(_10633_),
    .A2(_10638_),
    .B1(_10991_),
    .B2(_10995_),
    .Y(_11000_));
 sky130_fd_sc_hd__o211ai_4 _21081_ (.A1(_10635_),
    .A2(_10997_),
    .B1(_10996_),
    .C1(_10993_),
    .Y(_11001_));
 sky130_fd_sc_hd__o2bb2ai_4 _21082_ (.A1_N(_10993_),
    .A2_N(_10996_),
    .B1(_10997_),
    .B2(_10635_),
    .Y(_11002_));
 sky130_fd_sc_hd__o221ai_4 _21083_ (.A1(_10633_),
    .A2(_10638_),
    .B1(_10984_),
    .B2(_10994_),
    .C1(_10993_),
    .Y(_11004_));
 sky130_fd_sc_hd__a32oi_4 _21084_ (.A1(_10579_),
    .A2(_10580_),
    .A3(_10583_),
    .B1(_10551_),
    .B2(_10550_),
    .Y(_11005_));
 sky130_fd_sc_hd__o2bb2ai_4 _21085_ (.A1_N(_10586_),
    .A2_N(_11005_),
    .B1(_10550_),
    .B2(_10551_),
    .Y(_11006_));
 sky130_fd_sc_hd__a22oi_4 _21086_ (.A1(_10549_),
    .A2(_10556_),
    .B1(_11005_),
    .B2(_10586_),
    .Y(_11007_));
 sky130_fd_sc_hd__a32o_1 _21087_ (.A1(_10520_),
    .A2(_10531_),
    .A3(_10533_),
    .B1(_10534_),
    .B2(_10546_),
    .X(_11008_));
 sky130_fd_sc_hd__a32o_2 _21088_ (.A1(_05841_),
    .A2(_05863_),
    .A3(_08657_),
    .B1(_08659_),
    .B2(net29),
    .X(_11009_));
 sky130_fd_sc_hd__a31oi_4 _21089_ (.A1(net162),
    .A2(net33),
    .A3(net319),
    .B1(_11009_),
    .Y(_11010_));
 sky130_fd_sc_hd__and3_1 _21090_ (.A(_11009_),
    .B(net33),
    .C(net319),
    .X(_11011_));
 sky130_fd_sc_hd__nand3_2 _21091_ (.A(_11009_),
    .B(net33),
    .C(net319),
    .Y(_11012_));
 sky130_fd_sc_hd__o22a_2 _21092_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_11009_),
    .B2(_08877_),
    .X(_11013_));
 sky130_fd_sc_hd__o21ai_1 _21093_ (.A1(_11009_),
    .A2(_08877_),
    .B1(_09300_),
    .Y(_11015_));
 sky130_fd_sc_hd__o21ai_4 _21094_ (.A1(_11010_),
    .A2(_11011_),
    .B1(net148),
    .Y(_11016_));
 sky130_fd_sc_hd__o21ai_2 _21095_ (.A1(_11010_),
    .A2(_11011_),
    .B1(_09300_),
    .Y(_11017_));
 sky130_fd_sc_hd__nand3b_2 _21096_ (.A_N(_11010_),
    .B(_11012_),
    .C(net148),
    .Y(_11018_));
 sky130_fd_sc_hd__o211ai_1 _21097_ (.A1(net319),
    .A2(_04331_),
    .B1(_09298_),
    .C1(_10527_),
    .Y(_11019_));
 sky130_fd_sc_hd__o21ai_2 _21098_ (.A1(_10523_),
    .A2(_08877_),
    .B1(_11019_),
    .Y(_11020_));
 sky130_fd_sc_hd__a21boi_1 _21099_ (.A1(_11015_),
    .A2(_11016_),
    .B1_N(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__nand4_4 _21100_ (.A(_10527_),
    .B(_10530_),
    .C(_11017_),
    .D(_11018_),
    .Y(_11022_));
 sky130_fd_sc_hd__o21ai_2 _21101_ (.A1(_10526_),
    .A2(_10529_),
    .B1(_11016_),
    .Y(_11023_));
 sky130_fd_sc_hd__o221a_1 _21102_ (.A1(_10526_),
    .A2(_10529_),
    .B1(_11010_),
    .B2(net147),
    .C1(_11016_),
    .X(_11024_));
 sky130_fd_sc_hd__o221ai_4 _21103_ (.A1(_10526_),
    .A2(_10529_),
    .B1(_11010_),
    .B2(net147),
    .C1(_11016_),
    .Y(_11026_));
 sky130_fd_sc_hd__a22oi_4 _21104_ (.A1(_10541_),
    .A2(net134),
    .B1(_11022_),
    .B2(_11026_),
    .Y(_11027_));
 sky130_fd_sc_hd__a22o_1 _21105_ (.A1(_10541_),
    .A2(net134),
    .B1(_11022_),
    .B2(_11026_),
    .X(_11028_));
 sky130_fd_sc_hd__a311oi_4 _21106_ (.A1(_11017_),
    .A2(_11018_),
    .A3(_11020_),
    .B1(net137),
    .C1(_10540_),
    .Y(_11029_));
 sky130_fd_sc_hd__and3_1 _21107_ (.A(net133),
    .B(_11022_),
    .C(_11026_),
    .X(_11030_));
 sky130_fd_sc_hd__o2111ai_4 _21108_ (.A1(_11013_),
    .A2(_11023_),
    .B1(_11022_),
    .C1(_10541_),
    .D1(net134),
    .Y(_11031_));
 sky130_fd_sc_hd__a221oi_4 _21109_ (.A1(_10534_),
    .A2(_10548_),
    .B1(_11029_),
    .B2(_11026_),
    .C1(_11027_),
    .Y(_11032_));
 sky130_fd_sc_hd__a221o_4 _21110_ (.A1(_10534_),
    .A2(_10548_),
    .B1(_11029_),
    .B2(_11026_),
    .C1(_11027_),
    .X(_11033_));
 sky130_fd_sc_hd__a21boi_4 _21111_ (.A1(_11028_),
    .A2(_11031_),
    .B1_N(_11008_),
    .Y(_11034_));
 sky130_fd_sc_hd__o21ai_4 _21112_ (.A1(_11027_),
    .A2(_11030_),
    .B1(_11008_),
    .Y(_11035_));
 sky130_fd_sc_hd__a21o_1 _21113_ (.A1(_10562_),
    .A2(_10570_),
    .B1(_10571_),
    .X(_11037_));
 sky130_fd_sc_hd__a32o_2 _21114_ (.A1(net164),
    .A2(net162),
    .A3(_06826_),
    .B1(_06848_),
    .B2(net24),
    .X(_11038_));
 sky130_fd_sc_hd__nor2_1 _21115_ (.A(net25),
    .B(_05238_),
    .Y(_11039_));
 sky130_fd_sc_hd__o311a_4 _21116_ (.A1(net22),
    .A2(net24),
    .A3(_07503_),
    .B1(_05227_),
    .C1(net319),
    .X(_11040_));
 sky130_fd_sc_hd__a21oi_4 _21117_ (.A1(_08208_),
    .A2(_11039_),
    .B1(_10566_),
    .Y(_11041_));
 sky130_fd_sc_hd__a31o_4 _21118_ (.A1(net319),
    .A2(net163),
    .A3(_05227_),
    .B1(_10566_),
    .X(_11042_));
 sky130_fd_sc_hd__nor2_2 _21119_ (.A(_04277_),
    .B(_05720_),
    .Y(_11043_));
 sky130_fd_sc_hd__or3b_4 _21120_ (.A(net61),
    .B(_04277_),
    .C_N(net60),
    .X(_11044_));
 sky130_fd_sc_hd__a21oi_2 _21121_ (.A1(net151),
    .A2(net158),
    .B1(_05699_),
    .Y(_11045_));
 sky130_fd_sc_hd__o221ai_4 _21122_ (.A1(_04277_),
    .A2(_05720_),
    .B1(_05699_),
    .B2(_08669_),
    .C1(net142),
    .Y(_11046_));
 sky130_fd_sc_hd__o22a_2 _21123_ (.A1(_10566_),
    .A2(_11040_),
    .B1(_11043_),
    .B2(_11045_),
    .X(_11048_));
 sky130_fd_sc_hd__o22ai_2 _21124_ (.A1(_10566_),
    .A2(_11040_),
    .B1(_11043_),
    .B2(_11045_),
    .Y(_11049_));
 sky130_fd_sc_hd__o31a_4 _21125_ (.A1(_11042_),
    .A2(_11043_),
    .A3(_11045_),
    .B1(_11038_),
    .X(_11050_));
 sky130_fd_sc_hd__nand2_2 _21126_ (.A(_11038_),
    .B(_11046_),
    .Y(_11051_));
 sky130_fd_sc_hd__a21oi_4 _21127_ (.A1(_11046_),
    .A2(_11049_),
    .B1(_11038_),
    .Y(_11052_));
 sky130_fd_sc_hd__a21o_1 _21128_ (.A1(_11046_),
    .A2(_11049_),
    .B1(_11038_),
    .X(_11053_));
 sky130_fd_sc_hd__nand2_1 _21129_ (.A(_11053_),
    .B(net137),
    .Y(_11054_));
 sky130_fd_sc_hd__nor3_4 _21130_ (.A(net134),
    .B(_11050_),
    .C(_11052_),
    .Y(_11055_));
 sky130_fd_sc_hd__o2111ai_4 _21131_ (.A1(_09755_),
    .A2(_10296_),
    .B1(_10539_),
    .C1(_11051_),
    .D1(_11053_),
    .Y(_11056_));
 sky130_fd_sc_hd__o22a_2 _21132_ (.A1(_10297_),
    .A2(_10538_),
    .B1(_11050_),
    .B2(_11052_),
    .X(_11057_));
 sky130_fd_sc_hd__o22ai_4 _21133_ (.A1(_10297_),
    .A2(_10538_),
    .B1(_11050_),
    .B2(_11052_),
    .Y(_11059_));
 sky130_fd_sc_hd__a21o_1 _21134_ (.A1(_11056_),
    .A2(_11059_),
    .B1(_11037_),
    .X(_11060_));
 sky130_fd_sc_hd__o21ai_2 _21135_ (.A1(_10571_),
    .A2(_10575_),
    .B1(_11059_),
    .Y(_11061_));
 sky130_fd_sc_hd__nand4_4 _21136_ (.A(_10572_),
    .B(_10577_),
    .C(_11056_),
    .D(_11059_),
    .Y(_11062_));
 sky130_fd_sc_hd__o22ai_4 _21137_ (.A1(_10571_),
    .A2(_10575_),
    .B1(_11055_),
    .B2(_11057_),
    .Y(_11063_));
 sky130_fd_sc_hd__nand4_4 _21138_ (.A(_11033_),
    .B(_11035_),
    .C(_11062_),
    .D(_11063_),
    .Y(_11064_));
 sky130_fd_sc_hd__o221ai_4 _21139_ (.A1(_11055_),
    .A2(_11061_),
    .B1(_11032_),
    .B2(_11034_),
    .C1(_11060_),
    .Y(_11065_));
 sky130_fd_sc_hd__o211ai_4 _21140_ (.A1(_11032_),
    .A2(_11034_),
    .B1(_11062_),
    .C1(_11063_),
    .Y(_11066_));
 sky130_fd_sc_hd__o2111ai_4 _21141_ (.A1(_11061_),
    .A2(_11055_),
    .B1(_11035_),
    .C1(_11033_),
    .D1(_11060_),
    .Y(_11067_));
 sky130_fd_sc_hd__a21oi_2 _21142_ (.A1(_11066_),
    .A2(_11067_),
    .B1(_11006_),
    .Y(_11068_));
 sky130_fd_sc_hd__nand3_1 _21143_ (.A(_11007_),
    .B(_11064_),
    .C(_11065_),
    .Y(_11070_));
 sky130_fd_sc_hd__a21oi_2 _21144_ (.A1(_11064_),
    .A2(_11065_),
    .B1(_11007_),
    .Y(_11071_));
 sky130_fd_sc_hd__nand3_1 _21145_ (.A(_11006_),
    .B(_11066_),
    .C(_11067_),
    .Y(_11072_));
 sky130_fd_sc_hd__nand4_2 _21146_ (.A(_11000_),
    .B(_11001_),
    .C(_11070_),
    .D(_11072_),
    .Y(_11073_));
 sky130_fd_sc_hd__o2bb2ai_1 _21147_ (.A1_N(_11000_),
    .A2_N(_11001_),
    .B1(_11068_),
    .B2(_11071_),
    .Y(_11074_));
 sky130_fd_sc_hd__nand4_2 _21148_ (.A(_11002_),
    .B(_11004_),
    .C(_11070_),
    .D(_11072_),
    .Y(_11075_));
 sky130_fd_sc_hd__o2bb2ai_2 _21149_ (.A1_N(_11002_),
    .A2_N(_11004_),
    .B1(_11068_),
    .B2(_11071_),
    .Y(_11076_));
 sky130_fd_sc_hd__o211a_4 _21150_ (.A1(_10594_),
    .A2(_10932_),
    .B1(_11075_),
    .C1(_11076_),
    .X(_11077_));
 sky130_fd_sc_hd__o211ai_4 _21151_ (.A1(_10594_),
    .A2(_10932_),
    .B1(_11075_),
    .C1(_11076_),
    .Y(_11078_));
 sky130_fd_sc_hd__nand3_4 _21152_ (.A(_11074_),
    .B(_10933_),
    .C(_11073_),
    .Y(_11079_));
 sky130_fd_sc_hd__a21oi_1 _21153_ (.A1(_10421_),
    .A2(_10430_),
    .B1(_10427_),
    .Y(_11081_));
 sky130_fd_sc_hd__o21ai_1 _21154_ (.A1(_10420_),
    .A2(_10429_),
    .B1(_10428_),
    .Y(_11082_));
 sky130_fd_sc_hd__a21oi_2 _21155_ (.A1(_10597_),
    .A2(_10605_),
    .B1(_10603_),
    .Y(_11083_));
 sky130_fd_sc_hd__a21o_1 _21156_ (.A1(_10597_),
    .A2(_10605_),
    .B1(_10603_),
    .X(_11084_));
 sky130_fd_sc_hd__a32o_1 _21157_ (.A1(net182),
    .A2(net179),
    .A3(net281),
    .B1(_04217_),
    .B2(net14),
    .X(_11085_));
 sky130_fd_sc_hd__a211o_1 _21158_ (.A1(net177),
    .A2(net16),
    .B1(_02869_),
    .C1(net203),
    .X(_11086_));
 sky130_fd_sc_hd__or3b_2 _21159_ (.A(net38),
    .B(_04157_),
    .C_N(net37),
    .X(_11087_));
 sky130_fd_sc_hd__nor2_1 _21160_ (.A(_04146_),
    .B(_03737_),
    .Y(_11088_));
 sky130_fd_sc_hd__a31oi_4 _21161_ (.A1(net178),
    .A2(net177),
    .A3(net285),
    .B1(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__a21oi_4 _21162_ (.A1(_11086_),
    .A2(_11087_),
    .B1(_11089_),
    .Y(_11090_));
 sky130_fd_sc_hd__a21o_1 _21163_ (.A1(_11086_),
    .A2(_11087_),
    .B1(_11089_),
    .X(_11092_));
 sky130_fd_sc_hd__o311a_1 _21164_ (.A1(net37),
    .A2(_04037_),
    .A3(net155),
    .B1(_11087_),
    .C1(_11089_),
    .X(_11093_));
 sky130_fd_sc_hd__o221ai_4 _21165_ (.A1(_04157_),
    .A2(_02891_),
    .B1(net155),
    .B2(_02869_),
    .C1(_11089_),
    .Y(_11094_));
 sky130_fd_sc_hd__o21bai_4 _21166_ (.A1(_11090_),
    .A2(_11093_),
    .B1_N(_11085_),
    .Y(_11095_));
 sky130_fd_sc_hd__nand3_4 _21167_ (.A(_11085_),
    .B(_11092_),
    .C(_11094_),
    .Y(_11096_));
 sky130_fd_sc_hd__inv_2 _21168_ (.A(_11096_),
    .Y(_11097_));
 sky130_fd_sc_hd__nand2_1 _21169_ (.A(_11095_),
    .B(_11096_),
    .Y(_11098_));
 sky130_fd_sc_hd__a21oi_4 _21170_ (.A1(_11095_),
    .A2(_11096_),
    .B1(_11084_),
    .Y(_11099_));
 sky130_fd_sc_hd__a21o_1 _21171_ (.A1(_11095_),
    .A2(_11096_),
    .B1(_11084_),
    .X(_11100_));
 sky130_fd_sc_hd__o211a_4 _21172_ (.A1(_10603_),
    .A2(_10608_),
    .B1(_11095_),
    .C1(_11096_),
    .X(_11101_));
 sky130_fd_sc_hd__o211ai_1 _21173_ (.A1(_10603_),
    .A2(_10608_),
    .B1(_11095_),
    .C1(_11096_),
    .Y(_11103_));
 sky130_fd_sc_hd__o21ai_1 _21174_ (.A1(_11099_),
    .A2(_11101_),
    .B1(_11081_),
    .Y(_11104_));
 sky130_fd_sc_hd__a22oi_4 _21175_ (.A1(_10428_),
    .A2(_10435_),
    .B1(_11098_),
    .B2(_11083_),
    .Y(_11105_));
 sky130_fd_sc_hd__o2bb2ai_1 _21176_ (.A1_N(_11083_),
    .A2_N(_11098_),
    .B1(_10427_),
    .B2(_10434_),
    .Y(_11106_));
 sky130_fd_sc_hd__nand3_2 _21177_ (.A(_11100_),
    .B(_11103_),
    .C(_11081_),
    .Y(_11107_));
 sky130_fd_sc_hd__o22ai_4 _21178_ (.A1(_10427_),
    .A2(_10434_),
    .B1(_11099_),
    .B2(_11101_),
    .Y(_11108_));
 sky130_fd_sc_hd__o2111ai_4 _21179_ (.A1(_10417_),
    .A2(_10437_),
    .B1(_10439_),
    .C1(_11107_),
    .D1(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__inv_2 _21180_ (.A(_11109_),
    .Y(_11110_));
 sky130_fd_sc_hd__a2bb2oi_4 _21181_ (.A1_N(_10438_),
    .A2_N(_10440_),
    .B1(_11107_),
    .B2(_11108_),
    .Y(_11111_));
 sky130_fd_sc_hd__o221ai_4 _21182_ (.A1(_10438_),
    .A2(_10440_),
    .B1(_11101_),
    .B2(_11106_),
    .C1(_11104_),
    .Y(_11112_));
 sky130_fd_sc_hd__a21oi_1 _21183_ (.A1(_10454_),
    .A2(_10464_),
    .B1(_10462_),
    .Y(_11114_));
 sky130_fd_sc_hd__a21o_2 _21184_ (.A1(_10454_),
    .A2(_10464_),
    .B1(_10462_),
    .X(_11115_));
 sky130_fd_sc_hd__o211ai_4 _21185_ (.A1(_04787_),
    .A2(net208),
    .B1(net280),
    .C1(net210),
    .Y(_11116_));
 sky130_fd_sc_hd__or3b_4 _21186_ (.A(net41),
    .B(_04113_),
    .C_N(net40),
    .X(_11117_));
 sky130_fd_sc_hd__o221ai_4 _21187_ (.A1(net231),
    .A2(_04787_),
    .B1(_04091_),
    .B2(net216),
    .C1(net279),
    .Y(_11118_));
 sky130_fd_sc_hd__or3b_2 _21188_ (.A(net42),
    .B(_04091_),
    .C_N(net41),
    .X(_11119_));
 sky130_fd_sc_hd__a22oi_4 _21189_ (.A1(_11116_),
    .A2(_11117_),
    .B1(_11118_),
    .B2(_11119_),
    .Y(_11120_));
 sky130_fd_sc_hd__a22o_1 _21190_ (.A1(_11116_),
    .A2(_11117_),
    .B1(_11118_),
    .B2(_11119_),
    .X(_11121_));
 sky130_fd_sc_hd__o2111a_2 _21191_ (.A1(_04091_),
    .A2(_04483_),
    .B1(_11116_),
    .C1(_11117_),
    .D1(_11118_),
    .X(_11122_));
 sky130_fd_sc_hd__o2111ai_4 _21192_ (.A1(_04091_),
    .A2(_04483_),
    .B1(_11116_),
    .C1(_11117_),
    .D1(_11118_),
    .Y(_11123_));
 sky130_fd_sc_hd__a32o_4 _21193_ (.A1(net218),
    .A2(net186),
    .A3(net243),
    .B1(_04897_),
    .B2(net10),
    .X(_11125_));
 sky130_fd_sc_hd__o21bai_2 _21194_ (.A1(_11120_),
    .A2(_11122_),
    .B1_N(_11125_),
    .Y(_11126_));
 sky130_fd_sc_hd__nand3_1 _21195_ (.A(_11121_),
    .B(_11123_),
    .C(_11125_),
    .Y(_11127_));
 sky130_fd_sc_hd__o21ai_2 _21196_ (.A1(_11120_),
    .A2(_11122_),
    .B1(_11125_),
    .Y(_11128_));
 sky130_fd_sc_hd__nand3b_2 _21197_ (.A_N(_11125_),
    .B(_11123_),
    .C(_11121_),
    .Y(_11129_));
 sky130_fd_sc_hd__nand2_1 _21198_ (.A(_11128_),
    .B(_11129_),
    .Y(_11130_));
 sky130_fd_sc_hd__nand3_4 _21199_ (.A(_11128_),
    .B(_11129_),
    .C(_11114_),
    .Y(_11131_));
 sky130_fd_sc_hd__and3_1 _21200_ (.A(_11115_),
    .B(_11126_),
    .C(_11127_),
    .X(_11132_));
 sky130_fd_sc_hd__nand3_4 _21201_ (.A(_11115_),
    .B(_11126_),
    .C(_11127_),
    .Y(_11133_));
 sky130_fd_sc_hd__o32a_1 _21202_ (.A1(_05463_),
    .A2(_03957_),
    .A3(_03951_),
    .B1(_04048_),
    .B2(_05465_),
    .X(_11134_));
 sky130_fd_sc_hd__a32o_1 _21203_ (.A1(_03952_),
    .A2(net231),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net7),
    .X(_11136_));
 sky130_fd_sc_hd__nand4_4 _21204_ (.A(_04102_),
    .B(net222),
    .C(net45),
    .D(net188),
    .Y(_11137_));
 sky130_fd_sc_hd__or3_2 _21205_ (.A(net45),
    .B(_04102_),
    .C(_04069_),
    .X(_11138_));
 sky130_fd_sc_hd__nor2_1 _21206_ (.A(_04059_),
    .B(_05229_),
    .Y(_11139_));
 sky130_fd_sc_hd__a31oi_4 _21207_ (.A1(net229),
    .A2(net227),
    .A3(net276),
    .B1(_11139_),
    .Y(_11140_));
 sky130_fd_sc_hd__a21oi_2 _21208_ (.A1(_11137_),
    .A2(_11138_),
    .B1(_11140_),
    .Y(_11141_));
 sky130_fd_sc_hd__a21o_1 _21209_ (.A1(_11137_),
    .A2(_11138_),
    .B1(_11140_),
    .X(_11142_));
 sky130_fd_sc_hd__o211ai_1 _21210_ (.A1(_04069_),
    .A2(_04989_),
    .B1(_11137_),
    .C1(_11140_),
    .Y(_11143_));
 sky130_fd_sc_hd__nand4_1 _21211_ (.A(_11134_),
    .B(_11137_),
    .C(_11138_),
    .D(_11140_),
    .Y(_11144_));
 sky130_fd_sc_hd__a31oi_2 _21212_ (.A1(_11137_),
    .A2(_11140_),
    .A3(_11138_),
    .B1(_11134_),
    .Y(_11145_));
 sky130_fd_sc_hd__a21oi_2 _21213_ (.A1(_11136_),
    .A2(_11143_),
    .B1(_11141_),
    .Y(_11147_));
 sky130_fd_sc_hd__o2bb2ai_2 _21214_ (.A1_N(_11144_),
    .A2_N(_11147_),
    .B1(_11134_),
    .B2(_11142_),
    .Y(_11148_));
 sky130_fd_sc_hd__a22oi_1 _21215_ (.A1(_11141_),
    .A2(_11136_),
    .B1(_11147_),
    .B2(_11144_),
    .Y(_11149_));
 sky130_fd_sc_hd__a21oi_1 _21216_ (.A1(_11131_),
    .A2(_11133_),
    .B1(_11148_),
    .Y(_11150_));
 sky130_fd_sc_hd__a21o_1 _21217_ (.A1(_11131_),
    .A2(_11133_),
    .B1(_11148_),
    .X(_11151_));
 sky130_fd_sc_hd__nand2_2 _21218_ (.A(_11131_),
    .B(_11148_),
    .Y(_11152_));
 sky130_fd_sc_hd__and3_1 _21219_ (.A(_11131_),
    .B(_11133_),
    .C(_11148_),
    .X(_11153_));
 sky130_fd_sc_hd__o21a_1 _21220_ (.A1(_11132_),
    .A2(_11152_),
    .B1(_11151_),
    .X(_11154_));
 sky130_fd_sc_hd__o21ai_1 _21221_ (.A1(_11132_),
    .A2(_11152_),
    .B1(_11151_),
    .Y(_11155_));
 sky130_fd_sc_hd__a21o_1 _21222_ (.A1(_11109_),
    .A2(_11112_),
    .B1(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__o211ai_2 _21223_ (.A1(_11150_),
    .A2(_11153_),
    .B1(_11109_),
    .C1(_11112_),
    .Y(_11158_));
 sky130_fd_sc_hd__o2bb2ai_1 _21224_ (.A1_N(_11109_),
    .A2_N(_11112_),
    .B1(_11150_),
    .B2(_11153_),
    .Y(_11159_));
 sky130_fd_sc_hd__nand2_1 _21225_ (.A(_11109_),
    .B(_11154_),
    .Y(_11160_));
 sky130_fd_sc_hd__a31o_1 _21226_ (.A1(_10637_),
    .A2(_10643_),
    .A3(_10639_),
    .B1(_10648_),
    .X(_11161_));
 sky130_fd_sc_hd__nand2_1 _21227_ (.A(_10645_),
    .B(_11161_),
    .Y(_11162_));
 sky130_fd_sc_hd__nand3_4 _21228_ (.A(_11156_),
    .B(_11158_),
    .C(_11162_),
    .Y(_11163_));
 sky130_fd_sc_hd__o2111ai_4 _21229_ (.A1(_11111_),
    .A2(_11160_),
    .B1(_11161_),
    .C1(_11159_),
    .D1(_10645_),
    .Y(_11164_));
 sky130_fd_sc_hd__o21a_1 _21230_ (.A1(_10489_),
    .A2(_10492_),
    .B1(_10451_),
    .X(_11165_));
 sky130_fd_sc_hd__a32o_1 _21231_ (.A1(_10443_),
    .A2(_10445_),
    .A3(_10447_),
    .B1(_10451_),
    .B2(_10494_),
    .X(_11166_));
 sky130_fd_sc_hd__a21oi_1 _21232_ (.A1(_11163_),
    .A2(_11164_),
    .B1(_11166_),
    .Y(_11167_));
 sky130_fd_sc_hd__a22o_1 _21233_ (.A1(_10451_),
    .A2(_10495_),
    .B1(_11163_),
    .B2(_11164_),
    .X(_11169_));
 sky130_fd_sc_hd__and3_1 _21234_ (.A(_11163_),
    .B(_11164_),
    .C(_11166_),
    .X(_11170_));
 sky130_fd_sc_hd__o2111ai_4 _21235_ (.A1(_10494_),
    .A2(_10449_),
    .B1(_10451_),
    .C1(_11163_),
    .D1(_11164_),
    .Y(_11171_));
 sky130_fd_sc_hd__o2bb2a_1 _21236_ (.A1_N(_11163_),
    .A2_N(_11164_),
    .B1(_11165_),
    .B2(_10449_),
    .X(_11172_));
 sky130_fd_sc_hd__a21bo_1 _21237_ (.A1(_11163_),
    .A2(_11164_),
    .B1_N(_11166_),
    .X(_11173_));
 sky130_fd_sc_hd__and3b_1 _21238_ (.A_N(_11166_),
    .B(_11164_),
    .C(_11163_),
    .X(_11174_));
 sky130_fd_sc_hd__nand3b_2 _21239_ (.A_N(_11166_),
    .B(_11164_),
    .C(_11163_),
    .Y(_11175_));
 sky130_fd_sc_hd__nand2_2 _21240_ (.A(_11169_),
    .B(_11171_),
    .Y(_11176_));
 sky130_fd_sc_hd__o2bb2ai_4 _21241_ (.A1_N(_11078_),
    .A2_N(_11079_),
    .B1(_11172_),
    .B2(_11174_),
    .Y(_11177_));
 sky130_fd_sc_hd__nand3_2 _21242_ (.A(_11079_),
    .B(_11173_),
    .C(_11175_),
    .Y(_11178_));
 sky130_fd_sc_hd__nand4_4 _21243_ (.A(_11078_),
    .B(_11079_),
    .C(_11173_),
    .D(_11175_),
    .Y(_11180_));
 sky130_fd_sc_hd__nand4_4 _21244_ (.A(_11078_),
    .B(_11079_),
    .C(_11169_),
    .D(_11171_),
    .Y(_11181_));
 sky130_fd_sc_hd__o2bb2ai_4 _21245_ (.A1_N(_11078_),
    .A2_N(_11079_),
    .B1(_11167_),
    .B2(_11170_),
    .Y(_11182_));
 sky130_fd_sc_hd__a21oi_1 _21246_ (.A1(_10511_),
    .A2(_10665_),
    .B1(_10666_),
    .Y(_11183_));
 sky130_fd_sc_hd__o21bai_4 _21247_ (.A1(_10663_),
    .A2(_10512_),
    .B1_N(_10666_),
    .Y(_11184_));
 sky130_fd_sc_hd__a21oi_4 _21248_ (.A1(_11177_),
    .A2(_11180_),
    .B1(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__o2111ai_4 _21249_ (.A1(_10512_),
    .A2(_10663_),
    .B1(_10667_),
    .C1(_11181_),
    .D1(_11182_),
    .Y(_11186_));
 sky130_fd_sc_hd__o211a_4 _21250_ (.A1(_11178_),
    .A2(_11077_),
    .B1(_11177_),
    .C1(_11184_),
    .X(_11187_));
 sky130_fd_sc_hd__o211ai_4 _21251_ (.A1(_11077_),
    .A2(_11178_),
    .B1(_11184_),
    .C1(_11177_),
    .Y(_11188_));
 sky130_fd_sc_hd__a32oi_4 _21252_ (.A1(_11183_),
    .A2(_11182_),
    .A3(_11181_),
    .B1(_10929_),
    .B2(_10931_),
    .Y(_11189_));
 sky130_fd_sc_hd__o21ai_2 _21253_ (.A1(_10928_),
    .A2(_10930_),
    .B1(_11186_),
    .Y(_11191_));
 sky130_fd_sc_hd__o211a_1 _21254_ (.A1(_10928_),
    .A2(_10930_),
    .B1(_11186_),
    .C1(_11188_),
    .X(_11192_));
 sky130_fd_sc_hd__nand2_1 _21255_ (.A(_11189_),
    .B(_11188_),
    .Y(_11193_));
 sky130_fd_sc_hd__a2bb2oi_2 _21256_ (.A1_N(_10922_),
    .A2_N(_10925_),
    .B1(_11186_),
    .B2(_11188_),
    .Y(_11194_));
 sky130_fd_sc_hd__o22ai_4 _21257_ (.A1(_10922_),
    .A2(_10925_),
    .B1(_11185_),
    .B2(_11187_),
    .Y(_11195_));
 sky130_fd_sc_hd__o21ai_1 _21258_ (.A1(_11187_),
    .A2(_11191_),
    .B1(_11195_),
    .Y(_11196_));
 sky130_fd_sc_hd__a221oi_4 _21259_ (.A1(_11189_),
    .A2(_11188_),
    .B1(_10781_),
    .B2(_10674_),
    .C1(_11194_),
    .Y(_11197_));
 sky130_fd_sc_hd__o211ai_4 _21260_ (.A1(_11187_),
    .A2(_11191_),
    .B1(_11195_),
    .C1(_10822_),
    .Y(_11198_));
 sky130_fd_sc_hd__a21oi_1 _21261_ (.A1(_11193_),
    .A2(_11195_),
    .B1(_10822_),
    .Y(_11199_));
 sky130_fd_sc_hd__o21ai_2 _21262_ (.A1(_11192_),
    .A2(_11194_),
    .B1(_10821_),
    .Y(_11200_));
 sky130_fd_sc_hd__o211a_1 _21263_ (.A1(_10099_),
    .A2(_10059_),
    .B1(_10062_),
    .C1(_10768_),
    .X(_11202_));
 sky130_fd_sc_hd__a21oi_2 _21264_ (.A1(_10767_),
    .A2(_10770_),
    .B1(_10769_),
    .Y(_11203_));
 sky130_fd_sc_hd__o22ai_1 _21265_ (.A1(_10769_),
    .A2(_10777_),
    .B1(_11197_),
    .B2(_11199_),
    .Y(_11204_));
 sky130_fd_sc_hd__o211ai_1 _21266_ (.A1(_10766_),
    .A2(_11202_),
    .B1(_11200_),
    .C1(_11198_),
    .Y(_11205_));
 sky130_fd_sc_hd__o21ai_2 _21267_ (.A1(_11197_),
    .A2(_11199_),
    .B1(_11203_),
    .Y(_11206_));
 sky130_fd_sc_hd__a21oi_2 _21268_ (.A1(_11196_),
    .A2(_10821_),
    .B1(_11203_),
    .Y(_11207_));
 sky130_fd_sc_hd__o211ai_4 _21269_ (.A1(_10769_),
    .A2(_10777_),
    .B1(_11198_),
    .C1(_11200_),
    .Y(_11208_));
 sky130_fd_sc_hd__a22oi_1 _21270_ (.A1(_10789_),
    .A2(_10793_),
    .B1(_11204_),
    .B2(_11205_),
    .Y(_11209_));
 sky130_fd_sc_hd__nand4_4 _21271_ (.A(_10788_),
    .B(_10820_),
    .C(_11206_),
    .D(_11208_),
    .Y(_11210_));
 sky130_fd_sc_hd__a22oi_4 _21272_ (.A1(_10788_),
    .A2(_10820_),
    .B1(_11206_),
    .B2(_11208_),
    .Y(_11211_));
 sky130_fd_sc_hd__nand4_1 _21273_ (.A(_10789_),
    .B(_10793_),
    .C(_11204_),
    .D(_11205_),
    .Y(_11213_));
 sky130_fd_sc_hd__o21ai_1 _21274_ (.A1(_10819_),
    .A2(_11211_),
    .B1(_11210_),
    .Y(_11214_));
 sky130_fd_sc_hd__o22ai_1 _21275_ (.A1(_10753_),
    .A2(_10816_),
    .B1(_11209_),
    .B2(_11211_),
    .Y(_11215_));
 sky130_fd_sc_hd__o211ai_1 _21276_ (.A1(_10755_),
    .A2(_10815_),
    .B1(_11210_),
    .C1(_11213_),
    .Y(_11216_));
 sky130_fd_sc_hd__o22ai_1 _21277_ (.A1(_10755_),
    .A2(_10815_),
    .B1(_11209_),
    .B2(_11211_),
    .Y(_11217_));
 sky130_fd_sc_hd__o211ai_1 _21278_ (.A1(_10753_),
    .A2(_10816_),
    .B1(_11210_),
    .C1(_11213_),
    .Y(_11218_));
 sky130_fd_sc_hd__nand3_1 _21279_ (.A(_10813_),
    .B(_11215_),
    .C(_11216_),
    .Y(_11219_));
 sky130_fd_sc_hd__nand3_1 _21280_ (.A(_10814_),
    .B(_11217_),
    .C(_11218_),
    .Y(_11220_));
 sky130_fd_sc_hd__nand2_1 _21281_ (.A(_11219_),
    .B(_11220_),
    .Y(_11221_));
 sky130_fd_sc_hd__o21a_1 _21282_ (.A1(_10806_),
    .A2(_10812_),
    .B1(_10805_),
    .X(_11222_));
 sky130_fd_sc_hd__xor2_1 _21283_ (.A(_11221_),
    .B(_11222_),
    .X(net95));
 sky130_fd_sc_hd__o21a_1 _21284_ (.A1(_10825_),
    .A2(_10856_),
    .B1(_10855_),
    .X(_11224_));
 sky130_fd_sc_hd__o21ai_1 _21285_ (.A1(_10766_),
    .A2(_11202_),
    .B1(_11198_),
    .Y(_11225_));
 sky130_fd_sc_hd__a32o_1 _21286_ (.A1(_10674_),
    .A2(_10781_),
    .A3(_11196_),
    .B1(_11198_),
    .B2(_11203_),
    .X(_11226_));
 sky130_fd_sc_hd__a32oi_4 _21287_ (.A1(_11177_),
    .A2(_11180_),
    .A3(_11184_),
    .B1(_10927_),
    .B2(_10923_),
    .Y(_11227_));
 sky130_fd_sc_hd__o21ai_2 _21288_ (.A1(_10449_),
    .A2(_11165_),
    .B1(_11164_),
    .Y(_11228_));
 sky130_fd_sc_hd__and3_1 _21289_ (.A(_04266_),
    .B(net54),
    .C(net31),
    .X(_11229_));
 sky130_fd_sc_hd__and3_2 _21290_ (.A(_07242_),
    .B(net257),
    .C(_08005_),
    .X(_11230_));
 sky130_fd_sc_hd__a21oi_2 _21291_ (.A1(net31),
    .A2(_08006_),
    .B1(_11230_),
    .Y(_11231_));
 sky130_fd_sc_hd__a32o_1 _21292_ (.A1(net256),
    .A2(_08700_),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net32),
    .X(_11232_));
 sky130_fd_sc_hd__a21o_1 _21293_ (.A1(_10830_),
    .A2(_10838_),
    .B1(_10839_),
    .X(_11234_));
 sky130_fd_sc_hd__a32o_1 _21294_ (.A1(net255),
    .A2(_09698_),
    .A3(_07305_),
    .B1(_07308_),
    .B2(net2),
    .X(_11235_));
 sky130_fd_sc_hd__nand3_1 _21295_ (.A(net234),
    .B(net251),
    .C(net240),
    .Y(_11236_));
 sky130_fd_sc_hd__or3_1 _21296_ (.A(net51),
    .B(_04190_),
    .C(_04004_),
    .X(_11237_));
 sky130_fd_sc_hd__or3b_1 _21297_ (.A(_03982_),
    .B(net52),
    .C_N(net51),
    .X(_11238_));
 sky130_fd_sc_hd__o211ai_2 _21298_ (.A1(net259),
    .A2(_11387_),
    .B1(net269),
    .C1(_11354_),
    .Y(_11239_));
 sky130_fd_sc_hd__a22oi_1 _21299_ (.A1(_11236_),
    .A2(_11237_),
    .B1(_11238_),
    .B2(_11239_),
    .Y(_11240_));
 sky130_fd_sc_hd__a22o_1 _21300_ (.A1(_11236_),
    .A2(_11237_),
    .B1(_11238_),
    .B2(_11239_),
    .X(_11241_));
 sky130_fd_sc_hd__o2111a_1 _21301_ (.A1(_04004_),
    .A2(_06866_),
    .B1(_11236_),
    .C1(_11238_),
    .D1(_11239_),
    .X(_11242_));
 sky130_fd_sc_hd__o2111ai_1 _21302_ (.A1(_04004_),
    .A2(_06866_),
    .B1(_11236_),
    .C1(_11238_),
    .D1(_11239_),
    .Y(_11243_));
 sky130_fd_sc_hd__o21bai_1 _21303_ (.A1(_11240_),
    .A2(_11242_),
    .B1_N(_11235_),
    .Y(_11245_));
 sky130_fd_sc_hd__nand3_1 _21304_ (.A(_11235_),
    .B(_11241_),
    .C(_11243_),
    .Y(_11246_));
 sky130_fd_sc_hd__a21o_1 _21305_ (.A1(_11245_),
    .A2(_11246_),
    .B1(_11234_),
    .X(_11247_));
 sky130_fd_sc_hd__nand3_2 _21306_ (.A(_11234_),
    .B(_11245_),
    .C(_11246_),
    .Y(_11248_));
 sky130_fd_sc_hd__a21o_1 _21307_ (.A1(_11247_),
    .A2(_11248_),
    .B1(_11232_),
    .X(_11249_));
 sky130_fd_sc_hd__nand3_4 _21308_ (.A(_11232_),
    .B(_11247_),
    .C(_11248_),
    .Y(_11250_));
 sky130_fd_sc_hd__o2bb2ai_4 _21309_ (.A1_N(_10826_),
    .A2_N(_10846_),
    .B1(_10844_),
    .B2(_10841_),
    .Y(_11251_));
 sky130_fd_sc_hd__a21oi_2 _21310_ (.A1(_11249_),
    .A2(_11250_),
    .B1(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__a21o_1 _21311_ (.A1(_11249_),
    .A2(_11250_),
    .B1(_11251_),
    .X(_11253_));
 sky130_fd_sc_hd__and3_1 _21312_ (.A(_11249_),
    .B(_11250_),
    .C(_11251_),
    .X(_11254_));
 sky130_fd_sc_hd__nand3_2 _21313_ (.A(_11249_),
    .B(_11250_),
    .C(_11251_),
    .Y(_11256_));
 sky130_fd_sc_hd__or3_1 _21314_ (.A(_11231_),
    .B(_11252_),
    .C(_11254_),
    .X(_11257_));
 sky130_fd_sc_hd__a211o_1 _21315_ (.A1(_11253_),
    .A2(_11256_),
    .B1(_11229_),
    .C1(_11230_),
    .X(_11258_));
 sky130_fd_sc_hd__o22a_1 _21316_ (.A1(_11229_),
    .A2(_11230_),
    .B1(_11252_),
    .B2(_11254_),
    .X(_11259_));
 sky130_fd_sc_hd__and3_1 _21317_ (.A(_11253_),
    .B(_11256_),
    .C(_11231_),
    .X(_11260_));
 sky130_fd_sc_hd__o2bb2ai_1 _21318_ (.A1_N(_10865_),
    .A2_N(_10895_),
    .B1(_10887_),
    .B2(_10896_),
    .Y(_11261_));
 sky130_fd_sc_hd__a21oi_1 _21319_ (.A1(_10865_),
    .A2(_10895_),
    .B1(_10897_),
    .Y(_11262_));
 sky130_fd_sc_hd__a21o_1 _21320_ (.A1(_10880_),
    .A2(_10886_),
    .B1(_10883_),
    .X(_11263_));
 sky130_fd_sc_hd__nand2_2 _21321_ (.A(_11133_),
    .B(_11149_),
    .Y(_11264_));
 sky130_fd_sc_hd__a21oi_4 _21322_ (.A1(_10872_),
    .A2(_10875_),
    .B1(_10873_),
    .Y(_11265_));
 sky130_fd_sc_hd__o311a_1 _21323_ (.A1(net259),
    .A2(_11387_),
    .A3(_00646_),
    .B1(net273),
    .C1(_00625_),
    .X(_11267_));
 sky130_fd_sc_hd__and3_2 _21324_ (.A(_04190_),
    .B(net49),
    .C(net5),
    .X(_11268_));
 sky130_fd_sc_hd__a31oi_4 _21325_ (.A1(_00625_),
    .A2(net250),
    .A3(net273),
    .B1(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__nand2_1 _21326_ (.A(net248),
    .B(net274),
    .Y(_11270_));
 sky130_fd_sc_hd__o22a_1 _21327_ (.A1(_04026_),
    .A2(_06030_),
    .B1(_02410_),
    .B2(_11270_),
    .X(_11271_));
 sky130_fd_sc_hd__o22ai_4 _21328_ (.A1(_04026_),
    .A2(_06030_),
    .B1(_02410_),
    .B2(_11270_),
    .Y(_11272_));
 sky130_fd_sc_hd__nor2_2 _21329_ (.A(_04048_),
    .B(_05766_),
    .Y(_11273_));
 sky130_fd_sc_hd__a31oi_4 _21330_ (.A1(_03952_),
    .A2(net231),
    .A3(net275),
    .B1(_11273_),
    .Y(_11274_));
 sky130_fd_sc_hd__a31o_1 _21331_ (.A1(_03952_),
    .A2(net231),
    .A3(net275),
    .B1(_11273_),
    .X(_11275_));
 sky130_fd_sc_hd__a211oi_4 _21332_ (.A1(_03959_),
    .A2(net275),
    .B1(_11273_),
    .C1(_11272_),
    .Y(_11276_));
 sky130_fd_sc_hd__a211o_1 _21333_ (.A1(_03959_),
    .A2(net275),
    .B1(_11273_),
    .C1(_11272_),
    .X(_11278_));
 sky130_fd_sc_hd__nor2_2 _21334_ (.A(_11271_),
    .B(_11274_),
    .Y(_11279_));
 sky130_fd_sc_hd__nand2_2 _21335_ (.A(_11272_),
    .B(_11275_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand3_1 _21336_ (.A(_11269_),
    .B(_11271_),
    .C(_11274_),
    .Y(_11281_));
 sky130_fd_sc_hd__o21a_1 _21337_ (.A1(_11271_),
    .A2(_11274_),
    .B1(_11269_),
    .X(_11282_));
 sky130_fd_sc_hd__o22a_1 _21338_ (.A1(_11267_),
    .A2(_11268_),
    .B1(_11272_),
    .B2(_11275_),
    .X(_11283_));
 sky130_fd_sc_hd__o22ai_2 _21339_ (.A1(_11267_),
    .A2(_11268_),
    .B1(_11272_),
    .B2(_11275_),
    .Y(_11284_));
 sky130_fd_sc_hd__o211ai_2 _21340_ (.A1(_11271_),
    .A2(_11274_),
    .B1(_11281_),
    .C1(_11284_),
    .Y(_11285_));
 sky130_fd_sc_hd__o211ai_2 _21341_ (.A1(_11267_),
    .A2(_11268_),
    .B1(_11278_),
    .C1(_11280_),
    .Y(_11286_));
 sky130_fd_sc_hd__o21ai_2 _21342_ (.A1(_11276_),
    .A2(_11279_),
    .B1(_11269_),
    .Y(_11287_));
 sky130_fd_sc_hd__o211ai_4 _21343_ (.A1(_11141_),
    .A2(_11145_),
    .B1(_11286_),
    .C1(_11287_),
    .Y(_11289_));
 sky130_fd_sc_hd__o211ai_4 _21344_ (.A1(_11269_),
    .A2(_11280_),
    .B1(_11285_),
    .C1(_11147_),
    .Y(_11290_));
 sky130_fd_sc_hd__nand2_2 _21345_ (.A(_11289_),
    .B(_11290_),
    .Y(_11291_));
 sky130_fd_sc_hd__o211a_1 _21346_ (.A1(_10873_),
    .A2(_10879_),
    .B1(_11289_),
    .C1(_11290_),
    .X(_11292_));
 sky130_fd_sc_hd__o211ai_4 _21347_ (.A1(_10873_),
    .A2(_10879_),
    .B1(_11289_),
    .C1(_11290_),
    .Y(_11293_));
 sky130_fd_sc_hd__a21boi_1 _21348_ (.A1(_11289_),
    .A2(_11290_),
    .B1_N(_11265_),
    .Y(_11294_));
 sky130_fd_sc_hd__nand2_1 _21349_ (.A(_11291_),
    .B(_11265_),
    .Y(_11295_));
 sky130_fd_sc_hd__a22oi_4 _21350_ (.A1(_11291_),
    .A2(_11265_),
    .B1(_11152_),
    .B2(_11133_),
    .Y(_11296_));
 sky130_fd_sc_hd__o2111ai_4 _21351_ (.A1(_11115_),
    .A2(_11130_),
    .B1(_11264_),
    .C1(_11293_),
    .D1(_11295_),
    .Y(_11297_));
 sky130_fd_sc_hd__o2bb2ai_4 _21352_ (.A1_N(_11131_),
    .A2_N(_11264_),
    .B1(_11292_),
    .B2(_11294_),
    .Y(_11298_));
 sky130_fd_sc_hd__o211a_1 _21353_ (.A1(_10883_),
    .A2(_10890_),
    .B1(_11297_),
    .C1(_11298_),
    .X(_11300_));
 sky130_fd_sc_hd__a21oi_1 _21354_ (.A1(_11297_),
    .A2(_11298_),
    .B1(_11263_),
    .Y(_11301_));
 sky130_fd_sc_hd__a21o_1 _21355_ (.A1(_11297_),
    .A2(_11298_),
    .B1(_11263_),
    .X(_11302_));
 sky130_fd_sc_hd__nand3b_4 _21356_ (.A_N(_11300_),
    .B(_11302_),
    .C(_11261_),
    .Y(_11303_));
 sky130_fd_sc_hd__inv_2 _21357_ (.A(_11303_),
    .Y(_11304_));
 sky130_fd_sc_hd__o21ai_4 _21358_ (.A1(_11300_),
    .A2(_11301_),
    .B1(_11262_),
    .Y(_11305_));
 sky130_fd_sc_hd__o21ai_2 _21359_ (.A1(_11259_),
    .A2(_11260_),
    .B1(_11305_),
    .Y(_11306_));
 sky130_fd_sc_hd__o211a_1 _21360_ (.A1(_11259_),
    .A2(_11260_),
    .B1(_11303_),
    .C1(_11305_),
    .X(_11307_));
 sky130_fd_sc_hd__a22oi_2 _21361_ (.A1(_11257_),
    .A2(_11258_),
    .B1(_11303_),
    .B2(_11305_),
    .Y(_11308_));
 sky130_fd_sc_hd__a22o_1 _21362_ (.A1(_11257_),
    .A2(_11258_),
    .B1(_11303_),
    .B2(_11305_),
    .X(_11309_));
 sky130_fd_sc_hd__o2bb2a_1 _21363_ (.A1_N(_11163_),
    .A2_N(_11228_),
    .B1(_11307_),
    .B2(_11308_),
    .X(_11311_));
 sky130_fd_sc_hd__o2bb2ai_2 _21364_ (.A1_N(_11163_),
    .A2_N(_11228_),
    .B1(_11307_),
    .B2(_11308_),
    .Y(_11312_));
 sky130_fd_sc_hd__o2111ai_4 _21365_ (.A1(_11306_),
    .A2(_11304_),
    .B1(_11228_),
    .C1(_11163_),
    .D1(_11309_),
    .Y(_11313_));
 sky130_fd_sc_hd__a32o_2 _21366_ (.A1(_10863_),
    .A2(_10899_),
    .A3(_10900_),
    .B1(_10907_),
    .B2(_10862_),
    .X(_11314_));
 sky130_fd_sc_hd__o211a_1 _21367_ (.A1(_10906_),
    .A2(_10910_),
    .B1(_11312_),
    .C1(_11313_),
    .X(_11315_));
 sky130_fd_sc_hd__a21boi_2 _21368_ (.A1(_11312_),
    .A2(_11313_),
    .B1_N(_11314_),
    .Y(_11316_));
 sky130_fd_sc_hd__a21oi_1 _21369_ (.A1(_11312_),
    .A2(_11313_),
    .B1(_11314_),
    .Y(_11317_));
 sky130_fd_sc_hd__a2bb2o_1 _21370_ (.A1_N(_10906_),
    .A2_N(_10910_),
    .B1(_11312_),
    .B2(_11313_),
    .X(_11318_));
 sky130_fd_sc_hd__and3_1 _21371_ (.A(_11312_),
    .B(_11313_),
    .C(_11314_),
    .X(_11319_));
 sky130_fd_sc_hd__o2111ai_2 _21372_ (.A1(_10862_),
    .A2(_10908_),
    .B1(_11312_),
    .C1(_11313_),
    .D1(_10907_),
    .Y(_11320_));
 sky130_fd_sc_hd__nand2_1 _21373_ (.A(_11318_),
    .B(_11320_),
    .Y(_11322_));
 sky130_fd_sc_hd__o21ai_2 _21374_ (.A1(_11077_),
    .A2(_11176_),
    .B1(_11079_),
    .Y(_11323_));
 sky130_fd_sc_hd__nand2_1 _21375_ (.A(_11078_),
    .B(_11178_),
    .Y(_11324_));
 sky130_fd_sc_hd__nor2_1 _21376_ (.A(_11125_),
    .B(_11120_),
    .Y(_11325_));
 sky130_fd_sc_hd__a22oi_4 _21377_ (.A1(_04792_),
    .A2(net243),
    .B1(_04897_),
    .B2(net11),
    .Y(_11326_));
 sky130_fd_sc_hd__a32o_1 _21378_ (.A1(net184),
    .A2(net214),
    .A3(net243),
    .B1(_04897_),
    .B2(net11),
    .X(_11327_));
 sky130_fd_sc_hd__a41oi_4 _21379_ (.A1(_06519_),
    .A2(_03955_),
    .A3(net277),
    .A4(_04113_),
    .B1(_04481_),
    .Y(_11328_));
 sky130_fd_sc_hd__o21ai_2 _21380_ (.A1(_04113_),
    .A2(_04788_),
    .B1(_11328_),
    .Y(_11329_));
 sky130_fd_sc_hd__or3b_2 _21381_ (.A(net42),
    .B(_04113_),
    .C_N(net41),
    .X(_11330_));
 sky130_fd_sc_hd__a22oi_2 _21382_ (.A1(net13),
    .A2(_04482_),
    .B1(_11328_),
    .B2(net210),
    .Y(_11331_));
 sky130_fd_sc_hd__nand3_4 _21383_ (.A(net182),
    .B(net179),
    .C(_04267_),
    .Y(_11333_));
 sky130_fd_sc_hd__or3b_2 _21384_ (.A(net41),
    .B(_04135_),
    .C_N(net40),
    .X(_11334_));
 sky130_fd_sc_hd__a22oi_4 _21385_ (.A1(_11329_),
    .A2(_11330_),
    .B1(_11333_),
    .B2(_11334_),
    .Y(_11335_));
 sky130_fd_sc_hd__a22o_1 _21386_ (.A1(_11329_),
    .A2(_11330_),
    .B1(_11333_),
    .B2(_11334_),
    .X(_11336_));
 sky130_fd_sc_hd__o211a_1 _21387_ (.A1(_04135_),
    .A2(_04270_),
    .B1(_11333_),
    .C1(_11331_),
    .X(_11337_));
 sky130_fd_sc_hd__o211ai_4 _21388_ (.A1(_04135_),
    .A2(_04270_),
    .B1(_11333_),
    .C1(_11331_),
    .Y(_11338_));
 sky130_fd_sc_hd__nor3_4 _21389_ (.A(_11326_),
    .B(_11335_),
    .C(_11337_),
    .Y(_11339_));
 sky130_fd_sc_hd__nand3_2 _21390_ (.A(_11327_),
    .B(_11336_),
    .C(_11338_),
    .Y(_11340_));
 sky130_fd_sc_hd__a21oi_1 _21391_ (.A1(_11336_),
    .A2(_11338_),
    .B1(_11327_),
    .Y(_11341_));
 sky130_fd_sc_hd__o21ai_4 _21392_ (.A1(_11335_),
    .A2(_11337_),
    .B1(_11326_),
    .Y(_11342_));
 sky130_fd_sc_hd__o211ai_4 _21393_ (.A1(_11125_),
    .A2(_11120_),
    .B1(_11123_),
    .C1(_11342_),
    .Y(_11344_));
 sky130_fd_sc_hd__o2111ai_4 _21394_ (.A1(_11125_),
    .A2(_11120_),
    .B1(_11123_),
    .C1(_11340_),
    .D1(_11342_),
    .Y(_11345_));
 sky130_fd_sc_hd__a2bb2oi_2 _21395_ (.A1_N(_11122_),
    .A2_N(_11325_),
    .B1(_11340_),
    .B2(_11342_),
    .Y(_11346_));
 sky130_fd_sc_hd__o22ai_4 _21396_ (.A1(_11122_),
    .A2(_11325_),
    .B1(_11339_),
    .B2(_11341_),
    .Y(_11347_));
 sky130_fd_sc_hd__nor2_2 _21397_ (.A(_04059_),
    .B(_05465_),
    .Y(_11348_));
 sky130_fd_sc_hd__and3_1 _21398_ (.A(net229),
    .B(net227),
    .C(_05462_),
    .X(_11349_));
 sky130_fd_sc_hd__a31oi_2 _21399_ (.A1(net229),
    .A2(net227),
    .A3(_05462_),
    .B1(_11348_),
    .Y(_11350_));
 sky130_fd_sc_hd__o31a_1 _21400_ (.A1(net259),
    .A2(_03956_),
    .A3(_04407_),
    .B1(net276),
    .X(_11351_));
 sky130_fd_sc_hd__a22oi_4 _21401_ (.A1(net9),
    .A2(_05228_),
    .B1(_11351_),
    .B2(net221),
    .Y(_11352_));
 sky130_fd_sc_hd__o2111ai_4 _21402_ (.A1(net231),
    .A2(_04557_),
    .B1(net45),
    .C1(net218),
    .D1(_04102_),
    .Y(_11353_));
 sky130_fd_sc_hd__and3_1 _21403_ (.A(_04124_),
    .B(net43),
    .C(net10),
    .X(_11355_));
 sky130_fd_sc_hd__or3_2 _21404_ (.A(net45),
    .B(_04102_),
    .C(_04080_),
    .X(_11356_));
 sky130_fd_sc_hd__a31oi_2 _21405_ (.A1(net218),
    .A2(net186),
    .A3(net242),
    .B1(_11355_),
    .Y(_11357_));
 sky130_fd_sc_hd__a21oi_4 _21406_ (.A1(_11353_),
    .A2(_11356_),
    .B1(_11352_),
    .Y(_11358_));
 sky130_fd_sc_hd__a21o_1 _21407_ (.A1(_11353_),
    .A2(_11356_),
    .B1(_11352_),
    .X(_11359_));
 sky130_fd_sc_hd__o21ai_1 _21408_ (.A1(_04562_),
    .A2(_04986_),
    .B1(_11352_),
    .Y(_11360_));
 sky130_fd_sc_hd__o311a_2 _21409_ (.A1(_04080_),
    .A2(_04102_),
    .A3(net45),
    .B1(_11353_),
    .C1(_11352_),
    .X(_11361_));
 sky130_fd_sc_hd__o21ai_2 _21410_ (.A1(_11358_),
    .A2(_11361_),
    .B1(_11350_),
    .Y(_11362_));
 sky130_fd_sc_hd__o221ai_4 _21411_ (.A1(_11348_),
    .A2(_11349_),
    .B1(_11355_),
    .B2(_11360_),
    .C1(_11359_),
    .Y(_11363_));
 sky130_fd_sc_hd__nor4_2 _21412_ (.A(_11348_),
    .B(_11349_),
    .C(_11358_),
    .D(_11361_),
    .Y(_11364_));
 sky130_fd_sc_hd__o22a_1 _21413_ (.A1(_11348_),
    .A2(_11349_),
    .B1(_11358_),
    .B2(_11361_),
    .X(_11366_));
 sky130_fd_sc_hd__nand2_1 _21414_ (.A(_11362_),
    .B(_11363_),
    .Y(_11367_));
 sky130_fd_sc_hd__a22oi_4 _21415_ (.A1(_11345_),
    .A2(_11347_),
    .B1(_11362_),
    .B2(_11363_),
    .Y(_11368_));
 sky130_fd_sc_hd__a22o_2 _21416_ (.A1(_11345_),
    .A2(_11347_),
    .B1(_11362_),
    .B2(_11363_),
    .X(_11369_));
 sky130_fd_sc_hd__o221a_2 _21417_ (.A1(_11364_),
    .A2(_11366_),
    .B1(_11339_),
    .B2(_11344_),
    .C1(_11347_),
    .X(_11370_));
 sky130_fd_sc_hd__o211ai_4 _21418_ (.A1(_11364_),
    .A2(_11366_),
    .B1(_11345_),
    .C1(_11347_),
    .Y(_11371_));
 sky130_fd_sc_hd__nand2_1 _21419_ (.A(_11369_),
    .B(_11371_),
    .Y(_11372_));
 sky130_fd_sc_hd__a31oi_2 _21420_ (.A1(_11084_),
    .A2(_11095_),
    .A3(_11096_),
    .B1(_11082_),
    .Y(_11373_));
 sky130_fd_sc_hd__a21o_1 _21421_ (.A1(_11085_),
    .A2(_11094_),
    .B1(_11090_),
    .X(_11374_));
 sky130_fd_sc_hd__o311a_1 _21422_ (.A1(net231),
    .A2(_04787_),
    .A3(_05551_),
    .B1(net178),
    .C1(net281),
    .X(_11375_));
 sky130_fd_sc_hd__nor2_1 _21423_ (.A(_04146_),
    .B(_04218_),
    .Y(_11377_));
 sky130_fd_sc_hd__a31o_1 _21424_ (.A1(net178),
    .A2(net177),
    .A3(net281),
    .B1(_11377_),
    .X(_11378_));
 sky130_fd_sc_hd__o211ai_4 _21425_ (.A1(_05927_),
    .A2(_06220_),
    .B1(_02858_),
    .C1(net201),
    .Y(_11379_));
 sky130_fd_sc_hd__or3b_2 _21426_ (.A(net38),
    .B(_04168_),
    .C_N(net37),
    .X(_11380_));
 sky130_fd_sc_hd__nor2_1 _21427_ (.A(_04157_),
    .B(_03737_),
    .Y(_11381_));
 sky130_fd_sc_hd__a221oi_2 _21428_ (.A1(_03957_),
    .A2(_05926_),
    .B1(net177),
    .B2(net16),
    .C1(_03714_),
    .Y(_11382_));
 sky130_fd_sc_hd__o221ai_4 _21429_ (.A1(net231),
    .A2(_05927_),
    .B1(_04157_),
    .B2(net206),
    .C1(net285),
    .Y(_11383_));
 sky130_fd_sc_hd__o2111ai_4 _21430_ (.A1(_04157_),
    .A2(_03737_),
    .B1(_11379_),
    .C1(_11380_),
    .D1(_11383_),
    .Y(_11384_));
 sky130_fd_sc_hd__o2bb2a_2 _21431_ (.A1_N(_11379_),
    .A2_N(_11380_),
    .B1(_11381_),
    .B2(_11382_),
    .X(_11385_));
 sky130_fd_sc_hd__o2bb2ai_2 _21432_ (.A1_N(_11379_),
    .A2_N(_11380_),
    .B1(_11381_),
    .B2(_11382_),
    .Y(_11386_));
 sky130_fd_sc_hd__o211a_4 _21433_ (.A1(_11375_),
    .A2(_11377_),
    .B1(_11384_),
    .C1(_11386_),
    .X(_11388_));
 sky130_fd_sc_hd__a21oi_2 _21434_ (.A1(_11384_),
    .A2(_11386_),
    .B1(_11378_),
    .Y(_11389_));
 sky130_fd_sc_hd__a21o_1 _21435_ (.A1(_11384_),
    .A2(_11386_),
    .B1(_11378_),
    .X(_11390_));
 sky130_fd_sc_hd__nand2_1 _21436_ (.A(_11390_),
    .B(_10978_),
    .Y(_11391_));
 sky130_fd_sc_hd__nor3_2 _21437_ (.A(_10979_),
    .B(_11388_),
    .C(_11389_),
    .Y(_11392_));
 sky130_fd_sc_hd__nand3b_4 _21438_ (.A_N(_11388_),
    .B(_11390_),
    .C(_10978_),
    .Y(_11393_));
 sky130_fd_sc_hd__o22a_1 _21439_ (.A1(_10969_),
    .A2(_10977_),
    .B1(_11388_),
    .B2(_11389_),
    .X(_11394_));
 sky130_fd_sc_hd__o22ai_4 _21440_ (.A1(_10969_),
    .A2(_10977_),
    .B1(_11388_),
    .B2(_11389_),
    .Y(_11395_));
 sky130_fd_sc_hd__nand2_2 _21441_ (.A(_11374_),
    .B(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__a21o_1 _21442_ (.A1(_11393_),
    .A2(_11395_),
    .B1(_11374_),
    .X(_11397_));
 sky130_fd_sc_hd__nand4_4 _21443_ (.A(_11092_),
    .B(_11096_),
    .C(_11393_),
    .D(_11395_),
    .Y(_11399_));
 sky130_fd_sc_hd__o22ai_4 _21444_ (.A1(_11090_),
    .A2(_11097_),
    .B1(_11392_),
    .B2(_11394_),
    .Y(_11400_));
 sky130_fd_sc_hd__a2bb2oi_2 _21445_ (.A1_N(_11101_),
    .A2_N(_11105_),
    .B1(_11399_),
    .B2(_11400_),
    .Y(_11401_));
 sky130_fd_sc_hd__o221ai_4 _21446_ (.A1(_11392_),
    .A2(_11396_),
    .B1(_11101_),
    .B2(_11105_),
    .C1(_11397_),
    .Y(_11402_));
 sky130_fd_sc_hd__o211a_2 _21447_ (.A1(_11099_),
    .A2(_11373_),
    .B1(_11399_),
    .C1(_11400_),
    .X(_11403_));
 sky130_fd_sc_hd__o211ai_4 _21448_ (.A1(_11099_),
    .A2(_11373_),
    .B1(_11399_),
    .C1(_11400_),
    .Y(_11404_));
 sky130_fd_sc_hd__a21o_1 _21449_ (.A1(_11402_),
    .A2(_11404_),
    .B1(_11372_),
    .X(_11405_));
 sky130_fd_sc_hd__o211ai_4 _21450_ (.A1(_11368_),
    .A2(_11370_),
    .B1(_11402_),
    .C1(_11404_),
    .Y(_11406_));
 sky130_fd_sc_hd__o22ai_4 _21451_ (.A1(_11368_),
    .A2(_11370_),
    .B1(_11401_),
    .B2(_11403_),
    .Y(_11407_));
 sky130_fd_sc_hd__nand4_4 _21452_ (.A(_11369_),
    .B(_11371_),
    .C(_11402_),
    .D(_11404_),
    .Y(_11408_));
 sky130_fd_sc_hd__o21ai_2 _21453_ (.A1(_10633_),
    .A2(_10638_),
    .B1(_10993_),
    .Y(_11410_));
 sky130_fd_sc_hd__o22ai_4 _21454_ (.A1(_10984_),
    .A2(_10994_),
    .B1(_10999_),
    .B2(_10991_),
    .Y(_11411_));
 sky130_fd_sc_hd__a21oi_1 _21455_ (.A1(_10993_),
    .A2(_10998_),
    .B1(_10995_),
    .Y(_11412_));
 sky130_fd_sc_hd__a21oi_2 _21456_ (.A1(_11407_),
    .A2(_11408_),
    .B1(_11411_),
    .Y(_11413_));
 sky130_fd_sc_hd__nand3_2 _21457_ (.A(_11405_),
    .B(_11406_),
    .C(_11412_),
    .Y(_11414_));
 sky130_fd_sc_hd__and3_1 _21458_ (.A(_11407_),
    .B(_11411_),
    .C(_11408_),
    .X(_11415_));
 sky130_fd_sc_hd__nand3_4 _21459_ (.A(_11407_),
    .B(_11411_),
    .C(_11408_),
    .Y(_11416_));
 sky130_fd_sc_hd__o21a_1 _21460_ (.A1(_11150_),
    .A2(_11153_),
    .B1(_11112_),
    .X(_11417_));
 sky130_fd_sc_hd__a21o_1 _21461_ (.A1(_11109_),
    .A2(_11154_),
    .B1(_11111_),
    .X(_11418_));
 sky130_fd_sc_hd__a21oi_4 _21462_ (.A1(_11109_),
    .A2(_11154_),
    .B1(_11111_),
    .Y(_11419_));
 sky130_fd_sc_hd__nand3_4 _21463_ (.A(_11414_),
    .B(_11416_),
    .C(_11418_),
    .Y(_11421_));
 sky130_fd_sc_hd__o2bb2ai_4 _21464_ (.A1_N(_11414_),
    .A2_N(_11416_),
    .B1(_11417_),
    .B2(_11110_),
    .Y(_11422_));
 sky130_fd_sc_hd__nand2_1 _21465_ (.A(_11421_),
    .B(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__a32oi_4 _21466_ (.A1(_11006_),
    .A2(_11066_),
    .A3(_11067_),
    .B1(_11004_),
    .B2(_11002_),
    .Y(_11424_));
 sky130_fd_sc_hd__a32oi_4 _21467_ (.A1(_11007_),
    .A2(_11064_),
    .A3(_11065_),
    .B1(_11001_),
    .B2(_11000_),
    .Y(_11425_));
 sky130_fd_sc_hd__and3_1 _21468_ (.A(_03971_),
    .B(net21),
    .C(net64),
    .X(_11426_));
 sky130_fd_sc_hd__o311a_1 _21469_ (.A1(net246),
    .A2(_05928_),
    .A3(_07501_),
    .B1(net289),
    .C1(_07499_),
    .X(_11427_));
 sky130_fd_sc_hd__a31o_1 _21470_ (.A1(_07499_),
    .A2(net167),
    .A3(net289),
    .B1(_11426_),
    .X(_11428_));
 sky130_fd_sc_hd__o211ai_4 _21471_ (.A1(net168),
    .A2(_07765_),
    .B1(net291),
    .C1(_07771_),
    .Y(_11429_));
 sky130_fd_sc_hd__nor2_1 _21472_ (.A(_04245_),
    .B(_08283_),
    .Y(_11430_));
 sky130_fd_sc_hd__or3b_2 _21473_ (.A(net64),
    .B(_04245_),
    .C_N(net63),
    .X(_11432_));
 sky130_fd_sc_hd__a31oi_4 _21474_ (.A1(_07771_),
    .A2(net291),
    .A3(net165),
    .B1(_11430_),
    .Y(_11433_));
 sky130_fd_sc_hd__nor2_1 _21475_ (.A(_04256_),
    .B(_07691_),
    .Y(_11434_));
 sky130_fd_sc_hd__or3_1 _21476_ (.A(net63),
    .B(_04256_),
    .C(_03927_),
    .X(_11435_));
 sky130_fd_sc_hd__a211oi_1 _21477_ (.A1(_07075_),
    .A2(_08205_),
    .B1(_07669_),
    .C1(_08203_),
    .Y(_11436_));
 sky130_fd_sc_hd__a31oi_4 _21478_ (.A1(net164),
    .A2(net162),
    .A3(_07658_),
    .B1(_11434_),
    .Y(_11437_));
 sky130_fd_sc_hd__o311a_2 _21479_ (.A1(_07669_),
    .A2(_08203_),
    .A3(net154),
    .B1(_11435_),
    .C1(_11433_),
    .X(_11438_));
 sky130_fd_sc_hd__nand2_1 _21480_ (.A(_11433_),
    .B(_11437_),
    .Y(_11439_));
 sky130_fd_sc_hd__a21oi_4 _21481_ (.A1(_11429_),
    .A2(_11432_),
    .B1(_11437_),
    .Y(_11440_));
 sky130_fd_sc_hd__o2bb2ai_1 _21482_ (.A1_N(_11429_),
    .A2_N(_11432_),
    .B1(_11434_),
    .B2(_11436_),
    .Y(_11441_));
 sky130_fd_sc_hd__o22ai_4 _21483_ (.A1(_11426_),
    .A2(_11427_),
    .B1(_11433_),
    .B2(_11437_),
    .Y(_11443_));
 sky130_fd_sc_hd__a21oi_4 _21484_ (.A1(_11433_),
    .A2(_11437_),
    .B1(_11443_),
    .Y(_11444_));
 sky130_fd_sc_hd__a31o_1 _21485_ (.A1(_11429_),
    .A2(_11432_),
    .A3(_11437_),
    .B1(_11443_),
    .X(_11445_));
 sky130_fd_sc_hd__a21oi_2 _21486_ (.A1(_11439_),
    .A2(_11441_),
    .B1(_11428_),
    .Y(_11446_));
 sky130_fd_sc_hd__o21bai_4 _21487_ (.A1(_11438_),
    .A2(_11440_),
    .B1_N(_11428_),
    .Y(_11447_));
 sky130_fd_sc_hd__o211ai_4 _21488_ (.A1(_11443_),
    .A2(_11438_),
    .B1(_10957_),
    .C1(_11447_),
    .Y(_11448_));
 sky130_fd_sc_hd__inv_2 _21489_ (.A(_11448_),
    .Y(_11449_));
 sky130_fd_sc_hd__a21oi_4 _21490_ (.A1(_11445_),
    .A2(_11447_),
    .B1(_10957_),
    .Y(_11450_));
 sky130_fd_sc_hd__o21ai_4 _21491_ (.A1(_11444_),
    .A2(_11446_),
    .B1(_10956_),
    .Y(_11451_));
 sky130_fd_sc_hd__o211ai_4 _21492_ (.A1(net174),
    .A2(_06759_),
    .B1(_12330_),
    .C1(net193),
    .Y(_11452_));
 sky130_fd_sc_hd__or3_2 _21493_ (.A(net36),
    .B(_04201_),
    .C(_03993_),
    .X(_11454_));
 sky130_fd_sc_hd__a32oi_2 _21494_ (.A1(net194),
    .A2(net171),
    .A3(_12330_),
    .B1(_12352_),
    .B2(net19),
    .Y(_11455_));
 sky130_fd_sc_hd__and3_1 _21495_ (.A(_03993_),
    .B(net20),
    .C(net34),
    .X(_11456_));
 sky130_fd_sc_hd__a221oi_1 _21496_ (.A1(net203),
    .A2(net272),
    .B1(net171),
    .B2(net20),
    .C1(_11782_),
    .Y(_11457_));
 sky130_fd_sc_hd__a31oi_4 _21497_ (.A1(_07072_),
    .A2(net168),
    .A3(net252),
    .B1(_11456_),
    .Y(_11458_));
 sky130_fd_sc_hd__nand2_1 _21498_ (.A(_11455_),
    .B(_11458_),
    .Y(_11459_));
 sky130_fd_sc_hd__a32oi_4 _21499_ (.A1(net198),
    .A2(net172),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net18),
    .Y(_11460_));
 sky130_fd_sc_hd__a32o_1 _21500_ (.A1(net198),
    .A2(net172),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net18),
    .X(_11461_));
 sky130_fd_sc_hd__a21oi_2 _21501_ (.A1(_11452_),
    .A2(_11454_),
    .B1(_11458_),
    .Y(_11462_));
 sky130_fd_sc_hd__o2bb2ai_2 _21502_ (.A1_N(_11452_),
    .A2_N(_11454_),
    .B1(_11456_),
    .B2(_11457_),
    .Y(_11463_));
 sky130_fd_sc_hd__a21oi_1 _21503_ (.A1(_11455_),
    .A2(_11458_),
    .B1(_11460_),
    .Y(_11465_));
 sky130_fd_sc_hd__a32oi_4 _21504_ (.A1(_11452_),
    .A2(_11454_),
    .A3(_11458_),
    .B1(_11463_),
    .B2(_11460_),
    .Y(_11466_));
 sky130_fd_sc_hd__a21oi_1 _21505_ (.A1(_11459_),
    .A2(_11461_),
    .B1(_11462_),
    .Y(_11467_));
 sky130_fd_sc_hd__o21a_1 _21506_ (.A1(_11459_),
    .A2(_11461_),
    .B1(_11467_),
    .X(_11468_));
 sky130_fd_sc_hd__nor2_1 _21507_ (.A(_11460_),
    .B(_11463_),
    .Y(_11469_));
 sky130_fd_sc_hd__and3_1 _21508_ (.A(_11459_),
    .B(_11461_),
    .C(_11463_),
    .X(_11470_));
 sky130_fd_sc_hd__a21oi_2 _21509_ (.A1(_11459_),
    .A2(_11463_),
    .B1(_11461_),
    .Y(_11471_));
 sky130_fd_sc_hd__a21oi_1 _21510_ (.A1(_11461_),
    .A2(_11462_),
    .B1(_11468_),
    .Y(_11472_));
 sky130_fd_sc_hd__o2bb2ai_2 _21511_ (.A1_N(_11448_),
    .A2_N(_11451_),
    .B1(_11470_),
    .B2(_11471_),
    .Y(_11473_));
 sky130_fd_sc_hd__o21a_1 _21512_ (.A1(_11468_),
    .A2(_11469_),
    .B1(_11451_),
    .X(_11474_));
 sky130_fd_sc_hd__o211ai_2 _21513_ (.A1(_11468_),
    .A2(_11469_),
    .B1(_11448_),
    .C1(_11451_),
    .Y(_11476_));
 sky130_fd_sc_hd__o211ai_2 _21514_ (.A1(_11470_),
    .A2(_11471_),
    .B1(_11448_),
    .C1(_11451_),
    .Y(_11477_));
 sky130_fd_sc_hd__o2bb2ai_1 _21515_ (.A1_N(_11448_),
    .A2_N(_11451_),
    .B1(_11468_),
    .B2(_11469_),
    .Y(_11478_));
 sky130_fd_sc_hd__a31oi_4 _21516_ (.A1(_11053_),
    .A2(net137),
    .A3(_11051_),
    .B1(_11037_),
    .Y(_11479_));
 sky130_fd_sc_hd__o2bb2ai_2 _21517_ (.A1_N(_11037_),
    .A2_N(_11059_),
    .B1(_11050_),
    .B2(_11054_),
    .Y(_11480_));
 sky130_fd_sc_hd__o211ai_4 _21518_ (.A1(_11057_),
    .A2(_11479_),
    .B1(_11478_),
    .C1(_11477_),
    .Y(_11481_));
 sky130_fd_sc_hd__and3_1 _21519_ (.A(_11480_),
    .B(_11476_),
    .C(_11473_),
    .X(_11482_));
 sky130_fd_sc_hd__nand3_4 _21520_ (.A(_11480_),
    .B(_11476_),
    .C(_11473_),
    .Y(_11483_));
 sky130_fd_sc_hd__o32a_2 _21521_ (.A1(_10934_),
    .A2(_10951_),
    .A3(_10953_),
    .B1(_10980_),
    .B2(_10982_),
    .X(_11484_));
 sky130_fd_sc_hd__o31a_1 _21522_ (.A1(_10934_),
    .A2(_10951_),
    .A3(_10953_),
    .B1(_10986_),
    .X(_11485_));
 sky130_fd_sc_hd__o2bb2ai_2 _21523_ (.A1_N(_11481_),
    .A2_N(_11483_),
    .B1(_11484_),
    .B2(_10961_),
    .Y(_11487_));
 sky130_fd_sc_hd__o21ai_4 _21524_ (.A1(_10963_),
    .A2(_10987_),
    .B1(_11481_),
    .Y(_11488_));
 sky130_fd_sc_hd__o211ai_1 _21525_ (.A1(_10963_),
    .A2(_10987_),
    .B1(_11481_),
    .C1(_11483_),
    .Y(_11489_));
 sky130_fd_sc_hd__a21oi_1 _21526_ (.A1(_11481_),
    .A2(_11483_),
    .B1(_11485_),
    .Y(_11490_));
 sky130_fd_sc_hd__a22o_1 _21527_ (.A1(_10964_),
    .A2(_10986_),
    .B1(_11481_),
    .B2(_11483_),
    .X(_11491_));
 sky130_fd_sc_hd__and3_1 _21528_ (.A(_11481_),
    .B(_11483_),
    .C(_11485_),
    .X(_11492_));
 sky130_fd_sc_hd__o211ai_4 _21529_ (.A1(_10961_),
    .A2(_11484_),
    .B1(_11483_),
    .C1(_11481_),
    .Y(_11493_));
 sky130_fd_sc_hd__nor2_1 _21530_ (.A(_03916_),
    .B(_08660_),
    .Y(_11494_));
 sky130_fd_sc_hd__o311a_2 _21531_ (.A1(net26),
    .A2(_04452_),
    .A3(_06508_),
    .B1(_08657_),
    .C1(_06486_),
    .X(_11495_));
 sky130_fd_sc_hd__a31o_2 _21532_ (.A1(_06486_),
    .A2(net262),
    .A3(_08657_),
    .B1(_11494_),
    .X(_11496_));
 sky130_fd_sc_hd__a31oi_2 _21533_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_11496_),
    .Y(_11498_));
 sky130_fd_sc_hd__and3_1 _21534_ (.A(_11496_),
    .B(net33),
    .C(net319),
    .X(_11499_));
 sky130_fd_sc_hd__o211ai_4 _21535_ (.A1(_11494_),
    .A2(_11495_),
    .B1(net33),
    .C1(net319),
    .Y(_11500_));
 sky130_fd_sc_hd__o21ai_2 _21536_ (.A1(_11498_),
    .A2(_11499_),
    .B1(net148),
    .Y(_11501_));
 sky130_fd_sc_hd__o32a_1 _21537_ (.A1(_08877_),
    .A2(_11494_),
    .A3(_11495_),
    .B1(_08881_),
    .B2(_09297_),
    .X(_11502_));
 sky130_fd_sc_hd__o21ai_1 _21538_ (.A1(_11496_),
    .A2(_08877_),
    .B1(_09300_),
    .Y(_11503_));
 sky130_fd_sc_hd__nand3b_1 _21539_ (.A_N(_11498_),
    .B(_11500_),
    .C(net148),
    .Y(_11504_));
 sky130_fd_sc_hd__o22ai_1 _21540_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_11498_),
    .B2(_11499_),
    .Y(_11505_));
 sky130_fd_sc_hd__nand2_1 _21541_ (.A(net148),
    .B(_11012_),
    .Y(_11506_));
 sky130_fd_sc_hd__o21ai_2 _21542_ (.A1(net148),
    .A2(_11010_),
    .B1(_11012_),
    .Y(_11507_));
 sky130_fd_sc_hd__o21ai_1 _21543_ (.A1(_08877_),
    .A2(_11009_),
    .B1(_11506_),
    .Y(_11509_));
 sky130_fd_sc_hd__a21oi_2 _21544_ (.A1(_11501_),
    .A2(_11503_),
    .B1(_11507_),
    .Y(_11510_));
 sky130_fd_sc_hd__nand3_2 _21545_ (.A(_11504_),
    .B(_11505_),
    .C(_11509_),
    .Y(_11511_));
 sky130_fd_sc_hd__o21ai_1 _21546_ (.A1(_11011_),
    .A2(_11013_),
    .B1(_11501_),
    .Y(_11512_));
 sky130_fd_sc_hd__nand3_2 _21547_ (.A(_11501_),
    .B(_11503_),
    .C(_11507_),
    .Y(_11513_));
 sky130_fd_sc_hd__a22o_2 _21548_ (.A1(_10541_),
    .A2(net134),
    .B1(_11511_),
    .B2(_11513_),
    .X(_11514_));
 sky130_fd_sc_hd__nand4_4 _21549_ (.A(_10541_),
    .B(net134),
    .C(_11511_),
    .D(_11513_),
    .Y(_11515_));
 sky130_fd_sc_hd__o22ai_2 _21550_ (.A1(_11013_),
    .A2(_11023_),
    .B1(_10546_),
    .B2(_11021_),
    .Y(_11516_));
 sky130_fd_sc_hd__a21oi_4 _21551_ (.A1(_11514_),
    .A2(_11515_),
    .B1(_11516_),
    .Y(_11517_));
 sky130_fd_sc_hd__a21o_2 _21552_ (.A1(_11514_),
    .A2(_11515_),
    .B1(_11516_),
    .X(_11518_));
 sky130_fd_sc_hd__o211a_2 _21553_ (.A1(_11024_),
    .A2(_11029_),
    .B1(_11514_),
    .C1(_11515_),
    .X(_11520_));
 sky130_fd_sc_hd__o211ai_4 _21554_ (.A1(_11024_),
    .A2(_11029_),
    .B1(_11514_),
    .C1(_11515_),
    .Y(_11521_));
 sky130_fd_sc_hd__and3_2 _21555_ (.A(_03927_),
    .B(net25),
    .C(net61),
    .X(_11522_));
 sky130_fd_sc_hd__a21oi_2 _21556_ (.A1(net151),
    .A2(net158),
    .B1(_06837_),
    .Y(_11523_));
 sky130_fd_sc_hd__o21ai_1 _21557_ (.A1(_08664_),
    .A2(_08666_),
    .B1(_06826_),
    .Y(_11524_));
 sky130_fd_sc_hd__a31o_1 _21558_ (.A1(net61),
    .A2(_03927_),
    .A3(net25),
    .B1(_11523_),
    .X(_11525_));
 sky130_fd_sc_hd__a31oi_4 _21559_ (.A1(_04277_),
    .A2(net162),
    .A3(_05688_),
    .B1(_11043_),
    .Y(_11526_));
 sky130_fd_sc_hd__o221ai_4 _21560_ (.A1(_04277_),
    .A2(_05720_),
    .B1(net151),
    .B2(_05699_),
    .C1(_11041_),
    .Y(_11527_));
 sky130_fd_sc_hd__nand4b_4 _21561_ (.A_N(_11522_),
    .B(_11524_),
    .C(_11526_),
    .D(net142),
    .Y(_11528_));
 sky130_fd_sc_hd__o21ai_4 _21562_ (.A1(_11522_),
    .A2(_11523_),
    .B1(_11527_),
    .Y(_11529_));
 sky130_fd_sc_hd__a2bb2oi_4 _21563_ (.A1_N(_10297_),
    .A2_N(_10538_),
    .B1(_11528_),
    .B2(_11529_),
    .Y(_11531_));
 sky130_fd_sc_hd__a2bb2o_1 _21564_ (.A1_N(_10297_),
    .A2_N(_10538_),
    .B1(_11528_),
    .B2(_11529_),
    .X(_11532_));
 sky130_fd_sc_hd__o2111a_1 _21565_ (.A1(_09755_),
    .A2(_10296_),
    .B1(_10539_),
    .C1(_11528_),
    .D1(_11529_),
    .X(_11533_));
 sky130_fd_sc_hd__o2111ai_4 _21566_ (.A1(_09755_),
    .A2(_10296_),
    .B1(_10539_),
    .C1(_11528_),
    .D1(_11529_),
    .Y(_11534_));
 sky130_fd_sc_hd__a21oi_4 _21567_ (.A1(_11038_),
    .A2(_11046_),
    .B1(_11048_),
    .Y(_11535_));
 sky130_fd_sc_hd__o22ai_4 _21568_ (.A1(_11048_),
    .A2(_11050_),
    .B1(_11531_),
    .B2(_11533_),
    .Y(_11536_));
 sky130_fd_sc_hd__nand3_4 _21569_ (.A(_11532_),
    .B(_11534_),
    .C(_11535_),
    .Y(_11537_));
 sky130_fd_sc_hd__nand2_1 _21570_ (.A(_11536_),
    .B(_11537_),
    .Y(_11538_));
 sky130_fd_sc_hd__nand4_2 _21571_ (.A(_11518_),
    .B(_11521_),
    .C(_11536_),
    .D(_11537_),
    .Y(_11539_));
 sky130_fd_sc_hd__o21ai_1 _21572_ (.A1(_11517_),
    .A2(_11520_),
    .B1(_11538_),
    .Y(_11540_));
 sky130_fd_sc_hd__o21bai_4 _21573_ (.A1(_11517_),
    .A2(_11520_),
    .B1_N(_11538_),
    .Y(_11542_));
 sky130_fd_sc_hd__nand2_1 _21574_ (.A(_11518_),
    .B(_11538_),
    .Y(_11543_));
 sky130_fd_sc_hd__nand3_2 _21575_ (.A(_11518_),
    .B(_11521_),
    .C(_11538_),
    .Y(_11544_));
 sky130_fd_sc_hd__nand3_2 _21576_ (.A(_11033_),
    .B(_11062_),
    .C(_11063_),
    .Y(_11545_));
 sky130_fd_sc_hd__a22oi_4 _21577_ (.A1(_11542_),
    .A2(_11544_),
    .B1(_11545_),
    .B2(_11035_),
    .Y(_11546_));
 sky130_fd_sc_hd__nand4_4 _21578_ (.A(_11033_),
    .B(_11067_),
    .C(_11539_),
    .D(_11540_),
    .Y(_11547_));
 sky130_fd_sc_hd__o2111a_1 _21579_ (.A1(_11520_),
    .A2(_11543_),
    .B1(_11545_),
    .C1(_11542_),
    .D1(_11035_),
    .X(_11548_));
 sky130_fd_sc_hd__nand4_4 _21580_ (.A(_11035_),
    .B(_11542_),
    .C(_11544_),
    .D(_11545_),
    .Y(_11549_));
 sky130_fd_sc_hd__nand4_2 _21581_ (.A(_11491_),
    .B(_11493_),
    .C(_11547_),
    .D(_11549_),
    .Y(_11550_));
 sky130_fd_sc_hd__o22ai_2 _21582_ (.A1(_11490_),
    .A2(_11492_),
    .B1(_11546_),
    .B2(_11548_),
    .Y(_11551_));
 sky130_fd_sc_hd__o2111ai_4 _21583_ (.A1(_11488_),
    .A2(_11482_),
    .B1(_11487_),
    .C1(_11547_),
    .D1(_11549_),
    .Y(_11553_));
 sky130_fd_sc_hd__inv_2 _21584_ (.A(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__o2bb2ai_2 _21585_ (.A1_N(_11487_),
    .A2_N(_11489_),
    .B1(_11546_),
    .B2(_11548_),
    .Y(_11555_));
 sky130_fd_sc_hd__o21ai_1 _21586_ (.A1(_11071_),
    .A2(_11425_),
    .B1(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__a2bb2oi_2 _21587_ (.A1_N(_11071_),
    .A2_N(_11425_),
    .B1(_11550_),
    .B2(_11551_),
    .Y(_11557_));
 sky130_fd_sc_hd__o211ai_2 _21588_ (.A1(_11071_),
    .A2(_11425_),
    .B1(_11553_),
    .C1(_11555_),
    .Y(_11558_));
 sky130_fd_sc_hd__a2bb2oi_2 _21589_ (.A1_N(_11068_),
    .A2_N(_11424_),
    .B1(_11553_),
    .B2(_11555_),
    .Y(_11559_));
 sky130_fd_sc_hd__o211ai_2 _21590_ (.A1(_11068_),
    .A2(_11424_),
    .B1(_11550_),
    .C1(_11551_),
    .Y(_11560_));
 sky130_fd_sc_hd__nand3_1 _21591_ (.A(_11421_),
    .B(_11422_),
    .C(_11560_),
    .Y(_11561_));
 sky130_fd_sc_hd__nand4_4 _21592_ (.A(_11421_),
    .B(_11422_),
    .C(_11558_),
    .D(_11560_),
    .Y(_11562_));
 sky130_fd_sc_hd__o2bb2ai_4 _21593_ (.A1_N(_11421_),
    .A2_N(_11422_),
    .B1(_11557_),
    .B2(_11559_),
    .Y(_11564_));
 sky130_fd_sc_hd__o21ai_2 _21594_ (.A1(_11557_),
    .A2(_11561_),
    .B1(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__o2111a_2 _21595_ (.A1(_11176_),
    .A2(_11077_),
    .B1(_11079_),
    .C1(_11562_),
    .D1(_11564_),
    .X(_11566_));
 sky130_fd_sc_hd__o2111ai_4 _21596_ (.A1(_11176_),
    .A2(_11077_),
    .B1(_11079_),
    .C1(_11562_),
    .D1(_11564_),
    .Y(_11567_));
 sky130_fd_sc_hd__a21oi_4 _21597_ (.A1(_11562_),
    .A2(_11564_),
    .B1(_11324_),
    .Y(_11568_));
 sky130_fd_sc_hd__nand2_1 _21598_ (.A(_11565_),
    .B(_11323_),
    .Y(_11569_));
 sky130_fd_sc_hd__o211ai_2 _21599_ (.A1(_11315_),
    .A2(_11316_),
    .B1(_11567_),
    .C1(_11569_),
    .Y(_11570_));
 sky130_fd_sc_hd__o22ai_2 _21600_ (.A1(_11317_),
    .A2(_11319_),
    .B1(_11566_),
    .B2(_11568_),
    .Y(_11571_));
 sky130_fd_sc_hd__a22oi_2 _21601_ (.A1(_11318_),
    .A2(_11320_),
    .B1(_11565_),
    .B2(_11323_),
    .Y(_11572_));
 sky130_fd_sc_hd__and3_1 _21602_ (.A(_11569_),
    .B(_11322_),
    .C(_11567_),
    .X(_11573_));
 sky130_fd_sc_hd__o211ai_2 _21603_ (.A1(_11317_),
    .A2(_11319_),
    .B1(_11567_),
    .C1(_11569_),
    .Y(_11575_));
 sky130_fd_sc_hd__o22ai_4 _21604_ (.A1(_11315_),
    .A2(_11316_),
    .B1(_11566_),
    .B2(_11568_),
    .Y(_11576_));
 sky130_fd_sc_hd__o21ai_1 _21605_ (.A1(_11187_),
    .A2(_11189_),
    .B1(_11576_),
    .Y(_11577_));
 sky130_fd_sc_hd__o211a_1 _21606_ (.A1(_11187_),
    .A2(_11189_),
    .B1(_11575_),
    .C1(_11576_),
    .X(_11578_));
 sky130_fd_sc_hd__o211ai_4 _21607_ (.A1(_11187_),
    .A2(_11189_),
    .B1(_11575_),
    .C1(_11576_),
    .Y(_11579_));
 sky130_fd_sc_hd__o211ai_4 _21608_ (.A1(_11185_),
    .A2(_11227_),
    .B1(_11570_),
    .C1(_11571_),
    .Y(_11580_));
 sky130_fd_sc_hd__o31a_1 _21609_ (.A1(_10824_),
    .A2(_10911_),
    .A3(_10913_),
    .B1(_10921_),
    .X(_11581_));
 sky130_fd_sc_hd__o31a_1 _21610_ (.A1(_10720_),
    .A2(_10761_),
    .A3(_10916_),
    .B1(_10918_),
    .X(_11582_));
 sky130_fd_sc_hd__a22o_1 _21611_ (.A1(_10917_),
    .A2(_10927_),
    .B1(_11579_),
    .B2(_11580_),
    .X(_11583_));
 sky130_fd_sc_hd__o2111ai_1 _21612_ (.A1(_10921_),
    .A2(_10919_),
    .B1(_10917_),
    .C1(_11580_),
    .D1(_11579_),
    .Y(_11584_));
 sky130_fd_sc_hd__o2bb2ai_2 _21613_ (.A1_N(_11579_),
    .A2_N(_11580_),
    .B1(_11581_),
    .B2(_10919_),
    .Y(_11586_));
 sky130_fd_sc_hd__o21ai_2 _21614_ (.A1(_10916_),
    .A2(_10924_),
    .B1(_11580_),
    .Y(_11587_));
 sky130_fd_sc_hd__o211ai_1 _21615_ (.A1(_10916_),
    .A2(_10924_),
    .B1(_11579_),
    .C1(_11580_),
    .Y(_11588_));
 sky130_fd_sc_hd__a22oi_1 _21616_ (.A1(_11200_),
    .A2(_11225_),
    .B1(_11586_),
    .B2(_11588_),
    .Y(_11589_));
 sky130_fd_sc_hd__a22o_1 _21617_ (.A1(_11200_),
    .A2(_11225_),
    .B1(_11586_),
    .B2(_11588_),
    .X(_11590_));
 sky130_fd_sc_hd__o221a_2 _21618_ (.A1(_11578_),
    .A2(_11587_),
    .B1(_11197_),
    .B2(_11207_),
    .C1(_11586_),
    .X(_11591_));
 sky130_fd_sc_hd__o221ai_4 _21619_ (.A1(_11578_),
    .A2(_11587_),
    .B1(_11197_),
    .B2(_11207_),
    .C1(_11586_),
    .Y(_11592_));
 sky130_fd_sc_hd__a31oi_1 _21620_ (.A1(_11226_),
    .A2(_11583_),
    .A3(_11584_),
    .B1(_11224_),
    .Y(_11593_));
 sky130_fd_sc_hd__a31o_1 _21621_ (.A1(_11226_),
    .A2(_11583_),
    .A3(_11584_),
    .B1(_11224_),
    .X(_11594_));
 sky130_fd_sc_hd__o21ai_1 _21622_ (.A1(_11589_),
    .A2(_11591_),
    .B1(_11224_),
    .Y(_11595_));
 sky130_fd_sc_hd__o2bb2ai_1 _21623_ (.A1_N(_10855_),
    .A2_N(_10861_),
    .B1(_11589_),
    .B2(_11591_),
    .Y(_11597_));
 sky130_fd_sc_hd__o2111ai_4 _21624_ (.A1(_10856_),
    .A2(_10825_),
    .B1(_10855_),
    .C1(_11590_),
    .D1(_11592_),
    .Y(_11598_));
 sky130_fd_sc_hd__o2111ai_4 _21625_ (.A1(_11211_),
    .A2(_10819_),
    .B1(_11210_),
    .C1(_11597_),
    .D1(_11598_),
    .Y(_11599_));
 sky130_fd_sc_hd__o211ai_2 _21626_ (.A1(_11591_),
    .A2(_11594_),
    .B1(_11214_),
    .C1(_11595_),
    .Y(_11600_));
 sky130_fd_sc_hd__nand2_1 _21627_ (.A(_11599_),
    .B(_11600_),
    .Y(_11601_));
 sky130_fd_sc_hd__a21boi_2 _21628_ (.A1(_10805_),
    .A2(_11220_),
    .B1_N(_11219_),
    .Y(_11602_));
 sky130_fd_sc_hd__nand4_1 _21629_ (.A(_10804_),
    .B(_10805_),
    .C(_11219_),
    .D(_11220_),
    .Y(_11603_));
 sky130_fd_sc_hd__o21ba_1 _21630_ (.A1(_11603_),
    .A2(_10812_),
    .B1_N(_11602_),
    .X(_11604_));
 sky130_fd_sc_hd__xor2_1 _21631_ (.A(_11601_),
    .B(_11604_),
    .X(net96));
 sky130_fd_sc_hd__o211a_1 _21632_ (.A1(_10862_),
    .A2(_10908_),
    .B1(_11313_),
    .C1(_10907_),
    .X(_11605_));
 sky130_fd_sc_hd__o21a_1 _21633_ (.A1(_11314_),
    .A2(_11311_),
    .B1(_11313_),
    .X(_11607_));
 sky130_fd_sc_hd__o22a_1 _21634_ (.A1(_11315_),
    .A2(_11316_),
    .B1(_11323_),
    .B2(_11565_),
    .X(_11608_));
 sky130_fd_sc_hd__o21ai_1 _21635_ (.A1(_11322_),
    .A2(_11566_),
    .B1(_11569_),
    .Y(_11609_));
 sky130_fd_sc_hd__a31oi_1 _21636_ (.A1(_11407_),
    .A2(_11411_),
    .A3(_11408_),
    .B1(_11418_),
    .Y(_11610_));
 sky130_fd_sc_hd__a41oi_4 _21637_ (.A1(_10996_),
    .A2(_11405_),
    .A3(_11406_),
    .A4(_11410_),
    .B1(_11419_),
    .Y(_11611_));
 sky130_fd_sc_hd__nand2_1 _21638_ (.A(_11248_),
    .B(_11250_),
    .Y(_11612_));
 sky130_fd_sc_hd__a22oi_4 _21639_ (.A1(_09709_),
    .A2(_07642_),
    .B1(_07643_),
    .B2(net2),
    .Y(_11613_));
 sky130_fd_sc_hd__a21o_1 _21640_ (.A1(_11235_),
    .A2(_11243_),
    .B1(_11240_),
    .X(_11614_));
 sky130_fd_sc_hd__a22oi_4 _21641_ (.A1(_11442_),
    .A2(net239),
    .B1(_07308_),
    .B2(net3),
    .Y(_11615_));
 sky130_fd_sc_hd__a32o_1 _21642_ (.A1(_11354_),
    .A2(net253),
    .A3(net239),
    .B1(_07308_),
    .B2(net3),
    .X(_11616_));
 sky130_fd_sc_hd__nor2_1 _21643_ (.A(_04004_),
    .B(_07226_),
    .Y(_11618_));
 sky130_fd_sc_hd__a31oi_2 _21644_ (.A1(net234),
    .A2(net251),
    .A3(net269),
    .B1(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__or3_1 _21645_ (.A(net51),
    .B(_04190_),
    .C(_04015_),
    .X(_11620_));
 sky130_fd_sc_hd__o211ai_4 _21646_ (.A1(net253),
    .A2(_00646_),
    .B1(net240),
    .C1(_00625_),
    .Y(_11621_));
 sky130_fd_sc_hd__o211a_4 _21647_ (.A1(_04015_),
    .A2(_06866_),
    .B1(_11621_),
    .C1(_11619_),
    .X(_11622_));
 sky130_fd_sc_hd__o211ai_1 _21648_ (.A1(_04015_),
    .A2(_06866_),
    .B1(_11621_),
    .C1(_11619_),
    .Y(_11623_));
 sky130_fd_sc_hd__a21oi_1 _21649_ (.A1(_11620_),
    .A2(_11621_),
    .B1(_11619_),
    .Y(_11624_));
 sky130_fd_sc_hd__a21o_2 _21650_ (.A1(_11620_),
    .A2(_11621_),
    .B1(_11619_),
    .X(_11625_));
 sky130_fd_sc_hd__o21ai_4 _21651_ (.A1(_11622_),
    .A2(_11624_),
    .B1(_11615_),
    .Y(_11626_));
 sky130_fd_sc_hd__nand2_1 _21652_ (.A(_11616_),
    .B(_11625_),
    .Y(_11627_));
 sky130_fd_sc_hd__nand3_1 _21653_ (.A(_11616_),
    .B(_11623_),
    .C(_11625_),
    .Y(_11629_));
 sky130_fd_sc_hd__a21oi_2 _21654_ (.A1(_11626_),
    .A2(_11629_),
    .B1(_11614_),
    .Y(_11630_));
 sky130_fd_sc_hd__a21o_1 _21655_ (.A1(_11626_),
    .A2(_11629_),
    .B1(_11614_),
    .X(_11631_));
 sky130_fd_sc_hd__o211a_1 _21656_ (.A1(_11622_),
    .A2(_11627_),
    .B1(_11626_),
    .C1(_11614_),
    .X(_11632_));
 sky130_fd_sc_hd__o211ai_4 _21657_ (.A1(_11622_),
    .A2(_11627_),
    .B1(_11626_),
    .C1(_11614_),
    .Y(_11633_));
 sky130_fd_sc_hd__o21ai_1 _21658_ (.A1(_11630_),
    .A2(_11632_),
    .B1(_11613_),
    .Y(_11634_));
 sky130_fd_sc_hd__nand3b_1 _21659_ (.A_N(_11613_),
    .B(_11631_),
    .C(_11633_),
    .Y(_11635_));
 sky130_fd_sc_hd__o21bai_1 _21660_ (.A1(_11630_),
    .A2(_11632_),
    .B1_N(_11613_),
    .Y(_11636_));
 sky130_fd_sc_hd__nand3_1 _21661_ (.A(_11631_),
    .B(_11633_),
    .C(_11613_),
    .Y(_11637_));
 sky130_fd_sc_hd__nand4_2 _21662_ (.A(_11248_),
    .B(_11250_),
    .C(_11636_),
    .D(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__and3_1 _21663_ (.A(_11612_),
    .B(_11634_),
    .C(_11635_),
    .X(_11640_));
 sky130_fd_sc_hd__nand3_1 _21664_ (.A(_11612_),
    .B(_11634_),
    .C(_11635_),
    .Y(_11641_));
 sky130_fd_sc_hd__o311a_1 _21665_ (.A1(_04747_),
    .A2(net264),
    .A3(_08656_),
    .B1(_08005_),
    .C1(_08700_),
    .X(_11642_));
 sky130_fd_sc_hd__and3_1 _21666_ (.A(_04266_),
    .B(net54),
    .C(net32),
    .X(_11643_));
 sky130_fd_sc_hd__a31o_1 _21667_ (.A1(net256),
    .A2(_08700_),
    .A3(_08005_),
    .B1(_11643_),
    .X(_11644_));
 sky130_fd_sc_hd__a21oi_2 _21668_ (.A1(_11638_),
    .A2(_11641_),
    .B1(_11644_),
    .Y(_11645_));
 sky130_fd_sc_hd__a221o_1 _21669_ (.A1(net32),
    .A2(_08006_),
    .B1(_11638_),
    .B2(_11641_),
    .C1(_11642_),
    .X(_11646_));
 sky130_fd_sc_hd__o21ai_1 _21670_ (.A1(_11642_),
    .A2(_11643_),
    .B1(_11638_),
    .Y(_11647_));
 sky130_fd_sc_hd__and3_2 _21671_ (.A(_11638_),
    .B(_11641_),
    .C(_11644_),
    .X(_11648_));
 sky130_fd_sc_hd__nor2_1 _21672_ (.A(_11645_),
    .B(_11648_),
    .Y(_11649_));
 sky130_fd_sc_hd__o21ai_1 _21673_ (.A1(_11640_),
    .A2(_11647_),
    .B1(_11646_),
    .Y(_11651_));
 sky130_fd_sc_hd__a22oi_4 _21674_ (.A1(_11293_),
    .A2(_11296_),
    .B1(_11298_),
    .B2(_11263_),
    .Y(_11652_));
 sky130_fd_sc_hd__a22o_1 _21675_ (.A1(_11293_),
    .A2(_11296_),
    .B1(_11298_),
    .B2(_11263_),
    .X(_11653_));
 sky130_fd_sc_hd__o21a_2 _21676_ (.A1(_11265_),
    .A2(_11291_),
    .B1(_11289_),
    .X(_11654_));
 sky130_fd_sc_hd__o21ai_2 _21677_ (.A1(_11265_),
    .A2(_11291_),
    .B1(_11289_),
    .Y(_11655_));
 sky130_fd_sc_hd__o22a_1 _21678_ (.A1(_11339_),
    .A2(_11344_),
    .B1(_11367_),
    .B2(_11346_),
    .X(_11656_));
 sky130_fd_sc_hd__o22ai_4 _21679_ (.A1(_11339_),
    .A2(_11344_),
    .B1(_11367_),
    .B2(_11346_),
    .Y(_11657_));
 sky130_fd_sc_hd__o21a_1 _21680_ (.A1(_11352_),
    .A2(_11357_),
    .B1(_11350_),
    .X(_11658_));
 sky130_fd_sc_hd__a21oi_2 _21681_ (.A1(_11352_),
    .A2(_11357_),
    .B1(_11350_),
    .Y(_11659_));
 sky130_fd_sc_hd__a22oi_2 _21682_ (.A1(_02464_),
    .A2(net273),
    .B1(_06326_),
    .B2(net6),
    .Y(_11660_));
 sky130_fd_sc_hd__a32o_1 _21683_ (.A1(_02421_),
    .A2(net248),
    .A3(net273),
    .B1(_06326_),
    .B2(net6),
    .X(_11662_));
 sky130_fd_sc_hd__nor2_1 _21684_ (.A(_04059_),
    .B(_05766_),
    .Y(_11663_));
 sky130_fd_sc_hd__or3b_1 _21685_ (.A(_04059_),
    .B(net48),
    .C_N(net47),
    .X(_11664_));
 sky130_fd_sc_hd__nand3_1 _21686_ (.A(net229),
    .B(net227),
    .C(net275),
    .Y(_11665_));
 sky130_fd_sc_hd__a31oi_2 _21687_ (.A1(net229),
    .A2(net227),
    .A3(net275),
    .B1(_11663_),
    .Y(_11666_));
 sky130_fd_sc_hd__nor2_1 _21688_ (.A(_04048_),
    .B(_06030_),
    .Y(_11667_));
 sky130_fd_sc_hd__o311a_1 _21689_ (.A1(net259),
    .A2(_11387_),
    .A3(_03954_),
    .B1(net274),
    .C1(_03952_),
    .X(_11668_));
 sky130_fd_sc_hd__a31oi_2 _21690_ (.A1(_03952_),
    .A2(net231),
    .A3(net274),
    .B1(_11667_),
    .Y(_11669_));
 sky130_fd_sc_hd__nand2_2 _21691_ (.A(_11666_),
    .B(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__inv_2 _21692_ (.A(_11670_),
    .Y(_11671_));
 sky130_fd_sc_hd__o2bb2ai_2 _21693_ (.A1_N(_11664_),
    .A2_N(_11665_),
    .B1(_11667_),
    .B2(_11668_),
    .Y(_11673_));
 sky130_fd_sc_hd__nand3_2 _21694_ (.A(_11670_),
    .B(_11673_),
    .C(_11660_),
    .Y(_11674_));
 sky130_fd_sc_hd__a21o_1 _21695_ (.A1(_11670_),
    .A2(_11673_),
    .B1(_11660_),
    .X(_11675_));
 sky130_fd_sc_hd__o21a_1 _21696_ (.A1(_11666_),
    .A2(_11669_),
    .B1(_11660_),
    .X(_11676_));
 sky130_fd_sc_hd__a21oi_2 _21697_ (.A1(_11666_),
    .A2(_11669_),
    .B1(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__nand3_2 _21698_ (.A(_11662_),
    .B(_11670_),
    .C(_11673_),
    .Y(_11678_));
 sky130_fd_sc_hd__a21o_1 _21699_ (.A1(_11670_),
    .A2(_11673_),
    .B1(_11662_),
    .X(_11679_));
 sky130_fd_sc_hd__a2bb2oi_2 _21700_ (.A1_N(_11358_),
    .A2_N(_11659_),
    .B1(_11674_),
    .B2(_11675_),
    .Y(_11680_));
 sky130_fd_sc_hd__o211ai_4 _21701_ (.A1(_11358_),
    .A2(_11659_),
    .B1(_11678_),
    .C1(_11679_),
    .Y(_11681_));
 sky130_fd_sc_hd__a2bb2oi_2 _21702_ (.A1_N(_11361_),
    .A2_N(_11658_),
    .B1(_11678_),
    .B2(_11679_),
    .Y(_11682_));
 sky130_fd_sc_hd__o211ai_4 _21703_ (.A1(_11361_),
    .A2(_11658_),
    .B1(_11674_),
    .C1(_11675_),
    .Y(_11684_));
 sky130_fd_sc_hd__o21a_1 _21704_ (.A1(_11279_),
    .A2(_11283_),
    .B1(_11684_),
    .X(_11685_));
 sky130_fd_sc_hd__o211ai_1 _21705_ (.A1(_11279_),
    .A2(_11283_),
    .B1(_11681_),
    .C1(_11684_),
    .Y(_11686_));
 sky130_fd_sc_hd__o22ai_1 _21706_ (.A1(_11276_),
    .A2(_11282_),
    .B1(_11680_),
    .B2(_11682_),
    .Y(_11687_));
 sky130_fd_sc_hd__a2bb2oi_2 _21707_ (.A1_N(_11279_),
    .A2_N(_11283_),
    .B1(_11681_),
    .B2(_11684_),
    .Y(_11688_));
 sky130_fd_sc_hd__a22o_1 _21708_ (.A1(_11280_),
    .A2(_11284_),
    .B1(_11681_),
    .B2(_11684_),
    .X(_11689_));
 sky130_fd_sc_hd__o211a_1 _21709_ (.A1(_11276_),
    .A2(_11282_),
    .B1(_11681_),
    .C1(_11684_),
    .X(_11690_));
 sky130_fd_sc_hd__o2111ai_4 _21710_ (.A1(_11269_),
    .A2(_11276_),
    .B1(_11280_),
    .C1(_11681_),
    .D1(_11684_),
    .Y(_11691_));
 sky130_fd_sc_hd__a21oi_1 _21711_ (.A1(_11686_),
    .A2(_11687_),
    .B1(_11657_),
    .Y(_11692_));
 sky130_fd_sc_hd__nand4_1 _21712_ (.A(_11345_),
    .B(_11371_),
    .C(_11689_),
    .D(_11691_),
    .Y(_11693_));
 sky130_fd_sc_hd__o21a_2 _21713_ (.A1(_11688_),
    .A2(_11690_),
    .B1(_11657_),
    .X(_11695_));
 sky130_fd_sc_hd__o21ai_2 _21714_ (.A1(_11688_),
    .A2(_11690_),
    .B1(_11657_),
    .Y(_11696_));
 sky130_fd_sc_hd__a21oi_1 _21715_ (.A1(_11693_),
    .A2(_11696_),
    .B1(_11655_),
    .Y(_11697_));
 sky130_fd_sc_hd__o21ai_2 _21716_ (.A1(_11692_),
    .A2(_11695_),
    .B1(_11654_),
    .Y(_11698_));
 sky130_fd_sc_hd__o31ai_4 _21717_ (.A1(_11688_),
    .A2(_11690_),
    .A3(_11657_),
    .B1(_11655_),
    .Y(_11699_));
 sky130_fd_sc_hd__nor3_1 _21718_ (.A(_11654_),
    .B(_11692_),
    .C(_11695_),
    .Y(_11700_));
 sky130_fd_sc_hd__a31o_1 _21719_ (.A1(_11657_),
    .A2(_11686_),
    .A3(_11687_),
    .B1(_11699_),
    .X(_11701_));
 sky130_fd_sc_hd__o2bb2ai_1 _21720_ (.A1_N(_11289_),
    .A2_N(_11293_),
    .B1(_11692_),
    .B2(_11695_),
    .Y(_11702_));
 sky130_fd_sc_hd__nand4_1 _21721_ (.A(_11289_),
    .B(_11293_),
    .C(_11693_),
    .D(_11696_),
    .Y(_11703_));
 sky130_fd_sc_hd__o21ai_2 _21722_ (.A1(_11695_),
    .A2(_11699_),
    .B1(_11698_),
    .Y(_11704_));
 sky130_fd_sc_hd__nand3_2 _21723_ (.A(_11702_),
    .B(_11703_),
    .C(_11652_),
    .Y(_11706_));
 sky130_fd_sc_hd__and3_1 _21724_ (.A(_11653_),
    .B(_11698_),
    .C(_11701_),
    .X(_11707_));
 sky130_fd_sc_hd__o211ai_4 _21725_ (.A1(_11699_),
    .A2(_11695_),
    .B1(_11653_),
    .C1(_11698_),
    .Y(_11708_));
 sky130_fd_sc_hd__o211a_1 _21726_ (.A1(_11645_),
    .A2(_11648_),
    .B1(_11706_),
    .C1(_11708_),
    .X(_11709_));
 sky130_fd_sc_hd__a21oi_1 _21727_ (.A1(_11706_),
    .A2(_11708_),
    .B1(_11651_),
    .Y(_11710_));
 sky130_fd_sc_hd__a2bb2oi_2 _21728_ (.A1_N(_11645_),
    .A2_N(_11648_),
    .B1(_11706_),
    .B2(_11708_),
    .Y(_11711_));
 sky130_fd_sc_hd__o211a_1 _21729_ (.A1(_11647_),
    .A2(_11640_),
    .B1(_11646_),
    .C1(_11706_),
    .X(_11712_));
 sky130_fd_sc_hd__a31o_1 _21730_ (.A1(_11652_),
    .A2(_11702_),
    .A3(_11703_),
    .B1(_11651_),
    .X(_11713_));
 sky130_fd_sc_hd__o311a_1 _21731_ (.A1(_11652_),
    .A2(_11697_),
    .A3(_11700_),
    .B1(_11706_),
    .C1(_11649_),
    .X(_11714_));
 sky130_fd_sc_hd__o22a_1 _21732_ (.A1(_11413_),
    .A2(_11610_),
    .B1(_11711_),
    .B2(_11714_),
    .X(_11715_));
 sky130_fd_sc_hd__o221ai_4 _21733_ (.A1(_11413_),
    .A2(_11419_),
    .B1(_11711_),
    .B2(_11714_),
    .C1(_11416_),
    .Y(_11717_));
 sky130_fd_sc_hd__o22a_2 _21734_ (.A1(_11415_),
    .A2(_11611_),
    .B1(_11709_),
    .B2(_11710_),
    .X(_11718_));
 sky130_fd_sc_hd__o22ai_2 _21735_ (.A1(_11415_),
    .A2(_11611_),
    .B1(_11709_),
    .B2(_11710_),
    .Y(_11719_));
 sky130_fd_sc_hd__a31o_1 _21736_ (.A1(_11257_),
    .A2(_11258_),
    .A3(_11305_),
    .B1(_11304_),
    .X(_11720_));
 sky130_fd_sc_hd__o211a_2 _21737_ (.A1(_11715_),
    .A2(_11718_),
    .B1(_11303_),
    .C1(_11306_),
    .X(_11721_));
 sky130_fd_sc_hd__o21bai_1 _21738_ (.A1(_11715_),
    .A2(_11718_),
    .B1_N(_11720_),
    .Y(_11722_));
 sky130_fd_sc_hd__nand2_1 _21739_ (.A(_11717_),
    .B(_11720_),
    .Y(_11723_));
 sky130_fd_sc_hd__and3_2 _21740_ (.A(_11717_),
    .B(_11719_),
    .C(_11720_),
    .X(_11724_));
 sky130_fd_sc_hd__a211o_1 _21741_ (.A1(_11303_),
    .A2(_11306_),
    .B1(_11715_),
    .C1(_11718_),
    .X(_11725_));
 sky130_fd_sc_hd__o21ai_2 _21742_ (.A1(_11718_),
    .A2(_11723_),
    .B1(_11722_),
    .Y(_11726_));
 sky130_fd_sc_hd__o22ai_4 _21743_ (.A1(_11554_),
    .A2(_11556_),
    .B1(_11559_),
    .B2(_11423_),
    .Y(_11728_));
 sky130_fd_sc_hd__nand3_1 _21744_ (.A(_11521_),
    .B(_11536_),
    .C(_11537_),
    .Y(_11729_));
 sky130_fd_sc_hd__a31oi_4 _21745_ (.A1(_11521_),
    .A2(_11536_),
    .A3(_11537_),
    .B1(_11517_),
    .Y(_11730_));
 sky130_fd_sc_hd__a21oi_4 _21746_ (.A1(_06826_),
    .A2(_08664_),
    .B1(_11522_),
    .Y(_11731_));
 sky130_fd_sc_hd__a31o_4 _21747_ (.A1(_04277_),
    .A2(net162),
    .A3(_06826_),
    .B1(_11522_),
    .X(_11732_));
 sky130_fd_sc_hd__a21o_1 _21748_ (.A1(net142),
    .A2(_11526_),
    .B1(_11732_),
    .X(_11733_));
 sky130_fd_sc_hd__o2111ai_4 _21749_ (.A1(_05699_),
    .A2(net151),
    .B1(_11041_),
    .C1(_11044_),
    .D1(_11732_),
    .Y(_11734_));
 sky130_fd_sc_hd__o2111a_4 _21750_ (.A1(_05699_),
    .A2(net151),
    .B1(net142),
    .C1(_11044_),
    .D1(_11731_),
    .X(_11735_));
 sky130_fd_sc_hd__o2111ai_4 _21751_ (.A1(_05699_),
    .A2(net151),
    .B1(_11041_),
    .C1(_11044_),
    .D1(_11731_),
    .Y(_11736_));
 sky130_fd_sc_hd__and3_4 _21752_ (.A(net134),
    .B(_11733_),
    .C(_11734_),
    .X(_11737_));
 sky130_fd_sc_hd__o211ai_4 _21753_ (.A1(_10297_),
    .A2(_10538_),
    .B1(_11733_),
    .C1(_11734_),
    .Y(_11739_));
 sky130_fd_sc_hd__o211a_4 _21754_ (.A1(_09755_),
    .A2(_10296_),
    .B1(_10539_),
    .C1(_11736_),
    .X(_11740_));
 sky130_fd_sc_hd__a31o_4 _21755_ (.A1(net142),
    .A2(_11526_),
    .A3(_11731_),
    .B1(net134),
    .X(_11741_));
 sky130_fd_sc_hd__o31a_4 _21756_ (.A1(_10297_),
    .A2(_10538_),
    .A3(_11735_),
    .B1(_11739_),
    .X(_11742_));
 sky130_fd_sc_hd__o21ai_4 _21757_ (.A1(net134),
    .A2(_11735_),
    .B1(_11739_),
    .Y(_11743_));
 sky130_fd_sc_hd__a22oi_2 _21758_ (.A1(_11525_),
    .A2(_11527_),
    .B1(_11739_),
    .B2(_11741_),
    .Y(_11744_));
 sky130_fd_sc_hd__o221a_1 _21759_ (.A1(_11522_),
    .A2(_11523_),
    .B1(_11732_),
    .B2(net137),
    .C1(_11527_),
    .X(_11745_));
 sky130_fd_sc_hd__o311a_1 _21760_ (.A1(_10297_),
    .A2(_10538_),
    .A3(_11735_),
    .B1(_11739_),
    .C1(_11529_),
    .X(_11746_));
 sky130_fd_sc_hd__and4_2 _21761_ (.A(_11525_),
    .B(_11731_),
    .C(_11527_),
    .D(net134),
    .X(_11747_));
 sky130_fd_sc_hd__o21a_1 _21762_ (.A1(_10540_),
    .A2(net137),
    .B1(_11513_),
    .X(_11748_));
 sky130_fd_sc_hd__o22ai_1 _21763_ (.A1(_11502_),
    .A2(_11512_),
    .B1(_10546_),
    .B2(_11510_),
    .Y(_11750_));
 sky130_fd_sc_hd__o22a_2 _21764_ (.A1(_11502_),
    .A2(_11512_),
    .B1(_10546_),
    .B2(_11510_),
    .X(_11751_));
 sky130_fd_sc_hd__nor2_1 _21765_ (.A(_03938_),
    .B(_08660_),
    .Y(_11752_));
 sky130_fd_sc_hd__a31o_2 _21766_ (.A1(_07242_),
    .A2(_07253_),
    .A3(_08657_),
    .B1(_11752_),
    .X(_11753_));
 sky130_fd_sc_hd__a31oi_4 _21767_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_11753_),
    .Y(_11754_));
 sky130_fd_sc_hd__a31o_1 _21768_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_11753_),
    .X(_11755_));
 sky130_fd_sc_hd__o2111a_1 _21769_ (.A1(net169),
    .A2(net268),
    .B1(net33),
    .C1(_11753_),
    .D1(net319),
    .X(_11756_));
 sky130_fd_sc_hd__o2111ai_4 _21770_ (.A1(net169),
    .A2(net268),
    .B1(net33),
    .C1(_11753_),
    .D1(net319),
    .Y(_11757_));
 sky130_fd_sc_hd__a21oi_2 _21771_ (.A1(_11755_),
    .A2(_11757_),
    .B1(_09300_),
    .Y(_11758_));
 sky130_fd_sc_hd__o21ai_1 _21772_ (.A1(_11754_),
    .A2(_11756_),
    .B1(net148),
    .Y(_11759_));
 sky130_fd_sc_hd__o22ai_2 _21773_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_11754_),
    .B2(_11756_),
    .Y(_11761_));
 sky130_fd_sc_hd__nand3_1 _21774_ (.A(_11755_),
    .B(_11757_),
    .C(net148),
    .Y(_11762_));
 sky130_fd_sc_hd__o211ai_4 _21775_ (.A1(net319),
    .A2(_04331_),
    .B1(_09298_),
    .C1(_11500_),
    .Y(_11763_));
 sky130_fd_sc_hd__o21ai_1 _21776_ (.A1(net148),
    .A2(_11498_),
    .B1(_11500_),
    .Y(_11764_));
 sky130_fd_sc_hd__o21ai_1 _21777_ (.A1(_11496_),
    .A2(net157),
    .B1(_11763_),
    .Y(_11765_));
 sky130_fd_sc_hd__nand3_2 _21778_ (.A(_11761_),
    .B(_11762_),
    .C(_11765_),
    .Y(_11766_));
 sky130_fd_sc_hd__o221ai_4 _21779_ (.A1(_11496_),
    .A2(_08877_),
    .B1(net148),
    .B2(_11754_),
    .C1(_11763_),
    .Y(_11767_));
 sky130_fd_sc_hd__o211ai_2 _21780_ (.A1(net148),
    .A2(_11754_),
    .B1(_11764_),
    .C1(_11759_),
    .Y(_11768_));
 sky130_fd_sc_hd__o21ai_1 _21781_ (.A1(_11767_),
    .A2(_11758_),
    .B1(_11766_),
    .Y(_11769_));
 sky130_fd_sc_hd__a2bb2oi_1 _21782_ (.A1_N(_10540_),
    .A2_N(net137),
    .B1(_11766_),
    .B2(_11768_),
    .Y(_11770_));
 sky130_fd_sc_hd__o21ai_1 _21783_ (.A1(_10540_),
    .A2(net137),
    .B1(_11769_),
    .Y(_11772_));
 sky130_fd_sc_hd__nand3_1 _21784_ (.A(net138),
    .B(net134),
    .C(_11766_),
    .Y(_11773_));
 sky130_fd_sc_hd__o2111a_1 _21785_ (.A1(_11767_),
    .A2(_11758_),
    .B1(net134),
    .C1(net138),
    .D1(_11766_),
    .X(_11774_));
 sky130_fd_sc_hd__o2111ai_4 _21786_ (.A1(_11767_),
    .A2(_11758_),
    .B1(net134),
    .C1(net138),
    .D1(_11766_),
    .Y(_11775_));
 sky130_fd_sc_hd__nand2_2 _21787_ (.A(_11772_),
    .B(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__nand3_2 _21788_ (.A(_11750_),
    .B(_11772_),
    .C(_11775_),
    .Y(_11777_));
 sky130_fd_sc_hd__o221a_1 _21789_ (.A1(_10546_),
    .A2(_11510_),
    .B1(_11770_),
    .B2(_11774_),
    .C1(_11513_),
    .X(_11778_));
 sky130_fd_sc_hd__o22ai_2 _21790_ (.A1(_11510_),
    .A2(_11748_),
    .B1(_11770_),
    .B2(_11774_),
    .Y(_11779_));
 sky130_fd_sc_hd__a2bb2oi_1 _21791_ (.A1_N(_11745_),
    .A2_N(_11746_),
    .B1(_11751_),
    .B2(_11776_),
    .Y(_11780_));
 sky130_fd_sc_hd__o21ai_1 _21792_ (.A1(_11745_),
    .A2(_11746_),
    .B1(_11779_),
    .Y(_11781_));
 sky130_fd_sc_hd__o211a_1 _21793_ (.A1(_11745_),
    .A2(_11746_),
    .B1(_11777_),
    .C1(_11779_),
    .X(_11783_));
 sky130_fd_sc_hd__o21ai_2 _21794_ (.A1(_11751_),
    .A2(_11776_),
    .B1(_11780_),
    .Y(_11784_));
 sky130_fd_sc_hd__a2bb2oi_2 _21795_ (.A1_N(_11744_),
    .A2_N(_11747_),
    .B1(_11777_),
    .B2(_11779_),
    .Y(_11785_));
 sky130_fd_sc_hd__a2bb2o_1 _21796_ (.A1_N(_11744_),
    .A2_N(_11747_),
    .B1(_11777_),
    .B2(_11779_),
    .X(_11786_));
 sky130_fd_sc_hd__a21oi_1 _21797_ (.A1(_11780_),
    .A2(_11777_),
    .B1(_11785_),
    .Y(_11787_));
 sky130_fd_sc_hd__a311o_1 _21798_ (.A1(_11521_),
    .A2(_11536_),
    .A3(_11537_),
    .B1(_11785_),
    .C1(_11517_),
    .X(_11788_));
 sky130_fd_sc_hd__and3_1 _21799_ (.A(_11784_),
    .B(_11786_),
    .C(_11730_),
    .X(_11789_));
 sky130_fd_sc_hd__nand3_4 _21800_ (.A(_11784_),
    .B(_11786_),
    .C(_11730_),
    .Y(_11790_));
 sky130_fd_sc_hd__o2bb2ai_4 _21801_ (.A1_N(_11518_),
    .A2_N(_11729_),
    .B1(_11783_),
    .B2(_11785_),
    .Y(_11791_));
 sky130_fd_sc_hd__a21oi_1 _21802_ (.A1(_11428_),
    .A2(_11439_),
    .B1(_11440_),
    .Y(_11792_));
 sky130_fd_sc_hd__a32oi_4 _21803_ (.A1(_07771_),
    .A2(net289),
    .A3(net165),
    .B1(_10335_),
    .B2(net22),
    .Y(_11794_));
 sky130_fd_sc_hd__a32o_1 _21804_ (.A1(_07771_),
    .A2(net289),
    .A3(net165),
    .B1(_10335_),
    .B2(net22),
    .X(_11795_));
 sky130_fd_sc_hd__nor2_1 _21805_ (.A(_04256_),
    .B(_08283_),
    .Y(_11796_));
 sky130_fd_sc_hd__o311a_1 _21806_ (.A1(net174),
    .A2(_07074_),
    .A3(net268),
    .B1(net291),
    .C1(net164),
    .X(_11797_));
 sky130_fd_sc_hd__a31oi_4 _21807_ (.A1(net164),
    .A2(net162),
    .A3(net291),
    .B1(_11796_),
    .Y(_11798_));
 sky130_fd_sc_hd__nor2_1 _21808_ (.A(_04277_),
    .B(_07691_),
    .Y(_11799_));
 sky130_fd_sc_hd__or3_2 _21809_ (.A(net63),
    .B(_04277_),
    .C(_03927_),
    .X(_11800_));
 sky130_fd_sc_hd__a21oi_1 _21810_ (.A1(net150),
    .A2(_08668_),
    .B1(_07669_),
    .Y(_11801_));
 sky130_fd_sc_hd__o21ai_2 _21811_ (.A1(net159),
    .A2(_08666_),
    .B1(_07658_),
    .Y(_11802_));
 sky130_fd_sc_hd__a22oi_2 _21812_ (.A1(net25),
    .A2(_07680_),
    .B1(_08670_),
    .B2(_07658_),
    .Y(_11803_));
 sky130_fd_sc_hd__o22a_2 _21813_ (.A1(_11796_),
    .A2(_11797_),
    .B1(_11799_),
    .B2(_11801_),
    .X(_11805_));
 sky130_fd_sc_hd__o22ai_1 _21814_ (.A1(_11796_),
    .A2(_11797_),
    .B1(_11799_),
    .B2(_11801_),
    .Y(_11806_));
 sky130_fd_sc_hd__a211o_1 _21815_ (.A1(_11800_),
    .A2(_11802_),
    .B1(_11794_),
    .C1(_11798_),
    .X(_11807_));
 sky130_fd_sc_hd__o311a_1 _21816_ (.A1(_03927_),
    .A2(net63),
    .A3(_04277_),
    .B1(_11798_),
    .C1(_11802_),
    .X(_11808_));
 sky130_fd_sc_hd__o211ai_2 _21817_ (.A1(_04277_),
    .A2(_07691_),
    .B1(_11798_),
    .C1(_11802_),
    .Y(_11809_));
 sky130_fd_sc_hd__o2111ai_1 _21818_ (.A1(_07669_),
    .A2(_08669_),
    .B1(_11794_),
    .C1(_11798_),
    .D1(_11800_),
    .Y(_11810_));
 sky130_fd_sc_hd__a31oi_2 _21819_ (.A1(_11802_),
    .A2(_11798_),
    .A3(_11800_),
    .B1(_11794_),
    .Y(_11811_));
 sky130_fd_sc_hd__a31o_1 _21820_ (.A1(_11802_),
    .A2(_11798_),
    .A3(_11800_),
    .B1(_11794_),
    .X(_11812_));
 sky130_fd_sc_hd__a21oi_2 _21821_ (.A1(_11795_),
    .A2(_11809_),
    .B1(_11805_),
    .Y(_11813_));
 sky130_fd_sc_hd__o211ai_2 _21822_ (.A1(_11798_),
    .A2(_11803_),
    .B1(_11810_),
    .C1(_11812_),
    .Y(_11814_));
 sky130_fd_sc_hd__a21o_1 _21823_ (.A1(_11806_),
    .A2(_11809_),
    .B1(_11795_),
    .X(_11816_));
 sky130_fd_sc_hd__o21ai_2 _21824_ (.A1(_11798_),
    .A2(_11803_),
    .B1(_11795_),
    .Y(_11817_));
 sky130_fd_sc_hd__nand3_4 _21825_ (.A(_11814_),
    .B(_11792_),
    .C(_11807_),
    .Y(_11818_));
 sky130_fd_sc_hd__o221a_2 _21826_ (.A1(_11808_),
    .A2(_11817_),
    .B1(_11440_),
    .B2(_11444_),
    .C1(_11816_),
    .X(_11819_));
 sky130_fd_sc_hd__o221ai_4 _21827_ (.A1(_11808_),
    .A2(_11817_),
    .B1(_11440_),
    .B2(_11444_),
    .C1(_11816_),
    .Y(_11820_));
 sky130_fd_sc_hd__o32a_2 _21828_ (.A1(_01304_),
    .A2(_06756_),
    .A3(net189),
    .B1(_01326_),
    .B2(_04201_),
    .X(_11821_));
 sky130_fd_sc_hd__a32o_1 _21829_ (.A1(net194),
    .A2(net171),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net19),
    .X(_11822_));
 sky130_fd_sc_hd__o211ai_4 _21830_ (.A1(net174),
    .A2(_07074_),
    .B1(_12330_),
    .C1(_07072_),
    .Y(_11823_));
 sky130_fd_sc_hd__or3_4 _21831_ (.A(net36),
    .B(_04212_),
    .C(_03993_),
    .X(_11824_));
 sky130_fd_sc_hd__nand2_1 _21832_ (.A(net167),
    .B(net252),
    .Y(_11825_));
 sky130_fd_sc_hd__a21oi_1 _21833_ (.A1(net21),
    .A2(net168),
    .B1(_11825_),
    .Y(_11827_));
 sky130_fd_sc_hd__nand3_4 _21834_ (.A(_07499_),
    .B(net167),
    .C(net252),
    .Y(_11828_));
 sky130_fd_sc_hd__and3_1 _21835_ (.A(_03993_),
    .B(net21),
    .C(net34),
    .X(_11829_));
 sky130_fd_sc_hd__or3_4 _21836_ (.A(net35),
    .B(_04223_),
    .C(_03971_),
    .X(_11830_));
 sky130_fd_sc_hd__a22oi_4 _21837_ (.A1(_11823_),
    .A2(_11824_),
    .B1(_11828_),
    .B2(_11830_),
    .Y(_11831_));
 sky130_fd_sc_hd__o2bb2ai_2 _21838_ (.A1_N(_11823_),
    .A2_N(_11824_),
    .B1(_11827_),
    .B2(_11829_),
    .Y(_11832_));
 sky130_fd_sc_hd__and4_1 _21839_ (.A(_11823_),
    .B(_11824_),
    .C(_11828_),
    .D(_11830_),
    .X(_11833_));
 sky130_fd_sc_hd__nand4_4 _21840_ (.A(_11823_),
    .B(_11824_),
    .C(_11828_),
    .D(_11830_),
    .Y(_11834_));
 sky130_fd_sc_hd__a21oi_2 _21841_ (.A1(_11832_),
    .A2(_11834_),
    .B1(_11822_),
    .Y(_11835_));
 sky130_fd_sc_hd__and3_1 _21842_ (.A(_11822_),
    .B(_11832_),
    .C(_11834_),
    .X(_11836_));
 sky130_fd_sc_hd__and3_1 _21843_ (.A(_11832_),
    .B(_11834_),
    .C(_11821_),
    .X(_11838_));
 sky130_fd_sc_hd__a21oi_2 _21844_ (.A1(_11832_),
    .A2(_11834_),
    .B1(_11821_),
    .Y(_11839_));
 sky130_fd_sc_hd__o2bb2ai_1 _21845_ (.A1_N(_11818_),
    .A2_N(_11820_),
    .B1(_11835_),
    .B2(_11836_),
    .Y(_11840_));
 sky130_fd_sc_hd__o21a_2 _21846_ (.A1(_11838_),
    .A2(_11839_),
    .B1(_11818_),
    .X(_11841_));
 sky130_fd_sc_hd__o211ai_2 _21847_ (.A1(_11838_),
    .A2(_11839_),
    .B1(_11818_),
    .C1(_11820_),
    .Y(_11842_));
 sky130_fd_sc_hd__o211ai_4 _21848_ (.A1(_11835_),
    .A2(_11836_),
    .B1(_11818_),
    .C1(_11820_),
    .Y(_11843_));
 sky130_fd_sc_hd__o2bb2ai_2 _21849_ (.A1_N(_11818_),
    .A2_N(_11820_),
    .B1(_11838_),
    .B2(_11839_),
    .Y(_11844_));
 sky130_fd_sc_hd__nand2_2 _21850_ (.A(_11843_),
    .B(_11844_),
    .Y(_11845_));
 sky130_fd_sc_hd__o21ai_4 _21851_ (.A1(_11535_),
    .A2(_11531_),
    .B1(_11534_),
    .Y(_11846_));
 sky130_fd_sc_hd__o2111ai_4 _21852_ (.A1(_11535_),
    .A2(_11531_),
    .B1(_11534_),
    .C1(_11843_),
    .D1(_11844_),
    .Y(_11847_));
 sky130_fd_sc_hd__nand3_4 _21853_ (.A(_11840_),
    .B(_11842_),
    .C(_11846_),
    .Y(_11849_));
 sky130_fd_sc_hd__o31a_2 _21854_ (.A1(_10956_),
    .A2(_11444_),
    .A3(_11446_),
    .B1(_11472_),
    .X(_11850_));
 sky130_fd_sc_hd__o31a_1 _21855_ (.A1(_11450_),
    .A2(_11470_),
    .A3(_11471_),
    .B1(_11448_),
    .X(_11851_));
 sky130_fd_sc_hd__o211a_1 _21856_ (.A1(_11449_),
    .A2(_11474_),
    .B1(_11847_),
    .C1(_11849_),
    .X(_11852_));
 sky130_fd_sc_hd__o211ai_4 _21857_ (.A1(_11449_),
    .A2(_11474_),
    .B1(_11847_),
    .C1(_11849_),
    .Y(_11853_));
 sky130_fd_sc_hd__a21boi_1 _21858_ (.A1(_11847_),
    .A2(_11849_),
    .B1_N(_11851_),
    .Y(_11854_));
 sky130_fd_sc_hd__o2bb2ai_4 _21859_ (.A1_N(_11847_),
    .A2_N(_11849_),
    .B1(_11850_),
    .B2(_11450_),
    .Y(_11855_));
 sky130_fd_sc_hd__a21oi_1 _21860_ (.A1(_11847_),
    .A2(_11849_),
    .B1(_11851_),
    .Y(_11856_));
 sky130_fd_sc_hd__a21o_1 _21861_ (.A1(_11847_),
    .A2(_11849_),
    .B1(_11851_),
    .X(_11857_));
 sky130_fd_sc_hd__o211a_1 _21862_ (.A1(_11450_),
    .A2(_11850_),
    .B1(_11849_),
    .C1(_11847_),
    .X(_11858_));
 sky130_fd_sc_hd__o2111ai_1 _21863_ (.A1(_11450_),
    .A2(_11472_),
    .B1(_11847_),
    .C1(_11849_),
    .D1(_11448_),
    .Y(_11860_));
 sky130_fd_sc_hd__nand4_2 _21864_ (.A(_11790_),
    .B(_11791_),
    .C(_11857_),
    .D(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__o2bb2ai_1 _21865_ (.A1_N(_11790_),
    .A2_N(_11791_),
    .B1(_11856_),
    .B2(_11858_),
    .Y(_11862_));
 sky130_fd_sc_hd__o2bb2ai_4 _21866_ (.A1_N(_11790_),
    .A2_N(_11791_),
    .B1(_11852_),
    .B2(_11854_),
    .Y(_11863_));
 sky130_fd_sc_hd__nand4_4 _21867_ (.A(_11790_),
    .B(_11791_),
    .C(_11853_),
    .D(_11855_),
    .Y(_11864_));
 sky130_fd_sc_hd__inv_2 _21868_ (.A(_11864_),
    .Y(_11865_));
 sky130_fd_sc_hd__nand3_1 _21869_ (.A(_11491_),
    .B(_11493_),
    .C(_11549_),
    .Y(_11866_));
 sky130_fd_sc_hd__o211ai_2 _21870_ (.A1(_11488_),
    .A2(_11482_),
    .B1(_11487_),
    .C1(_11547_),
    .Y(_11867_));
 sky130_fd_sc_hd__a31oi_4 _21871_ (.A1(_11491_),
    .A2(_11493_),
    .A3(_11549_),
    .B1(_11546_),
    .Y(_11868_));
 sky130_fd_sc_hd__a21oi_4 _21872_ (.A1(_11863_),
    .A2(_11864_),
    .B1(_11868_),
    .Y(_11869_));
 sky130_fd_sc_hd__nand4_4 _21873_ (.A(_11549_),
    .B(_11861_),
    .C(_11862_),
    .D(_11867_),
    .Y(_11871_));
 sky130_fd_sc_hd__nand2_1 _21874_ (.A(_11868_),
    .B(_11863_),
    .Y(_11872_));
 sky130_fd_sc_hd__nand4_4 _21875_ (.A(_11547_),
    .B(_11863_),
    .C(_11864_),
    .D(_11866_),
    .Y(_11873_));
 sky130_fd_sc_hd__o21ai_2 _21876_ (.A1(_10961_),
    .A2(_11484_),
    .B1(_11483_),
    .Y(_11874_));
 sky130_fd_sc_hd__a21oi_1 _21877_ (.A1(_11378_),
    .A2(_11384_),
    .B1(_11385_),
    .Y(_11875_));
 sky130_fd_sc_hd__nand3_2 _21878_ (.A(net198),
    .B(net172),
    .C(_02858_),
    .Y(_11876_));
 sky130_fd_sc_hd__or3b_2 _21879_ (.A(net38),
    .B(_04179_),
    .C_N(net37),
    .X(_11877_));
 sky130_fd_sc_hd__nor2_1 _21880_ (.A(_04168_),
    .B(_03737_),
    .Y(_11878_));
 sky130_fd_sc_hd__a31oi_4 _21881_ (.A1(net201),
    .A2(net173),
    .A3(net285),
    .B1(_11878_),
    .Y(_11879_));
 sky130_fd_sc_hd__a21oi_4 _21882_ (.A1(_11876_),
    .A2(_11877_),
    .B1(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__a21o_1 _21883_ (.A1(_11876_),
    .A2(_11877_),
    .B1(_11879_),
    .X(_11882_));
 sky130_fd_sc_hd__o211a_1 _21884_ (.A1(_04179_),
    .A2(_02891_),
    .B1(_11876_),
    .C1(_11879_),
    .X(_11883_));
 sky130_fd_sc_hd__o221ai_4 _21885_ (.A1(_04179_),
    .A2(_02891_),
    .B1(_06454_),
    .B2(_02869_),
    .C1(_11879_),
    .Y(_11884_));
 sky130_fd_sc_hd__a32o_1 _21886_ (.A1(_05933_),
    .A2(net281),
    .A3(net174),
    .B1(_04217_),
    .B2(net16),
    .X(_11885_));
 sky130_fd_sc_hd__o21bai_4 _21887_ (.A1(_11880_),
    .A2(_11883_),
    .B1_N(_11885_),
    .Y(_11886_));
 sky130_fd_sc_hd__nand3_4 _21888_ (.A(_11882_),
    .B(_11884_),
    .C(_11885_),
    .Y(_11887_));
 sky130_fd_sc_hd__inv_2 _21889_ (.A(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__a21oi_4 _21890_ (.A1(_11886_),
    .A2(_11887_),
    .B1(_11466_),
    .Y(_11889_));
 sky130_fd_sc_hd__a21o_1 _21891_ (.A1(_11886_),
    .A2(_11887_),
    .B1(_11466_),
    .X(_11890_));
 sky130_fd_sc_hd__o211a_2 _21892_ (.A1(_11462_),
    .A2(_11465_),
    .B1(_11886_),
    .C1(_11887_),
    .X(_11891_));
 sky130_fd_sc_hd__o211ai_2 _21893_ (.A1(_11462_),
    .A2(_11465_),
    .B1(_11886_),
    .C1(_11887_),
    .Y(_11893_));
 sky130_fd_sc_hd__o21ai_1 _21894_ (.A1(_11889_),
    .A2(_11891_),
    .B1(_11875_),
    .Y(_11894_));
 sky130_fd_sc_hd__o211ai_2 _21895_ (.A1(_11385_),
    .A2(_11388_),
    .B1(_11890_),
    .C1(_11893_),
    .Y(_11895_));
 sky130_fd_sc_hd__o22ai_2 _21896_ (.A1(_11385_),
    .A2(_11388_),
    .B1(_11889_),
    .B2(_11891_),
    .Y(_11896_));
 sky130_fd_sc_hd__nand3_1 _21897_ (.A(_11890_),
    .B(_11893_),
    .C(_11875_),
    .Y(_11897_));
 sky130_fd_sc_hd__o2bb2ai_1 _21898_ (.A1_N(_11374_),
    .A2_N(_11395_),
    .B1(_11391_),
    .B2(_11388_),
    .Y(_11898_));
 sky130_fd_sc_hd__nand3_4 _21899_ (.A(_11894_),
    .B(_11898_),
    .C(_11895_),
    .Y(_11899_));
 sky130_fd_sc_hd__and4_2 _21900_ (.A(_11393_),
    .B(_11396_),
    .C(_11896_),
    .D(_11897_),
    .X(_11900_));
 sky130_fd_sc_hd__nand4_4 _21901_ (.A(_11393_),
    .B(_11396_),
    .C(_11896_),
    .D(_11897_),
    .Y(_11901_));
 sky130_fd_sc_hd__nor2_1 _21902_ (.A(_04069_),
    .B(_05465_),
    .Y(_11902_));
 sky130_fd_sc_hd__o311a_1 _21903_ (.A1(net7),
    .A2(net248),
    .A3(_04407_),
    .B1(_05462_),
    .C1(net221),
    .X(_11904_));
 sky130_fd_sc_hd__a21oi_2 _21904_ (.A1(net9),
    .A2(_05464_),
    .B1(_11904_),
    .Y(_11905_));
 sky130_fd_sc_hd__and3_1 _21905_ (.A(_04124_),
    .B(net43),
    .C(net11),
    .X(_11906_));
 sky130_fd_sc_hd__a31oi_4 _21906_ (.A1(net184),
    .A2(net214),
    .A3(net242),
    .B1(_11906_),
    .Y(_11907_));
 sky130_fd_sc_hd__a32oi_4 _21907_ (.A1(net217),
    .A2(net186),
    .A3(net276),
    .B1(_05228_),
    .B2(net10),
    .Y(_11908_));
 sky130_fd_sc_hd__nor2_2 _21908_ (.A(_11907_),
    .B(_11908_),
    .Y(_11909_));
 sky130_fd_sc_hd__o221a_1 _21909_ (.A1(_04562_),
    .A2(_05226_),
    .B1(_05229_),
    .B2(_04080_),
    .C1(_11907_),
    .X(_11910_));
 sky130_fd_sc_hd__nand2_1 _21910_ (.A(_11907_),
    .B(_11908_),
    .Y(_11911_));
 sky130_fd_sc_hd__o22ai_4 _21911_ (.A1(_11902_),
    .A2(_11904_),
    .B1(_11909_),
    .B2(_11910_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand3b_4 _21912_ (.A_N(_11909_),
    .B(_11911_),
    .C(_11905_),
    .Y(_11913_));
 sky130_fd_sc_hd__nand2_2 _21913_ (.A(_11912_),
    .B(_11913_),
    .Y(_11915_));
 sky130_fd_sc_hd__a21oi_4 _21914_ (.A1(_11327_),
    .A2(_11338_),
    .B1(_11335_),
    .Y(_11916_));
 sky130_fd_sc_hd__nor2_1 _21915_ (.A(_04146_),
    .B(_04270_),
    .Y(_11917_));
 sky130_fd_sc_hd__or3b_1 _21916_ (.A(net41),
    .B(_04146_),
    .C_N(net40),
    .X(_11918_));
 sky130_fd_sc_hd__a211oi_2 _21917_ (.A1(_04788_),
    .A2(_05550_),
    .B1(_04268_),
    .C1(_05548_),
    .Y(_11919_));
 sky130_fd_sc_hd__o211ai_2 _21918_ (.A1(net184),
    .A2(_05551_),
    .B1(_04267_),
    .C1(net178),
    .Y(_11920_));
 sky130_fd_sc_hd__nand3_2 _21919_ (.A(net182),
    .B(net179),
    .C(net279),
    .Y(_11921_));
 sky130_fd_sc_hd__or3b_1 _21920_ (.A(net42),
    .B(_04135_),
    .C_N(net41),
    .X(_11922_));
 sky130_fd_sc_hd__o21ai_1 _21921_ (.A1(_04135_),
    .A2(_04483_),
    .B1(_11921_),
    .Y(_11923_));
 sky130_fd_sc_hd__o2111ai_4 _21922_ (.A1(_04146_),
    .A2(_04270_),
    .B1(_11920_),
    .C1(_11921_),
    .D1(_11922_),
    .Y(_11924_));
 sky130_fd_sc_hd__a22oi_1 _21923_ (.A1(_11918_),
    .A2(_11920_),
    .B1(_11921_),
    .B2(_11922_),
    .Y(_11926_));
 sky130_fd_sc_hd__o21ai_4 _21924_ (.A1(_11917_),
    .A2(_11919_),
    .B1(_11923_),
    .Y(_11927_));
 sky130_fd_sc_hd__nand2_1 _21925_ (.A(_11924_),
    .B(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__and3_1 _21926_ (.A(_04102_),
    .B(net13),
    .C(net42),
    .X(_11929_));
 sky130_fd_sc_hd__o311a_1 _21927_ (.A1(net11),
    .A2(_04557_),
    .A3(net208),
    .B1(_04895_),
    .C1(net210),
    .X(_11930_));
 sky130_fd_sc_hd__o22a_1 _21928_ (.A1(_04113_),
    .A2(_04898_),
    .B1(_05077_),
    .B2(_04896_),
    .X(_11931_));
 sky130_fd_sc_hd__a31o_1 _21929_ (.A1(net210),
    .A2(net183),
    .A3(_04895_),
    .B1(_11929_),
    .X(_11932_));
 sky130_fd_sc_hd__o211a_2 _21930_ (.A1(_11929_),
    .A2(_11930_),
    .B1(_11924_),
    .C1(_11927_),
    .X(_11933_));
 sky130_fd_sc_hd__o211ai_4 _21931_ (.A1(_11929_),
    .A2(_11930_),
    .B1(_11924_),
    .C1(_11927_),
    .Y(_11934_));
 sky130_fd_sc_hd__a21oi_4 _21932_ (.A1(_11924_),
    .A2(_11927_),
    .B1(_11932_),
    .Y(_11935_));
 sky130_fd_sc_hd__a21oi_1 _21933_ (.A1(_11928_),
    .A2(_11931_),
    .B1(_11916_),
    .Y(_11937_));
 sky130_fd_sc_hd__o2bb2ai_1 _21934_ (.A1_N(_11928_),
    .A2_N(_11931_),
    .B1(_11335_),
    .B2(_11339_),
    .Y(_11938_));
 sky130_fd_sc_hd__o21a_1 _21935_ (.A1(_11928_),
    .A2(_11931_),
    .B1(_11937_),
    .X(_11939_));
 sky130_fd_sc_hd__a211o_1 _21936_ (.A1(_11336_),
    .A2(_11340_),
    .B1(_11933_),
    .C1(_11935_),
    .X(_11940_));
 sky130_fd_sc_hd__o21ai_4 _21937_ (.A1(_11933_),
    .A2(_11935_),
    .B1(_11916_),
    .Y(_11941_));
 sky130_fd_sc_hd__o2111a_1 _21938_ (.A1(_11933_),
    .A2(_11938_),
    .B1(_11941_),
    .C1(_11913_),
    .D1(_11912_),
    .X(_11942_));
 sky130_fd_sc_hd__o2111ai_1 _21939_ (.A1(_11933_),
    .A2(_11938_),
    .B1(_11941_),
    .C1(_11913_),
    .D1(_11912_),
    .Y(_11943_));
 sky130_fd_sc_hd__a22oi_4 _21940_ (.A1(_11912_),
    .A2(_11913_),
    .B1(_11940_),
    .B2(_11941_),
    .Y(_11944_));
 sky130_fd_sc_hd__a22o_1 _21941_ (.A1(_11912_),
    .A2(_11913_),
    .B1(_11940_),
    .B2(_11941_),
    .X(_11945_));
 sky130_fd_sc_hd__o311a_1 _21942_ (.A1(_11916_),
    .A2(_11933_),
    .A3(_11935_),
    .B1(_11915_),
    .C1(_11941_),
    .X(_11946_));
 sky130_fd_sc_hd__a21oi_2 _21943_ (.A1(_11940_),
    .A2(_11941_),
    .B1(_11915_),
    .Y(_11948_));
 sky130_fd_sc_hd__o2bb2ai_4 _21944_ (.A1_N(_11899_),
    .A2_N(_11901_),
    .B1(_11942_),
    .B2(_11944_),
    .Y(_11949_));
 sky130_fd_sc_hd__o211ai_4 _21945_ (.A1(_11946_),
    .A2(_11948_),
    .B1(_11899_),
    .C1(_11901_),
    .Y(_11950_));
 sky130_fd_sc_hd__o2bb2ai_1 _21946_ (.A1_N(_11899_),
    .A2_N(_11901_),
    .B1(_11946_),
    .B2(_11948_),
    .Y(_11951_));
 sky130_fd_sc_hd__o211ai_2 _21947_ (.A1(_11942_),
    .A2(_11944_),
    .B1(_11899_),
    .C1(_11901_),
    .Y(_11952_));
 sky130_fd_sc_hd__nand4_4 _21948_ (.A(_11483_),
    .B(_11488_),
    .C(_11949_),
    .D(_11950_),
    .Y(_11953_));
 sky130_fd_sc_hd__a22oi_4 _21949_ (.A1(_11483_),
    .A2(_11488_),
    .B1(_11949_),
    .B2(_11950_),
    .Y(_11954_));
 sky130_fd_sc_hd__nand4_4 _21950_ (.A(_11481_),
    .B(_11874_),
    .C(_11951_),
    .D(_11952_),
    .Y(_11955_));
 sky130_fd_sc_hd__o21a_1 _21951_ (.A1(_11368_),
    .A2(_11370_),
    .B1(_11402_),
    .X(_11956_));
 sky130_fd_sc_hd__a31o_1 _21952_ (.A1(_11369_),
    .A2(_11371_),
    .A3(_11404_),
    .B1(_11401_),
    .X(_11957_));
 sky130_fd_sc_hd__a31oi_2 _21953_ (.A1(_11369_),
    .A2(_11371_),
    .A3(_11404_),
    .B1(_11401_),
    .Y(_11959_));
 sky130_fd_sc_hd__and3_1 _21954_ (.A(_11953_),
    .B(_11955_),
    .C(_11957_),
    .X(_11960_));
 sky130_fd_sc_hd__nand3_2 _21955_ (.A(_11953_),
    .B(_11955_),
    .C(_11957_),
    .Y(_11961_));
 sky130_fd_sc_hd__o2bb2a_1 _21956_ (.A1_N(_11953_),
    .A2_N(_11955_),
    .B1(_11956_),
    .B2(_11403_),
    .X(_11962_));
 sky130_fd_sc_hd__o2bb2ai_4 _21957_ (.A1_N(_11953_),
    .A2_N(_11955_),
    .B1(_11956_),
    .B2(_11403_),
    .Y(_11963_));
 sky130_fd_sc_hd__nand2_1 _21958_ (.A(_11961_),
    .B(_11963_),
    .Y(_11964_));
 sky130_fd_sc_hd__nand4_4 _21959_ (.A(_11871_),
    .B(_11873_),
    .C(_11961_),
    .D(_11963_),
    .Y(_11965_));
 sky130_fd_sc_hd__inv_2 _21960_ (.A(_11965_),
    .Y(_11966_));
 sky130_fd_sc_hd__o2bb2ai_4 _21961_ (.A1_N(_11871_),
    .A2_N(_11873_),
    .B1(_11960_),
    .B2(_11962_),
    .Y(_11967_));
 sky130_fd_sc_hd__a21oi_4 _21962_ (.A1(_11965_),
    .A2(_11967_),
    .B1(_11728_),
    .Y(_11968_));
 sky130_fd_sc_hd__a21o_1 _21963_ (.A1(_11965_),
    .A2(_11967_),
    .B1(_11728_),
    .X(_11970_));
 sky130_fd_sc_hd__nand2_1 _21964_ (.A(_11728_),
    .B(_11967_),
    .Y(_11971_));
 sky130_fd_sc_hd__and3_1 _21965_ (.A(_11728_),
    .B(_11965_),
    .C(_11967_),
    .X(_11972_));
 sky130_fd_sc_hd__nand3_2 _21966_ (.A(_11728_),
    .B(_11965_),
    .C(_11967_),
    .Y(_11973_));
 sky130_fd_sc_hd__nand3b_2 _21967_ (.A_N(_11726_),
    .B(_11970_),
    .C(_11973_),
    .Y(_11974_));
 sky130_fd_sc_hd__o22ai_4 _21968_ (.A1(_11721_),
    .A2(_11724_),
    .B1(_11968_),
    .B2(_11972_),
    .Y(_11975_));
 sky130_fd_sc_hd__o221ai_4 _21969_ (.A1(_11966_),
    .A2(_11971_),
    .B1(_11721_),
    .B2(_11724_),
    .C1(_11970_),
    .Y(_11976_));
 sky130_fd_sc_hd__a21o_1 _21970_ (.A1(_11970_),
    .A2(_11973_),
    .B1(_11726_),
    .X(_11977_));
 sky130_fd_sc_hd__a2bb2oi_1 _21971_ (.A1_N(_11568_),
    .A2_N(_11608_),
    .B1(_11974_),
    .B2(_11975_),
    .Y(_11978_));
 sky130_fd_sc_hd__o211ai_4 _21972_ (.A1(_11568_),
    .A2(_11608_),
    .B1(_11976_),
    .C1(_11977_),
    .Y(_11979_));
 sky130_fd_sc_hd__o211a_2 _21973_ (.A1(_11566_),
    .A2(_11572_),
    .B1(_11974_),
    .C1(_11975_),
    .X(_11981_));
 sky130_fd_sc_hd__o211ai_4 _21974_ (.A1(_11566_),
    .A2(_11572_),
    .B1(_11974_),
    .C1(_11975_),
    .Y(_11982_));
 sky130_fd_sc_hd__o21ai_1 _21975_ (.A1(_11978_),
    .A2(_11981_),
    .B1(_11607_),
    .Y(_11983_));
 sky130_fd_sc_hd__a31oi_1 _21976_ (.A1(_11977_),
    .A2(_11609_),
    .A3(_11976_),
    .B1(_11607_),
    .Y(_11984_));
 sky130_fd_sc_hd__a31o_1 _21977_ (.A1(_11977_),
    .A2(_11609_),
    .A3(_11976_),
    .B1(_11607_),
    .X(_11985_));
 sky130_fd_sc_hd__o21bai_1 _21978_ (.A1(_11978_),
    .A2(_11981_),
    .B1_N(_11607_),
    .Y(_11986_));
 sky130_fd_sc_hd__o2111ai_4 _21979_ (.A1(_11314_),
    .A2(_11311_),
    .B1(_11313_),
    .C1(_11979_),
    .D1(_11982_),
    .Y(_11987_));
 sky130_fd_sc_hd__o2bb2ai_2 _21980_ (.A1_N(_11580_),
    .A2_N(_11582_),
    .B1(_11573_),
    .B2(_11577_),
    .Y(_11988_));
 sky130_fd_sc_hd__a21oi_1 _21981_ (.A1(_11580_),
    .A2(_11582_),
    .B1(_11578_),
    .Y(_11989_));
 sky130_fd_sc_hd__nand3_4 _21982_ (.A(_11986_),
    .B(_11987_),
    .C(_11989_),
    .Y(_11990_));
 sky130_fd_sc_hd__o211ai_4 _21983_ (.A1(_11981_),
    .A2(_11985_),
    .B1(_11988_),
    .C1(_11983_),
    .Y(_11992_));
 sky130_fd_sc_hd__a311oi_2 _21984_ (.A1(net31),
    .A2(net54),
    .A3(_04266_),
    .B1(_11230_),
    .C1(_11254_),
    .Y(_11993_));
 sky130_fd_sc_hd__o21a_1 _21985_ (.A1(_11229_),
    .A2(_11230_),
    .B1(_11253_),
    .X(_11994_));
 sky130_fd_sc_hd__o21a_1 _21986_ (.A1(_11231_),
    .A2(_11252_),
    .B1(_11256_),
    .X(_11995_));
 sky130_fd_sc_hd__o211a_1 _21987_ (.A1(_11254_),
    .A2(_11994_),
    .B1(_11992_),
    .C1(_11990_),
    .X(_11996_));
 sky130_fd_sc_hd__o2bb2ai_1 _21988_ (.A1_N(_11990_),
    .A2_N(_11992_),
    .B1(_11993_),
    .B2(_11252_),
    .Y(_11997_));
 sky130_fd_sc_hd__o2bb2ai_1 _21989_ (.A1_N(_11990_),
    .A2_N(_11992_),
    .B1(_11994_),
    .B2(_11254_),
    .Y(_11998_));
 sky130_fd_sc_hd__o2111ai_2 _21990_ (.A1(_11231_),
    .A2(_11252_),
    .B1(_11256_),
    .C1(_11990_),
    .D1(_11992_),
    .Y(_11999_));
 sky130_fd_sc_hd__nand4_2 _21991_ (.A(_11592_),
    .B(_11594_),
    .C(_11998_),
    .D(_11999_),
    .Y(_12000_));
 sky130_fd_sc_hd__o21ai_2 _21992_ (.A1(_11591_),
    .A2(_11593_),
    .B1(_11997_),
    .Y(_12001_));
 sky130_fd_sc_hd__o21ai_1 _21993_ (.A1(_11996_),
    .A2(_12001_),
    .B1(_12000_),
    .Y(_12003_));
 sky130_fd_sc_hd__o21a_1 _21994_ (.A1(_11601_),
    .A2(_11604_),
    .B1(_11600_),
    .X(_12004_));
 sky130_fd_sc_hd__xor2_1 _21995_ (.A(_12003_),
    .B(_12004_),
    .X(net97));
 sky130_fd_sc_hd__o21ai_1 _21996_ (.A1(_11311_),
    .A2(_11605_),
    .B1(_11982_),
    .Y(_12005_));
 sky130_fd_sc_hd__a32oi_4 _21997_ (.A1(_11868_),
    .A2(_11864_),
    .A3(_11863_),
    .B1(_11963_),
    .B2(_11961_),
    .Y(_12006_));
 sky130_fd_sc_hd__o22ai_2 _21998_ (.A1(_11865_),
    .A2(_11872_),
    .B1(_11964_),
    .B2(_11869_),
    .Y(_12007_));
 sky130_fd_sc_hd__o22a_1 _21999_ (.A1(_11865_),
    .A2(_11872_),
    .B1(_11964_),
    .B2(_11869_),
    .X(_12008_));
 sky130_fd_sc_hd__o211ai_1 _22000_ (.A1(_11730_),
    .A2(_11787_),
    .B1(_11853_),
    .C1(_11855_),
    .Y(_12009_));
 sky130_fd_sc_hd__o21ai_2 _22001_ (.A1(_11783_),
    .A2(_11788_),
    .B1(_12009_),
    .Y(_12010_));
 sky130_fd_sc_hd__a31oi_4 _22002_ (.A1(_11791_),
    .A2(_11853_),
    .A3(_11855_),
    .B1(_11789_),
    .Y(_12011_));
 sky130_fd_sc_hd__a22o_1 _22003_ (.A1(_11736_),
    .A2(net137),
    .B1(_11525_),
    .B2(_11527_),
    .X(_12013_));
 sky130_fd_sc_hd__a31o_2 _22004_ (.A1(_11525_),
    .A2(_11527_),
    .A3(_11739_),
    .B1(_11740_),
    .X(_12014_));
 sky130_fd_sc_hd__and3_1 _22005_ (.A(_03927_),
    .B(_04277_),
    .C(net63),
    .X(_12015_));
 sky130_fd_sc_hd__or3b_4 _22006_ (.A(net62),
    .B(net25),
    .C_N(net63),
    .X(_12016_));
 sky130_fd_sc_hd__a31o_1 _22007_ (.A1(_07502_),
    .A2(_04256_),
    .A3(_04245_),
    .B1(_12016_),
    .X(_12017_));
 sky130_fd_sc_hd__a21oi_2 _22008_ (.A1(net162),
    .A2(_12015_),
    .B1(_11799_),
    .Y(_12018_));
 sky130_fd_sc_hd__a21oi_2 _22009_ (.A1(net150),
    .A2(_08668_),
    .B1(_08261_),
    .Y(_12019_));
 sky130_fd_sc_hd__o21ai_1 _22010_ (.A1(net159),
    .A2(_08666_),
    .B1(net291),
    .Y(_12020_));
 sky130_fd_sc_hd__nor2_1 _22011_ (.A(_04277_),
    .B(_08283_),
    .Y(_12021_));
 sky130_fd_sc_hd__or3b_4 _22012_ (.A(net64),
    .B(_04277_),
    .C_N(net63),
    .X(_12022_));
 sky130_fd_sc_hd__o221ai_4 _22013_ (.A1(_04277_),
    .A2(_07691_),
    .B1(_12016_),
    .B2(net154),
    .C1(_12022_),
    .Y(_12024_));
 sky130_fd_sc_hd__a21oi_4 _22014_ (.A1(_08670_),
    .A2(net291),
    .B1(_12024_),
    .Y(_12025_));
 sky130_fd_sc_hd__o32a_4 _22015_ (.A1(_10324_),
    .A2(_08203_),
    .A3(net154),
    .B1(_10346_),
    .B2(_04256_),
    .X(_12026_));
 sky130_fd_sc_hd__a32o_1 _22016_ (.A1(net164),
    .A2(net162),
    .A3(net289),
    .B1(_10335_),
    .B2(net24),
    .X(_12027_));
 sky130_fd_sc_hd__a22oi_2 _22017_ (.A1(_11800_),
    .A2(_12017_),
    .B1(_12020_),
    .B2(_12022_),
    .Y(_12028_));
 sky130_fd_sc_hd__o21bai_4 _22018_ (.A1(_12019_),
    .A2(_12021_),
    .B1_N(_12018_),
    .Y(_12029_));
 sky130_fd_sc_hd__o211ai_2 _22019_ (.A1(_12019_),
    .A2(_12024_),
    .B1(_12026_),
    .C1(_12029_),
    .Y(_12030_));
 sky130_fd_sc_hd__o21ai_1 _22020_ (.A1(_12025_),
    .A2(_12028_),
    .B1(_12027_),
    .Y(_12031_));
 sky130_fd_sc_hd__o21a_1 _22021_ (.A1(_12024_),
    .A2(_12019_),
    .B1(_12027_),
    .X(_12032_));
 sky130_fd_sc_hd__o21ai_1 _22022_ (.A1(_12024_),
    .A2(_12019_),
    .B1(_12027_),
    .Y(_12033_));
 sky130_fd_sc_hd__o21a_1 _22023_ (.A1(_12025_),
    .A2(_12028_),
    .B1(_12026_),
    .X(_12035_));
 sky130_fd_sc_hd__o21ai_2 _22024_ (.A1(_12025_),
    .A2(_12028_),
    .B1(_12026_),
    .Y(_12036_));
 sky130_fd_sc_hd__o221a_1 _22025_ (.A1(_11805_),
    .A2(_11811_),
    .B1(_12025_),
    .B2(_12026_),
    .C1(_12036_),
    .X(_12037_));
 sky130_fd_sc_hd__o221ai_4 _22026_ (.A1(_11805_),
    .A2(_11811_),
    .B1(_12025_),
    .B2(_12026_),
    .C1(_12036_),
    .Y(_12038_));
 sky130_fd_sc_hd__nand3_4 _22027_ (.A(_12031_),
    .B(_11813_),
    .C(_12030_),
    .Y(_12039_));
 sky130_fd_sc_hd__nor2_1 _22028_ (.A(_04212_),
    .B(_01326_),
    .Y(_12040_));
 sky130_fd_sc_hd__o311a_1 _22029_ (.A1(net246),
    .A2(_05928_),
    .A3(_07074_),
    .B1(_01293_),
    .C1(_07072_),
    .X(_12041_));
 sky130_fd_sc_hd__a31o_1 _22030_ (.A1(_07072_),
    .A2(net168),
    .A3(_01293_),
    .B1(_12040_),
    .X(_12042_));
 sky130_fd_sc_hd__nor2_1 _22031_ (.A(_04223_),
    .B(_12363_),
    .Y(_12043_));
 sky130_fd_sc_hd__a31oi_4 _22032_ (.A1(_07499_),
    .A2(net167),
    .A3(_12330_),
    .B1(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__and3_1 _22033_ (.A(_03993_),
    .B(net22),
    .C(net34),
    .X(_12046_));
 sky130_fd_sc_hd__and3_1 _22034_ (.A(_07771_),
    .B(net252),
    .C(net165),
    .X(_12047_));
 sky130_fd_sc_hd__a31oi_2 _22035_ (.A1(_07771_),
    .A2(net252),
    .A3(net165),
    .B1(_12046_),
    .Y(_12048_));
 sky130_fd_sc_hd__nand2_2 _22036_ (.A(_12044_),
    .B(_12048_),
    .Y(_12049_));
 sky130_fd_sc_hd__o21bai_2 _22037_ (.A1(_12046_),
    .A2(_12047_),
    .B1_N(_12044_),
    .Y(_12050_));
 sky130_fd_sc_hd__a21oi_1 _22038_ (.A1(_12049_),
    .A2(_12050_),
    .B1(_12042_),
    .Y(_12051_));
 sky130_fd_sc_hd__a221o_1 _22039_ (.A1(net20),
    .A2(_01315_),
    .B1(_12049_),
    .B2(_12050_),
    .C1(_12041_),
    .X(_12052_));
 sky130_fd_sc_hd__and3_1 _22040_ (.A(_12042_),
    .B(_12049_),
    .C(_12050_),
    .X(_12053_));
 sky130_fd_sc_hd__o211ai_4 _22041_ (.A1(_12040_),
    .A2(_12041_),
    .B1(_12049_),
    .C1(_12050_),
    .Y(_12054_));
 sky130_fd_sc_hd__o2bb2ai_4 _22042_ (.A1_N(_12038_),
    .A2_N(_12039_),
    .B1(_12051_),
    .B2(_12053_),
    .Y(_12055_));
 sky130_fd_sc_hd__nand3_4 _22043_ (.A(_12039_),
    .B(_12052_),
    .C(_12054_),
    .Y(_12057_));
 sky130_fd_sc_hd__nand4_2 _22044_ (.A(_12038_),
    .B(_12039_),
    .C(_12052_),
    .D(_12054_),
    .Y(_12058_));
 sky130_fd_sc_hd__o21a_1 _22045_ (.A1(_12037_),
    .A2(_12057_),
    .B1(_12055_),
    .X(_12059_));
 sky130_fd_sc_hd__a22oi_4 _22046_ (.A1(_11739_),
    .A2(_12013_),
    .B1(_12055_),
    .B2(_12058_),
    .Y(_12060_));
 sky130_fd_sc_hd__o221a_1 _22047_ (.A1(_11740_),
    .A2(_11747_),
    .B1(_12037_),
    .B2(_12057_),
    .C1(_12055_),
    .X(_12061_));
 sky130_fd_sc_hd__o221ai_4 _22048_ (.A1(_11740_),
    .A2(_11747_),
    .B1(_12037_),
    .B2(_12057_),
    .C1(_12055_),
    .Y(_12062_));
 sky130_fd_sc_hd__nor2_2 _22049_ (.A(_11819_),
    .B(_11841_),
    .Y(_12063_));
 sky130_fd_sc_hd__o22ai_4 _22050_ (.A1(_11819_),
    .A2(_11841_),
    .B1(_12060_),
    .B2(_12061_),
    .Y(_12064_));
 sky130_fd_sc_hd__nand2_2 _22051_ (.A(_12062_),
    .B(_12063_),
    .Y(_12065_));
 sky130_fd_sc_hd__o21ai_1 _22052_ (.A1(_12060_),
    .A2(_12061_),
    .B1(_12063_),
    .Y(_12066_));
 sky130_fd_sc_hd__o221ai_4 _22053_ (.A1(_11819_),
    .A2(_11841_),
    .B1(_12014_),
    .B2(_12059_),
    .C1(_12062_),
    .Y(_12068_));
 sky130_fd_sc_hd__o21ai_1 _22054_ (.A1(_12060_),
    .A2(_12065_),
    .B1(_12064_),
    .Y(_12069_));
 sky130_fd_sc_hd__o22a_1 _22055_ (.A1(_11744_),
    .A2(_11747_),
    .B1(_11751_),
    .B2(_11776_),
    .X(_12070_));
 sky130_fd_sc_hd__o21ai_2 _22056_ (.A1(_11751_),
    .A2(_11776_),
    .B1(_11781_),
    .Y(_12071_));
 sky130_fd_sc_hd__a31o_1 _22057_ (.A1(net309),
    .A2(net295),
    .A3(_08645_),
    .B1(_08658_),
    .X(_12072_));
 sky130_fd_sc_hd__o22ai_4 _22058_ (.A1(_03949_),
    .A2(_08660_),
    .B1(_08689_),
    .B2(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__a31oi_4 _22059_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_12073_),
    .Y(_12074_));
 sky130_fd_sc_hd__and4_1 _22060_ (.A(net161),
    .B(net33),
    .C(net319),
    .D(_12073_),
    .X(_12075_));
 sky130_fd_sc_hd__o2111ai_4 _22061_ (.A1(net169),
    .A2(net268),
    .B1(_12073_),
    .C1(net319),
    .D1(net33),
    .Y(_12076_));
 sky130_fd_sc_hd__o21ai_4 _22062_ (.A1(_12074_),
    .A2(_12075_),
    .B1(net147),
    .Y(_12077_));
 sky130_fd_sc_hd__o21ai_4 _22063_ (.A1(_12073_),
    .A2(net156),
    .B1(_09300_),
    .Y(_12079_));
 sky130_fd_sc_hd__o21ai_2 _22064_ (.A1(_12074_),
    .A2(_12075_),
    .B1(_09300_),
    .Y(_12080_));
 sky130_fd_sc_hd__nand3b_2 _22065_ (.A_N(_12074_),
    .B(_12076_),
    .C(net147),
    .Y(_12081_));
 sky130_fd_sc_hd__o21ai_4 _22066_ (.A1(net148),
    .A2(_11754_),
    .B1(_11757_),
    .Y(_12082_));
 sky130_fd_sc_hd__o21a_1 _22067_ (.A1(net148),
    .A2(_11754_),
    .B1(_11757_),
    .X(_12083_));
 sky130_fd_sc_hd__a21oi_1 _22068_ (.A1(_12077_),
    .A2(_12079_),
    .B1(_12082_),
    .Y(_12084_));
 sky130_fd_sc_hd__nand3_2 _22069_ (.A(_12080_),
    .B(_12081_),
    .C(_12083_),
    .Y(_12085_));
 sky130_fd_sc_hd__o211ai_4 _22070_ (.A1(net147),
    .A2(_12074_),
    .B1(_12082_),
    .C1(_12077_),
    .Y(_12086_));
 sky130_fd_sc_hd__a22o_1 _22071_ (.A1(net138),
    .A2(net134),
    .B1(_12085_),
    .B2(_12086_),
    .X(_12087_));
 sky130_fd_sc_hd__nand4_1 _22072_ (.A(net138),
    .B(net134),
    .C(_12085_),
    .D(_12086_),
    .Y(_12088_));
 sky130_fd_sc_hd__o211ai_2 _22073_ (.A1(_10540_),
    .A2(net137),
    .B1(_12085_),
    .C1(_12086_),
    .Y(_12090_));
 sky130_fd_sc_hd__a21o_1 _22074_ (.A1(_12085_),
    .A2(_12086_),
    .B1(_10546_),
    .X(_12091_));
 sky130_fd_sc_hd__o21ai_1 _22075_ (.A1(_11758_),
    .A2(_11767_),
    .B1(_11773_),
    .Y(_12092_));
 sky130_fd_sc_hd__a32o_1 _22076_ (.A1(_11761_),
    .A2(_11762_),
    .A3(_11765_),
    .B1(_11768_),
    .B2(_10546_),
    .X(_12093_));
 sky130_fd_sc_hd__nand3_4 _22077_ (.A(_12090_),
    .B(_12091_),
    .C(_12093_),
    .Y(_12094_));
 sky130_fd_sc_hd__a32oi_2 _22078_ (.A1(net133),
    .A2(_12085_),
    .A3(_12086_),
    .B1(_11768_),
    .B2(_11773_),
    .Y(_12095_));
 sky130_fd_sc_hd__and3_1 _22079_ (.A(_12087_),
    .B(_12092_),
    .C(_12088_),
    .X(_12096_));
 sky130_fd_sc_hd__nand3_2 _22080_ (.A(_12087_),
    .B(_12092_),
    .C(_12088_),
    .Y(_12097_));
 sky130_fd_sc_hd__a21oi_4 _22081_ (.A1(_11739_),
    .A2(_11741_),
    .B1(_11042_),
    .Y(_12098_));
 sky130_fd_sc_hd__a21o_4 _22082_ (.A1(_11739_),
    .A2(_11741_),
    .B1(_11042_),
    .X(_12099_));
 sky130_fd_sc_hd__o211ai_2 _22083_ (.A1(_11742_),
    .A2(_11042_),
    .B1(_12097_),
    .C1(_12094_),
    .Y(_12101_));
 sky130_fd_sc_hd__a21o_1 _22084_ (.A1(_12094_),
    .A2(_12097_),
    .B1(_12099_),
    .X(_12102_));
 sky130_fd_sc_hd__o2bb2ai_1 _22085_ (.A1_N(_12094_),
    .A2_N(_12097_),
    .B1(_11042_),
    .B2(_11742_),
    .Y(_12103_));
 sky130_fd_sc_hd__o2111ai_4 _22086_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net142),
    .C1(_12094_),
    .D1(_12097_),
    .Y(_12104_));
 sky130_fd_sc_hd__nand3_4 _22087_ (.A(_12102_),
    .B(_12071_),
    .C(_12101_),
    .Y(_12105_));
 sky130_fd_sc_hd__o211ai_4 _22088_ (.A1(_11778_),
    .A2(_12070_),
    .B1(_12103_),
    .C1(_12104_),
    .Y(_12106_));
 sky130_fd_sc_hd__nand2_1 _22089_ (.A(_12105_),
    .B(_12106_),
    .Y(_12107_));
 sky130_fd_sc_hd__o211ai_2 _22090_ (.A1(_12065_),
    .A2(_12060_),
    .B1(_12064_),
    .C1(_12107_),
    .Y(_12108_));
 sky130_fd_sc_hd__nand3_2 _22091_ (.A(_12066_),
    .B(_12068_),
    .C(_12106_),
    .Y(_12109_));
 sky130_fd_sc_hd__nand4_2 _22092_ (.A(_12066_),
    .B(_12068_),
    .C(_12105_),
    .D(_12106_),
    .Y(_12110_));
 sky130_fd_sc_hd__nand2_2 _22093_ (.A(_12069_),
    .B(_12107_),
    .Y(_12112_));
 sky130_fd_sc_hd__o2111ai_4 _22094_ (.A1(_12060_),
    .A2(_12065_),
    .B1(_12105_),
    .C1(_12106_),
    .D1(_12064_),
    .Y(_12113_));
 sky130_fd_sc_hd__a21oi_4 _22095_ (.A1(_12112_),
    .A2(_12113_),
    .B1(_12011_),
    .Y(_12114_));
 sky130_fd_sc_hd__nand3_4 _22096_ (.A(_12010_),
    .B(_12108_),
    .C(_12110_),
    .Y(_12115_));
 sky130_fd_sc_hd__nand3_4 _22097_ (.A(_12011_),
    .B(_12112_),
    .C(_12113_),
    .Y(_12116_));
 sky130_fd_sc_hd__and3_1 _22098_ (.A(_11899_),
    .B(_11943_),
    .C(_11945_),
    .X(_12117_));
 sky130_fd_sc_hd__nor2_2 _22099_ (.A(_11900_),
    .B(_12117_),
    .Y(_12118_));
 sky130_fd_sc_hd__a31o_1 _22100_ (.A1(_11899_),
    .A2(_11943_),
    .A3(_11945_),
    .B1(_11900_),
    .X(_12119_));
 sky130_fd_sc_hd__o21ai_4 _22101_ (.A1(_11450_),
    .A2(_11850_),
    .B1(_11849_),
    .Y(_12120_));
 sky130_fd_sc_hd__o21ai_2 _22102_ (.A1(_11845_),
    .A2(_11846_),
    .B1(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__a21oi_2 _22103_ (.A1(_11924_),
    .A2(_11932_),
    .B1(_11926_),
    .Y(_12123_));
 sky130_fd_sc_hd__and3_1 _22104_ (.A(_04102_),
    .B(net14),
    .C(net42),
    .X(_12124_));
 sky130_fd_sc_hd__and3_1 _22105_ (.A(net182),
    .B(net179),
    .C(_04895_),
    .X(_12125_));
 sky130_fd_sc_hd__a31oi_4 _22106_ (.A1(net182),
    .A2(net179),
    .A3(_04895_),
    .B1(_12124_),
    .Y(_12126_));
 sky130_fd_sc_hd__a31o_1 _22107_ (.A1(net182),
    .A2(net179),
    .A3(_04895_),
    .B1(_12124_),
    .X(_12127_));
 sky130_fd_sc_hd__o211ai_4 _22108_ (.A1(net184),
    .A2(_05551_),
    .B1(net279),
    .C1(net178),
    .Y(_12128_));
 sky130_fd_sc_hd__nor2_1 _22109_ (.A(_04146_),
    .B(_04483_),
    .Y(_12129_));
 sky130_fd_sc_hd__or3b_2 _22110_ (.A(net42),
    .B(_04146_),
    .C_N(net41),
    .X(_12130_));
 sky130_fd_sc_hd__a31oi_4 _22111_ (.A1(net178),
    .A2(net177),
    .A3(net279),
    .B1(_12129_),
    .Y(_12131_));
 sky130_fd_sc_hd__nor2_2 _22112_ (.A(_04157_),
    .B(_04270_),
    .Y(_12132_));
 sky130_fd_sc_hd__o311a_1 _22113_ (.A1(net7),
    .A2(net248),
    .A3(_05927_),
    .B1(_04267_),
    .C1(_05933_),
    .X(_12134_));
 sky130_fd_sc_hd__a31oi_4 _22114_ (.A1(_05933_),
    .A2(_04267_),
    .A3(net174),
    .B1(_12132_),
    .Y(_12135_));
 sky130_fd_sc_hd__nand2_2 _22115_ (.A(_12131_),
    .B(_12135_),
    .Y(_12136_));
 sky130_fd_sc_hd__a21oi_1 _22116_ (.A1(_12128_),
    .A2(_12130_),
    .B1(_12135_),
    .Y(_12137_));
 sky130_fd_sc_hd__o2bb2ai_4 _22117_ (.A1_N(_12128_),
    .A2_N(_12130_),
    .B1(_12132_),
    .B2(_12134_),
    .Y(_12138_));
 sky130_fd_sc_hd__nand2_1 _22118_ (.A(_12136_),
    .B(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__nand3_1 _22119_ (.A(_12126_),
    .B(_12131_),
    .C(_12135_),
    .Y(_12140_));
 sky130_fd_sc_hd__o21ai_1 _22120_ (.A1(_12131_),
    .A2(_12135_),
    .B1(_12126_),
    .Y(_12141_));
 sky130_fd_sc_hd__o2bb2ai_1 _22121_ (.A1_N(_12131_),
    .A2_N(_12135_),
    .B1(_12124_),
    .B2(_12125_),
    .Y(_12142_));
 sky130_fd_sc_hd__a21oi_1 _22122_ (.A1(_12127_),
    .A2(_12136_),
    .B1(_12137_),
    .Y(_12143_));
 sky130_fd_sc_hd__o211ai_4 _22123_ (.A1(_12131_),
    .A2(_12135_),
    .B1(_12140_),
    .C1(_12142_),
    .Y(_12145_));
 sky130_fd_sc_hd__a211o_1 _22124_ (.A1(_12128_),
    .A2(_12130_),
    .B1(_12135_),
    .C1(_12126_),
    .X(_12146_));
 sky130_fd_sc_hd__o221a_1 _22125_ (.A1(_12124_),
    .A2(_12125_),
    .B1(_12131_),
    .B2(_12135_),
    .C1(_12136_),
    .X(_12147_));
 sky130_fd_sc_hd__a311o_1 _22126_ (.A1(_12128_),
    .A2(_12135_),
    .A3(_12130_),
    .B1(_12126_),
    .C1(_12137_),
    .X(_12148_));
 sky130_fd_sc_hd__a21oi_1 _22127_ (.A1(_12136_),
    .A2(_12138_),
    .B1(_12127_),
    .Y(_12149_));
 sky130_fd_sc_hd__o2111ai_4 _22128_ (.A1(_12138_),
    .A2(_12126_),
    .B1(_11934_),
    .C1(_11927_),
    .D1(_12145_),
    .Y(_12150_));
 sky130_fd_sc_hd__a32o_1 _22129_ (.A1(net217),
    .A2(net186),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net10),
    .X(_12151_));
 sky130_fd_sc_hd__o311a_1 _22130_ (.A1(net7),
    .A2(net248),
    .A3(_04787_),
    .B1(net276),
    .C1(net213),
    .X(_12152_));
 sky130_fd_sc_hd__o211ai_2 _22131_ (.A1(net231),
    .A2(_04787_),
    .B1(net276),
    .C1(net213),
    .Y(_12153_));
 sky130_fd_sc_hd__nor2_1 _22132_ (.A(_04091_),
    .B(_05229_),
    .Y(_12154_));
 sky130_fd_sc_hd__or3_1 _22133_ (.A(net46),
    .B(_04124_),
    .C(_04091_),
    .X(_12156_));
 sky130_fd_sc_hd__a31o_1 _22134_ (.A1(net184),
    .A2(net213),
    .A3(net276),
    .B1(_12154_),
    .X(_12157_));
 sky130_fd_sc_hd__o211ai_4 _22135_ (.A1(_04787_),
    .A2(net208),
    .B1(net242),
    .C1(net210),
    .Y(_12158_));
 sky130_fd_sc_hd__or3_1 _22136_ (.A(net45),
    .B(_04113_),
    .C(_04102_),
    .X(_12159_));
 sky130_fd_sc_hd__o21ai_2 _22137_ (.A1(_04113_),
    .A2(_04989_),
    .B1(_12158_),
    .Y(_12160_));
 sky130_fd_sc_hd__o311a_1 _22138_ (.A1(_04091_),
    .A2(net46),
    .A3(_04124_),
    .B1(_12159_),
    .C1(_12153_),
    .X(_12161_));
 sky130_fd_sc_hd__a22oi_2 _22139_ (.A1(_12153_),
    .A2(_12156_),
    .B1(_12158_),
    .B2(_12159_),
    .Y(_12162_));
 sky130_fd_sc_hd__a22o_1 _22140_ (.A1(_12153_),
    .A2(_12156_),
    .B1(_12158_),
    .B2(_12159_),
    .X(_12163_));
 sky130_fd_sc_hd__nand3b_1 _22141_ (.A_N(_12151_),
    .B(_12161_),
    .C(_12158_),
    .Y(_12164_));
 sky130_fd_sc_hd__o21ai_1 _22142_ (.A1(_12157_),
    .A2(_12160_),
    .B1(_12151_),
    .Y(_12165_));
 sky130_fd_sc_hd__o32ai_4 _22143_ (.A1(_12152_),
    .A2(_12154_),
    .A3(_12160_),
    .B1(_12151_),
    .B2(_12162_),
    .Y(_12167_));
 sky130_fd_sc_hd__and3_1 _22144_ (.A(_12151_),
    .B(_12157_),
    .C(_12160_),
    .X(_12168_));
 sky130_fd_sc_hd__a21oi_1 _22145_ (.A1(_12164_),
    .A2(_12167_),
    .B1(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__a31o_2 _22146_ (.A1(_12163_),
    .A2(_12164_),
    .A3(_12165_),
    .B1(_12168_),
    .X(_12170_));
 sky130_fd_sc_hd__o2111ai_1 _22147_ (.A1(_12138_),
    .A2(_12126_),
    .B1(_12123_),
    .C1(_12145_),
    .D1(_12169_),
    .Y(_12171_));
 sky130_fd_sc_hd__a21oi_1 _22148_ (.A1(_12139_),
    .A2(_12126_),
    .B1(_12123_),
    .Y(_12172_));
 sky130_fd_sc_hd__a22o_1 _22149_ (.A1(_11927_),
    .A2(_11934_),
    .B1(_12145_),
    .B2(_12146_),
    .X(_12173_));
 sky130_fd_sc_hd__o31ai_2 _22150_ (.A1(_12123_),
    .A2(_12147_),
    .A3(_12149_),
    .B1(_12169_),
    .Y(_12174_));
 sky130_fd_sc_hd__nand2_1 _22151_ (.A(_12150_),
    .B(_12170_),
    .Y(_12175_));
 sky130_fd_sc_hd__a22oi_4 _22152_ (.A1(_12172_),
    .A2(_12148_),
    .B1(_12150_),
    .B2(_12170_),
    .Y(_12176_));
 sky130_fd_sc_hd__o311a_2 _22153_ (.A1(_12123_),
    .A2(_12147_),
    .A3(_12149_),
    .B1(_12171_),
    .C1(_12175_),
    .X(_12178_));
 sky130_fd_sc_hd__and3_2 _22154_ (.A(_12172_),
    .B(_12170_),
    .C(_12148_),
    .X(_12179_));
 sky130_fd_sc_hd__and3_2 _22155_ (.A(_12150_),
    .B(_12170_),
    .C(_12173_),
    .X(_12180_));
 sky130_fd_sc_hd__a21oi_2 _22156_ (.A1(_12150_),
    .A2(_12173_),
    .B1(_12170_),
    .Y(_12181_));
 sky130_fd_sc_hd__o2bb2a_1 _22157_ (.A1_N(_12171_),
    .A2_N(_12176_),
    .B1(_12173_),
    .B2(_12169_),
    .X(_12182_));
 sky130_fd_sc_hd__a311oi_4 _22158_ (.A1(_11466_),
    .A2(_11886_),
    .A3(_11887_),
    .B1(_11388_),
    .C1(_11385_),
    .Y(_12183_));
 sky130_fd_sc_hd__nor2_1 _22159_ (.A(_11875_),
    .B(_11889_),
    .Y(_12184_));
 sky130_fd_sc_hd__a21o_1 _22160_ (.A1(_11884_),
    .A2(_11885_),
    .B1(_11880_),
    .X(_12185_));
 sky130_fd_sc_hd__nor2_1 _22161_ (.A(_04179_),
    .B(_03737_),
    .Y(_12186_));
 sky130_fd_sc_hd__a31oi_4 _22162_ (.A1(net198),
    .A2(net172),
    .A3(_03704_),
    .B1(_12186_),
    .Y(_12187_));
 sky130_fd_sc_hd__o211ai_2 _22163_ (.A1(net174),
    .A2(_06759_),
    .B1(_02858_),
    .C1(net193),
    .Y(_12189_));
 sky130_fd_sc_hd__or3b_2 _22164_ (.A(net38),
    .B(_04201_),
    .C_N(net37),
    .X(_12190_));
 sky130_fd_sc_hd__a21oi_4 _22165_ (.A1(_12189_),
    .A2(_12190_),
    .B1(_12187_),
    .Y(_12191_));
 sky130_fd_sc_hd__a21o_1 _22166_ (.A1(_12189_),
    .A2(_12190_),
    .B1(_12187_),
    .X(_12192_));
 sky130_fd_sc_hd__o311a_1 _22167_ (.A1(_02869_),
    .A2(_06756_),
    .A3(net189),
    .B1(_12190_),
    .C1(_12187_),
    .X(_12193_));
 sky130_fd_sc_hd__o221ai_4 _22168_ (.A1(_04201_),
    .A2(_02891_),
    .B1(_06764_),
    .B2(_02869_),
    .C1(_12187_),
    .Y(_12194_));
 sky130_fd_sc_hd__a32o_1 _22169_ (.A1(net201),
    .A2(net173),
    .A3(net281),
    .B1(_04217_),
    .B2(net17),
    .X(_12195_));
 sky130_fd_sc_hd__o21bai_4 _22170_ (.A1(_12191_),
    .A2(_12193_),
    .B1_N(_12195_),
    .Y(_12196_));
 sky130_fd_sc_hd__and3_4 _22171_ (.A(_12192_),
    .B(_12194_),
    .C(_12195_),
    .X(_12197_));
 sky130_fd_sc_hd__nand3_2 _22172_ (.A(_12192_),
    .B(_12194_),
    .C(_12195_),
    .Y(_12198_));
 sky130_fd_sc_hd__o221a_1 _22173_ (.A1(_04201_),
    .A2(_01326_),
    .B1(_06764_),
    .B2(_01304_),
    .C1(_11832_),
    .X(_12200_));
 sky130_fd_sc_hd__a41oi_4 _22174_ (.A1(_11823_),
    .A2(_11824_),
    .A3(_11828_),
    .A4(_11830_),
    .B1(_11821_),
    .Y(_12201_));
 sky130_fd_sc_hd__a21oi_1 _22175_ (.A1(_11822_),
    .A2(_11834_),
    .B1(_11831_),
    .Y(_12202_));
 sky130_fd_sc_hd__a21boi_1 _22176_ (.A1(_12196_),
    .A2(_12198_),
    .B1_N(_12202_),
    .Y(_12203_));
 sky130_fd_sc_hd__o2bb2ai_4 _22177_ (.A1_N(_12196_),
    .A2_N(_12198_),
    .B1(_12200_),
    .B2(_11833_),
    .Y(_12204_));
 sky130_fd_sc_hd__o21ai_4 _22178_ (.A1(_11831_),
    .A2(_12201_),
    .B1(_12196_),
    .Y(_12205_));
 sky130_fd_sc_hd__o211a_1 _22179_ (.A1(_11831_),
    .A2(_12201_),
    .B1(_12198_),
    .C1(_12196_),
    .X(_12206_));
 sky130_fd_sc_hd__o211ai_1 _22180_ (.A1(_11831_),
    .A2(_12201_),
    .B1(_12198_),
    .C1(_12196_),
    .Y(_12207_));
 sky130_fd_sc_hd__o221a_2 _22181_ (.A1(_11880_),
    .A2(_11888_),
    .B1(_12197_),
    .B2(_12205_),
    .C1(_12204_),
    .X(_12208_));
 sky130_fd_sc_hd__o221ai_4 _22182_ (.A1(_11880_),
    .A2(_11888_),
    .B1(_12197_),
    .B2(_12205_),
    .C1(_12204_),
    .Y(_12209_));
 sky130_fd_sc_hd__a21oi_2 _22183_ (.A1(_12204_),
    .A2(_12207_),
    .B1(_12185_),
    .Y(_12211_));
 sky130_fd_sc_hd__o21bai_2 _22184_ (.A1(_12203_),
    .A2(_12206_),
    .B1_N(_12185_),
    .Y(_12212_));
 sky130_fd_sc_hd__o211a_2 _22185_ (.A1(_11891_),
    .A2(_12184_),
    .B1(_12209_),
    .C1(_12212_),
    .X(_12213_));
 sky130_fd_sc_hd__o211ai_4 _22186_ (.A1(_11891_),
    .A2(_12184_),
    .B1(_12209_),
    .C1(_12212_),
    .Y(_12214_));
 sky130_fd_sc_hd__o22a_2 _22187_ (.A1(_11889_),
    .A2(_12183_),
    .B1(_12208_),
    .B2(_12211_),
    .X(_12215_));
 sky130_fd_sc_hd__o22ai_4 _22188_ (.A1(_11889_),
    .A2(_12183_),
    .B1(_12208_),
    .B2(_12211_),
    .Y(_12216_));
 sky130_fd_sc_hd__o41a_1 _22189_ (.A1(_11889_),
    .A2(_12183_),
    .A3(_12208_),
    .A4(_12211_),
    .B1(_12182_),
    .X(_12217_));
 sky130_fd_sc_hd__o21a_1 _22190_ (.A1(_12178_),
    .A2(_12179_),
    .B1(_12216_),
    .X(_12218_));
 sky130_fd_sc_hd__o31a_1 _22191_ (.A1(_12178_),
    .A2(_12179_),
    .A3(_12213_),
    .B1(_12216_),
    .X(_12219_));
 sky130_fd_sc_hd__o211ai_2 _22192_ (.A1(_12180_),
    .A2(_12181_),
    .B1(_12214_),
    .C1(_12216_),
    .Y(_12220_));
 sky130_fd_sc_hd__o22ai_2 _22193_ (.A1(_12178_),
    .A2(_12179_),
    .B1(_12213_),
    .B2(_12215_),
    .Y(_12222_));
 sky130_fd_sc_hd__a2bb2oi_4 _22194_ (.A1_N(_12180_),
    .A2_N(_12181_),
    .B1(_12214_),
    .B2(_12216_),
    .Y(_12223_));
 sky130_fd_sc_hd__o22ai_2 _22195_ (.A1(_12180_),
    .A2(_12181_),
    .B1(_12213_),
    .B2(_12215_),
    .Y(_12224_));
 sky130_fd_sc_hd__o211a_1 _22196_ (.A1(_12178_),
    .A2(_12179_),
    .B1(_12214_),
    .C1(_12216_),
    .X(_12225_));
 sky130_fd_sc_hd__o211ai_4 _22197_ (.A1(_12178_),
    .A2(_12179_),
    .B1(_12214_),
    .C1(_12216_),
    .Y(_12226_));
 sky130_fd_sc_hd__o211ai_4 _22198_ (.A1(_11845_),
    .A2(_11846_),
    .B1(_12120_),
    .C1(_12226_),
    .Y(_12227_));
 sky130_fd_sc_hd__nand4_4 _22199_ (.A(_11847_),
    .B(_12120_),
    .C(_12224_),
    .D(_12226_),
    .Y(_12228_));
 sky130_fd_sc_hd__nand3_4 _22200_ (.A(_12121_),
    .B(_12220_),
    .C(_12222_),
    .Y(_12229_));
 sky130_fd_sc_hd__o211a_1 _22201_ (.A1(_12223_),
    .A2(_12227_),
    .B1(_12118_),
    .C1(_12229_),
    .X(_12230_));
 sky130_fd_sc_hd__o211ai_2 _22202_ (.A1(_12223_),
    .A2(_12227_),
    .B1(_12118_),
    .C1(_12229_),
    .Y(_12231_));
 sky130_fd_sc_hd__a21oi_2 _22203_ (.A1(_12228_),
    .A2(_12229_),
    .B1(_12118_),
    .Y(_12233_));
 sky130_fd_sc_hd__a21o_1 _22204_ (.A1(_12228_),
    .A2(_12229_),
    .B1(_12118_),
    .X(_12234_));
 sky130_fd_sc_hd__nor2_1 _22205_ (.A(_12119_),
    .B(_12228_),
    .Y(_12235_));
 sky130_fd_sc_hd__o211a_1 _22206_ (.A1(_12223_),
    .A2(_12225_),
    .B1(_12119_),
    .C1(_12121_),
    .X(_12236_));
 sky130_fd_sc_hd__o22ai_4 _22207_ (.A1(_11900_),
    .A2(_12117_),
    .B1(_12223_),
    .B2(_12227_),
    .Y(_12237_));
 sky130_fd_sc_hd__o2bb2ai_2 _22208_ (.A1_N(_12118_),
    .A2_N(_12229_),
    .B1(_12227_),
    .B2(_12223_),
    .Y(_12238_));
 sky130_fd_sc_hd__a21oi_1 _22209_ (.A1(_12229_),
    .A2(_12237_),
    .B1(_12236_),
    .Y(_12239_));
 sky130_fd_sc_hd__o22ai_2 _22210_ (.A1(_12119_),
    .A2(_12228_),
    .B1(_12236_),
    .B2(_12238_),
    .Y(_12240_));
 sky130_fd_sc_hd__o2bb2ai_2 _22211_ (.A1_N(_12115_),
    .A2_N(_12116_),
    .B1(_12230_),
    .B2(_12233_),
    .Y(_12241_));
 sky130_fd_sc_hd__nand3_1 _22212_ (.A(_12116_),
    .B(_12231_),
    .C(_12234_),
    .Y(_12242_));
 sky130_fd_sc_hd__nand4_2 _22213_ (.A(_12115_),
    .B(_12116_),
    .C(_12231_),
    .D(_12234_),
    .Y(_12244_));
 sky130_fd_sc_hd__o211ai_4 _22214_ (.A1(_12230_),
    .A2(_12233_),
    .B1(_12115_),
    .C1(_12116_),
    .Y(_12245_));
 sky130_fd_sc_hd__o2bb2ai_4 _22215_ (.A1_N(_12115_),
    .A2_N(_12116_),
    .B1(_12235_),
    .B2(_12239_),
    .Y(_12246_));
 sky130_fd_sc_hd__nand2_1 _22216_ (.A(_12241_),
    .B(_12244_),
    .Y(_12247_));
 sky130_fd_sc_hd__and3_1 _22217_ (.A(_12007_),
    .B(_12241_),
    .C(_12244_),
    .X(_12248_));
 sky130_fd_sc_hd__nand3_2 _22218_ (.A(_12007_),
    .B(_12241_),
    .C(_12244_),
    .Y(_12249_));
 sky130_fd_sc_hd__a21oi_1 _22219_ (.A1(_12241_),
    .A2(_12244_),
    .B1(_12007_),
    .Y(_12250_));
 sky130_fd_sc_hd__o211ai_4 _22220_ (.A1(_11869_),
    .A2(_12006_),
    .B1(_12245_),
    .C1(_12246_),
    .Y(_12251_));
 sky130_fd_sc_hd__o21ai_2 _22221_ (.A1(_11403_),
    .A2(_11956_),
    .B1(_11955_),
    .Y(_12252_));
 sky130_fd_sc_hd__a41oi_4 _22222_ (.A1(_11483_),
    .A2(_11488_),
    .A3(_11949_),
    .A4(_11950_),
    .B1(_11959_),
    .Y(_12253_));
 sky130_fd_sc_hd__o2bb2a_1 _22223_ (.A1_N(_09709_),
    .A2_N(_08005_),
    .B1(_08007_),
    .B2(_03960_),
    .X(_12254_));
 sky130_fd_sc_hd__a32o_2 _22224_ (.A1(net255),
    .A2(_09698_),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net2),
    .X(_12255_));
 sky130_fd_sc_hd__a32o_1 _22225_ (.A1(_11354_),
    .A2(net253),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net3),
    .X(_12256_));
 sky130_fd_sc_hd__o21ai_2 _22226_ (.A1(_11615_),
    .A2(_11622_),
    .B1(_11625_),
    .Y(_12257_));
 sky130_fd_sc_hd__and3_1 _22227_ (.A(_04234_),
    .B(net52),
    .C(net4),
    .X(_12258_));
 sky130_fd_sc_hd__a21oi_1 _22228_ (.A1(_13010_),
    .A2(net239),
    .B1(_12258_),
    .Y(_12259_));
 sky130_fd_sc_hd__a31o_1 _22229_ (.A1(net234),
    .A2(net251),
    .A3(net239),
    .B1(_12258_),
    .X(_12260_));
 sky130_fd_sc_hd__or3_1 _22230_ (.A(net51),
    .B(_04190_),
    .C(_04026_),
    .X(_12261_));
 sky130_fd_sc_hd__o211ai_4 _22231_ (.A1(net253),
    .A2(_02442_),
    .B1(net240),
    .C1(_02421_),
    .Y(_12262_));
 sky130_fd_sc_hd__or3b_2 _22232_ (.A(_04015_),
    .B(net52),
    .C_N(net51),
    .X(_12263_));
 sky130_fd_sc_hd__o211ai_4 _22233_ (.A1(net253),
    .A2(_00646_),
    .B1(net269),
    .C1(_00625_),
    .Y(_12265_));
 sky130_fd_sc_hd__a22oi_2 _22234_ (.A1(_12261_),
    .A2(_12262_),
    .B1(_12263_),
    .B2(_12265_),
    .Y(_12266_));
 sky130_fd_sc_hd__a22o_1 _22235_ (.A1(_12261_),
    .A2(_12262_),
    .B1(_12263_),
    .B2(_12265_),
    .X(_12267_));
 sky130_fd_sc_hd__o2111a_1 _22236_ (.A1(_04026_),
    .A2(_06866_),
    .B1(_12262_),
    .C1(_12263_),
    .D1(_12265_),
    .X(_12268_));
 sky130_fd_sc_hd__o2111ai_2 _22237_ (.A1(_04026_),
    .A2(_06866_),
    .B1(_12262_),
    .C1(_12263_),
    .D1(_12265_),
    .Y(_12269_));
 sky130_fd_sc_hd__nand3_1 _22238_ (.A(_12260_),
    .B(_12267_),
    .C(_12269_),
    .Y(_12270_));
 sky130_fd_sc_hd__o21ai_1 _22239_ (.A1(_12266_),
    .A2(_12268_),
    .B1(_12259_),
    .Y(_12271_));
 sky130_fd_sc_hd__nand3_1 _22240_ (.A(_12267_),
    .B(_12269_),
    .C(_12259_),
    .Y(_12272_));
 sky130_fd_sc_hd__o21ai_2 _22241_ (.A1(_12266_),
    .A2(_12268_),
    .B1(_12260_),
    .Y(_12273_));
 sky130_fd_sc_hd__o2111a_1 _22242_ (.A1(_11615_),
    .A2(_11622_),
    .B1(_11625_),
    .C1(_12272_),
    .D1(_12273_),
    .X(_12274_));
 sky130_fd_sc_hd__o2111ai_4 _22243_ (.A1(_11615_),
    .A2(_11622_),
    .B1(_11625_),
    .C1(_12272_),
    .D1(_12273_),
    .Y(_12276_));
 sky130_fd_sc_hd__nand3_2 _22244_ (.A(_12271_),
    .B(_12257_),
    .C(_12270_),
    .Y(_12277_));
 sky130_fd_sc_hd__a21o_1 _22245_ (.A1(_12276_),
    .A2(_12277_),
    .B1(_12256_),
    .X(_12278_));
 sky130_fd_sc_hd__nand3_1 _22246_ (.A(_12256_),
    .B(_12276_),
    .C(_12277_),
    .Y(_12279_));
 sky130_fd_sc_hd__nand3b_2 _22247_ (.A_N(_12256_),
    .B(_12276_),
    .C(_12277_),
    .Y(_12280_));
 sky130_fd_sc_hd__a21bo_1 _22248_ (.A1(_12276_),
    .A2(_12277_),
    .B1_N(_12256_),
    .X(_12281_));
 sky130_fd_sc_hd__nand2_1 _22249_ (.A(_11633_),
    .B(_11613_),
    .Y(_12282_));
 sky130_fd_sc_hd__nand4_4 _22250_ (.A(_11631_),
    .B(_12278_),
    .C(_12279_),
    .D(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__inv_2 _22251_ (.A(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__o2111a_1 _22252_ (.A1(_11613_),
    .A2(_11630_),
    .B1(_11633_),
    .C1(_12280_),
    .D1(_12281_),
    .X(_12285_));
 sky130_fd_sc_hd__o2111ai_4 _22253_ (.A1(_11613_),
    .A2(_11630_),
    .B1(_11633_),
    .C1(_12280_),
    .D1(_12281_),
    .Y(_12287_));
 sky130_fd_sc_hd__a21oi_1 _22254_ (.A1(_12283_),
    .A2(_12287_),
    .B1(_12255_),
    .Y(_12288_));
 sky130_fd_sc_hd__a21o_1 _22255_ (.A1(_12283_),
    .A2(_12287_),
    .B1(_12255_),
    .X(_12289_));
 sky130_fd_sc_hd__and3_1 _22256_ (.A(_12255_),
    .B(_12283_),
    .C(_12287_),
    .X(_12290_));
 sky130_fd_sc_hd__nand3_1 _22257_ (.A(_12255_),
    .B(_12283_),
    .C(_12287_),
    .Y(_12291_));
 sky130_fd_sc_hd__nor2_1 _22258_ (.A(_12288_),
    .B(_12290_),
    .Y(_12292_));
 sky130_fd_sc_hd__nand2_1 _22259_ (.A(_12289_),
    .B(_12291_),
    .Y(_12293_));
 sky130_fd_sc_hd__and3_1 _22260_ (.A(_11280_),
    .B(_11284_),
    .C(_11681_),
    .X(_12294_));
 sky130_fd_sc_hd__o31a_1 _22261_ (.A1(_11279_),
    .A2(_11283_),
    .A3(_11680_),
    .B1(_11684_),
    .X(_12295_));
 sky130_fd_sc_hd__o311ai_4 _22262_ (.A1(_11916_),
    .A2(_11933_),
    .A3(_11935_),
    .B1(_11913_),
    .C1(_11912_),
    .Y(_12296_));
 sky130_fd_sc_hd__a22oi_2 _22263_ (.A1(_11934_),
    .A2(_11937_),
    .B1(_11941_),
    .B2(_11915_),
    .Y(_12298_));
 sky130_fd_sc_hd__a32o_1 _22264_ (.A1(_03952_),
    .A2(net231),
    .A3(net273),
    .B1(_06326_),
    .B2(net7),
    .X(_12299_));
 sky130_fd_sc_hd__nand3_2 _22265_ (.A(_04409_),
    .B(net221),
    .C(_05762_),
    .Y(_12300_));
 sky130_fd_sc_hd__or3b_2 _22266_ (.A(_04069_),
    .B(net48),
    .C_N(net47),
    .X(_12301_));
 sky130_fd_sc_hd__nor2_1 _22267_ (.A(_04059_),
    .B(_06030_),
    .Y(_12302_));
 sky130_fd_sc_hd__a31oi_4 _22268_ (.A1(net229),
    .A2(net227),
    .A3(net274),
    .B1(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__a21oi_4 _22269_ (.A1(_12300_),
    .A2(_12301_),
    .B1(_12303_),
    .Y(_12304_));
 sky130_fd_sc_hd__a21o_1 _22270_ (.A1(_12300_),
    .A2(_12301_),
    .B1(_12303_),
    .X(_12305_));
 sky130_fd_sc_hd__o211a_1 _22271_ (.A1(_04069_),
    .A2(_05766_),
    .B1(_12300_),
    .C1(_12303_),
    .X(_12306_));
 sky130_fd_sc_hd__o221ai_4 _22272_ (.A1(net187),
    .A2(_05763_),
    .B1(_05766_),
    .B2(_04069_),
    .C1(_12303_),
    .Y(_12307_));
 sky130_fd_sc_hd__o21bai_4 _22273_ (.A1(_12304_),
    .A2(_12306_),
    .B1_N(_12299_),
    .Y(_12309_));
 sky130_fd_sc_hd__and3_1 _22274_ (.A(_12299_),
    .B(_12305_),
    .C(_12307_),
    .X(_12310_));
 sky130_fd_sc_hd__nand3_4 _22275_ (.A(_12299_),
    .B(_12305_),
    .C(_12307_),
    .Y(_12311_));
 sky130_fd_sc_hd__o21a_1 _22276_ (.A1(_11907_),
    .A2(_11908_),
    .B1(_11905_),
    .X(_12312_));
 sky130_fd_sc_hd__a21oi_2 _22277_ (.A1(_11907_),
    .A2(_11908_),
    .B1(_11905_),
    .Y(_12313_));
 sky130_fd_sc_hd__o2bb2ai_1 _22278_ (.A1_N(_11907_),
    .A2_N(_11908_),
    .B1(_11902_),
    .B2(_11904_),
    .Y(_12314_));
 sky130_fd_sc_hd__o21ai_1 _22279_ (.A1(_11907_),
    .A2(_11908_),
    .B1(_12314_),
    .Y(_12315_));
 sky130_fd_sc_hd__a21oi_4 _22280_ (.A1(_12309_),
    .A2(_12311_),
    .B1(_12315_),
    .Y(_12316_));
 sky130_fd_sc_hd__o2bb2ai_1 _22281_ (.A1_N(_12309_),
    .A2_N(_12311_),
    .B1(_12312_),
    .B2(_11910_),
    .Y(_12317_));
 sky130_fd_sc_hd__o211a_1 _22282_ (.A1(_11909_),
    .A2(_12313_),
    .B1(_12311_),
    .C1(_12309_),
    .X(_12318_));
 sky130_fd_sc_hd__o211ai_4 _22283_ (.A1(_11909_),
    .A2(_12313_),
    .B1(_12311_),
    .C1(_12309_),
    .Y(_12320_));
 sky130_fd_sc_hd__a21oi_1 _22284_ (.A1(_12317_),
    .A2(_12320_),
    .B1(_11677_),
    .Y(_12321_));
 sky130_fd_sc_hd__o22ai_4 _22285_ (.A1(_11671_),
    .A2(_11676_),
    .B1(_12316_),
    .B2(_12318_),
    .Y(_12322_));
 sky130_fd_sc_hd__nand2_1 _22286_ (.A(_12320_),
    .B(_11677_),
    .Y(_12323_));
 sky130_fd_sc_hd__and3_1 _22287_ (.A(_12317_),
    .B(_12320_),
    .C(_11677_),
    .X(_12324_));
 sky130_fd_sc_hd__nand3_2 _22288_ (.A(_12317_),
    .B(_12320_),
    .C(_11677_),
    .Y(_12325_));
 sky130_fd_sc_hd__o21ai_1 _22289_ (.A1(_12316_),
    .A2(_12323_),
    .B1(_12322_),
    .Y(_12326_));
 sky130_fd_sc_hd__o2111a_2 _22290_ (.A1(_12316_),
    .A2(_12323_),
    .B1(_12322_),
    .C1(_11941_),
    .D1(_12296_),
    .X(_12327_));
 sky130_fd_sc_hd__o2111ai_4 _22291_ (.A1(_12316_),
    .A2(_12323_),
    .B1(_12322_),
    .C1(_11941_),
    .D1(_12296_),
    .Y(_12328_));
 sky130_fd_sc_hd__a221oi_2 _22292_ (.A1(_11915_),
    .A2(_11941_),
    .B1(_12322_),
    .B2(_12325_),
    .C1(_11939_),
    .Y(_12329_));
 sky130_fd_sc_hd__o21ai_2 _22293_ (.A1(_12321_),
    .A2(_12324_),
    .B1(_12298_),
    .Y(_12331_));
 sky130_fd_sc_hd__a21oi_1 _22294_ (.A1(_12328_),
    .A2(_12331_),
    .B1(_12295_),
    .Y(_12332_));
 sky130_fd_sc_hd__o22ai_2 _22295_ (.A1(_11682_),
    .A2(_12294_),
    .B1(_12327_),
    .B2(_12329_),
    .Y(_12333_));
 sky130_fd_sc_hd__a2bb2oi_1 _22296_ (.A1_N(_11680_),
    .A2_N(_11685_),
    .B1(_12298_),
    .B2(_12326_),
    .Y(_12334_));
 sky130_fd_sc_hd__o211ai_2 _22297_ (.A1(_11680_),
    .A2(_11685_),
    .B1(_12328_),
    .C1(_12331_),
    .Y(_12335_));
 sky130_fd_sc_hd__o22ai_1 _22298_ (.A1(_11680_),
    .A2(_11685_),
    .B1(_12327_),
    .B2(_12329_),
    .Y(_12336_));
 sky130_fd_sc_hd__o211ai_1 _22299_ (.A1(_11682_),
    .A2(_12294_),
    .B1(_12328_),
    .C1(_12331_),
    .Y(_12337_));
 sky130_fd_sc_hd__a32oi_4 _22300_ (.A1(_11656_),
    .A2(_11689_),
    .A3(_11691_),
    .B1(_11696_),
    .B2(_11654_),
    .Y(_12338_));
 sky130_fd_sc_hd__a32o_1 _22301_ (.A1(_11656_),
    .A2(_11689_),
    .A3(_11691_),
    .B1(_11696_),
    .B2(_11654_),
    .X(_12339_));
 sky130_fd_sc_hd__and3_2 _22302_ (.A(_12336_),
    .B(_12337_),
    .C(_12339_),
    .X(_12340_));
 sky130_fd_sc_hd__nand3_2 _22303_ (.A(_12336_),
    .B(_12337_),
    .C(_12339_),
    .Y(_12342_));
 sky130_fd_sc_hd__nand2_1 _22304_ (.A(_12335_),
    .B(_12338_),
    .Y(_12343_));
 sky130_fd_sc_hd__and3_1 _22305_ (.A(_12333_),
    .B(_12335_),
    .C(_12338_),
    .X(_12344_));
 sky130_fd_sc_hd__nand3_2 _22306_ (.A(_12333_),
    .B(_12335_),
    .C(_12338_),
    .Y(_12345_));
 sky130_fd_sc_hd__a31o_1 _22307_ (.A1(_12333_),
    .A2(_12335_),
    .A3(_12338_),
    .B1(_12293_),
    .X(_12346_));
 sky130_fd_sc_hd__o211a_1 _22308_ (.A1(_12332_),
    .A2(_12343_),
    .B1(_12292_),
    .C1(_12342_),
    .X(_12347_));
 sky130_fd_sc_hd__a21oi_2 _22309_ (.A1(_12342_),
    .A2(_12345_),
    .B1(_12292_),
    .Y(_12348_));
 sky130_fd_sc_hd__a22o_1 _22310_ (.A1(_12289_),
    .A2(_12291_),
    .B1(_12342_),
    .B2(_12345_),
    .X(_12349_));
 sky130_fd_sc_hd__o221ai_4 _22311_ (.A1(_11954_),
    .A2(_12253_),
    .B1(_12340_),
    .B2(_12346_),
    .C1(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__o2bb2ai_4 _22312_ (.A1_N(_11953_),
    .A2_N(_12252_),
    .B1(_12347_),
    .B2(_12348_),
    .Y(_12351_));
 sky130_fd_sc_hd__a31o_1 _22313_ (.A1(_11653_),
    .A2(_11698_),
    .A3(_11701_),
    .B1(_11712_),
    .X(_12353_));
 sky130_fd_sc_hd__a2bb2oi_1 _22314_ (.A1_N(_11707_),
    .A2_N(_11712_),
    .B1(_12350_),
    .B2(_12351_),
    .Y(_12354_));
 sky130_fd_sc_hd__a22o_1 _22315_ (.A1(_11708_),
    .A2(_11713_),
    .B1(_12350_),
    .B2(_12351_),
    .X(_12355_));
 sky130_fd_sc_hd__o2111a_1 _22316_ (.A1(_11652_),
    .A2(_11704_),
    .B1(_11713_),
    .C1(_12350_),
    .D1(_12351_),
    .X(_12356_));
 sky130_fd_sc_hd__o2111ai_4 _22317_ (.A1(_11652_),
    .A2(_11704_),
    .B1(_11713_),
    .C1(_12350_),
    .D1(_12351_),
    .Y(_12357_));
 sky130_fd_sc_hd__a21oi_1 _22318_ (.A1(_12350_),
    .A2(_12351_),
    .B1(_12353_),
    .Y(_12358_));
 sky130_fd_sc_hd__and3_1 _22319_ (.A(_12350_),
    .B(_12351_),
    .C(_12353_),
    .X(_12359_));
 sky130_fd_sc_hd__nor2_1 _22320_ (.A(_12354_),
    .B(_12356_),
    .Y(_12360_));
 sky130_fd_sc_hd__a32oi_4 _22321_ (.A1(_12008_),
    .A2(_12245_),
    .A3(_12246_),
    .B1(_12355_),
    .B2(_12357_),
    .Y(_12361_));
 sky130_fd_sc_hd__o211ai_1 _22322_ (.A1(_12354_),
    .A2(_12356_),
    .B1(_12249_),
    .C1(_12251_),
    .Y(_12362_));
 sky130_fd_sc_hd__o2bb2ai_1 _22323_ (.A1_N(_12249_),
    .A2_N(_12251_),
    .B1(_12358_),
    .B2(_12359_),
    .Y(_12364_));
 sky130_fd_sc_hd__nand4_2 _22324_ (.A(_12249_),
    .B(_12251_),
    .C(_12355_),
    .D(_12357_),
    .Y(_12365_));
 sky130_fd_sc_hd__o2bb2ai_1 _22325_ (.A1_N(_12249_),
    .A2_N(_12251_),
    .B1(_12354_),
    .B2(_12356_),
    .Y(_12366_));
 sky130_fd_sc_hd__o22ai_1 _22326_ (.A1(_11966_),
    .A2(_11971_),
    .B1(_11726_),
    .B2(_11968_),
    .Y(_12367_));
 sky130_fd_sc_hd__o2111ai_4 _22327_ (.A1(_11726_),
    .A2(_11968_),
    .B1(_11973_),
    .C1(_12365_),
    .D1(_12366_),
    .Y(_12368_));
 sky130_fd_sc_hd__nand3_2 _22328_ (.A(_12367_),
    .B(_12364_),
    .C(_12362_),
    .Y(_12369_));
 sky130_fd_sc_hd__a21o_1 _22329_ (.A1(_11717_),
    .A2(_11720_),
    .B1(_11718_),
    .X(_12370_));
 sky130_fd_sc_hd__a21o_1 _22330_ (.A1(_12368_),
    .A2(_12369_),
    .B1(_12370_),
    .X(_12371_));
 sky130_fd_sc_hd__o211ai_2 _22331_ (.A1(_11718_),
    .A2(_11724_),
    .B1(_12368_),
    .C1(_12369_),
    .Y(_12372_));
 sky130_fd_sc_hd__nand4_1 _22332_ (.A(_11719_),
    .B(_11725_),
    .C(_12368_),
    .D(_12369_),
    .Y(_12373_));
 sky130_fd_sc_hd__a22o_1 _22333_ (.A1(_11719_),
    .A2(_11725_),
    .B1(_12368_),
    .B2(_12369_),
    .X(_12375_));
 sky130_fd_sc_hd__a22oi_1 _22334_ (.A1(_11979_),
    .A2(_12005_),
    .B1(_12371_),
    .B2(_12372_),
    .Y(_12376_));
 sky130_fd_sc_hd__nand4_2 _22335_ (.A(_11982_),
    .B(_11985_),
    .C(_12373_),
    .D(_12375_),
    .Y(_12377_));
 sky130_fd_sc_hd__a2bb2oi_1 _22336_ (.A1_N(_11981_),
    .A2_N(_11984_),
    .B1(_12373_),
    .B2(_12375_),
    .Y(_12378_));
 sky130_fd_sc_hd__nand4_2 _22337_ (.A(_11979_),
    .B(_12005_),
    .C(_12371_),
    .D(_12372_),
    .Y(_12379_));
 sky130_fd_sc_hd__a31o_1 _22338_ (.A1(_11612_),
    .A2(_11634_),
    .A3(_11635_),
    .B1(_11648_),
    .X(_12380_));
 sky130_fd_sc_hd__o21ai_2 _22339_ (.A1(_11640_),
    .A2(_11648_),
    .B1(_12377_),
    .Y(_12381_));
 sky130_fd_sc_hd__o22ai_1 _22340_ (.A1(_11640_),
    .A2(_11648_),
    .B1(_12376_),
    .B2(_12378_),
    .Y(_12382_));
 sky130_fd_sc_hd__nand3b_1 _22341_ (.A_N(_12380_),
    .B(_12379_),
    .C(_12377_),
    .Y(_12383_));
 sky130_fd_sc_hd__nand2_2 _22342_ (.A(_12382_),
    .B(_12383_),
    .Y(_12384_));
 sky130_fd_sc_hd__o21ai_2 _22343_ (.A1(_11252_),
    .A2(_11993_),
    .B1(_11992_),
    .Y(_12386_));
 sky130_fd_sc_hd__a21boi_2 _22344_ (.A1(_11992_),
    .A2(_11995_),
    .B1_N(_11990_),
    .Y(_12387_));
 sky130_fd_sc_hd__a21o_1 _22345_ (.A1(_11990_),
    .A2(_12386_),
    .B1(_12384_),
    .X(_12388_));
 sky130_fd_sc_hd__nand2_1 _22346_ (.A(_12384_),
    .B(_12387_),
    .Y(_12389_));
 sky130_fd_sc_hd__nand2_1 _22347_ (.A(_12388_),
    .B(_12389_),
    .Y(_12390_));
 sky130_fd_sc_hd__o2111a_1 _22348_ (.A1(_11996_),
    .A2(_12001_),
    .B1(_12000_),
    .C1(_11599_),
    .D1(_11600_),
    .X(_12391_));
 sky130_fd_sc_hd__o2111ai_2 _22349_ (.A1(_11996_),
    .A2(_12001_),
    .B1(_12000_),
    .C1(_11599_),
    .D1(_11600_),
    .Y(_12392_));
 sky130_fd_sc_hd__nor2_2 _22350_ (.A(_11603_),
    .B(_12392_),
    .Y(_12393_));
 sky130_fd_sc_hd__nand2_4 _22351_ (.A(_10810_),
    .B(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__o2111ai_1 _22352_ (.A1(_11591_),
    .A2(_11594_),
    .B1(_11214_),
    .C1(_11595_),
    .D1(_12000_),
    .Y(_12395_));
 sky130_fd_sc_hd__o21ai_1 _22353_ (.A1(_11996_),
    .A2(_12001_),
    .B1(_12395_),
    .Y(_12397_));
 sky130_fd_sc_hd__a21oi_4 _22354_ (.A1(_12391_),
    .A2(_11602_),
    .B1(_12397_),
    .Y(_12398_));
 sky130_fd_sc_hd__nand2_1 _22355_ (.A(_12394_),
    .B(_12398_),
    .Y(_12399_));
 sky130_fd_sc_hd__nand2_2 _22356_ (.A(_10811_),
    .B(_12393_),
    .Y(_12400_));
 sky130_fd_sc_hd__a21oi_4 _22357_ (.A1(_09167_),
    .A2(_09169_),
    .B1(_12400_),
    .Y(_12401_));
 sky130_fd_sc_hd__nor2_1 _22358_ (.A(_12399_),
    .B(_12401_),
    .Y(_12402_));
 sky130_fd_sc_hd__xor2_1 _22359_ (.A(_12390_),
    .B(_12402_),
    .X(net99));
 sky130_fd_sc_hd__a21boi_1 _22360_ (.A1(_12368_),
    .A2(_12370_),
    .B1_N(_12369_),
    .Y(_12403_));
 sky130_fd_sc_hd__o32ai_4 _22361_ (.A1(_11869_),
    .A2(_12006_),
    .A3(_12247_),
    .B1(_12250_),
    .B2(_12360_),
    .Y(_12404_));
 sky130_fd_sc_hd__a31oi_2 _22362_ (.A1(_12116_),
    .A2(_12231_),
    .A3(_12234_),
    .B1(_12114_),
    .Y(_12405_));
 sky130_fd_sc_hd__o311a_1 _22363_ (.A1(_03286_),
    .A2(net44),
    .A3(net319),
    .B1(_09298_),
    .C1(_12076_),
    .X(_12407_));
 sky130_fd_sc_hd__o21ai_2 _22364_ (.A1(net147),
    .A2(_12074_),
    .B1(_12076_),
    .Y(_12408_));
 sky130_fd_sc_hd__a31o_1 _22365_ (.A1(net307),
    .A2(net293),
    .A3(_09654_),
    .B1(_08658_),
    .X(_12409_));
 sky130_fd_sc_hd__o32a_2 _22366_ (.A1(_03960_),
    .A2(_04266_),
    .A3(net57),
    .B1(_09687_),
    .B2(_12409_),
    .X(_12410_));
 sky130_fd_sc_hd__o22ai_4 _22367_ (.A1(_03960_),
    .A2(_08660_),
    .B1(_09687_),
    .B2(_12409_),
    .Y(_12411_));
 sky130_fd_sc_hd__a31oi_4 _22368_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_12411_),
    .Y(_12412_));
 sky130_fd_sc_hd__a31o_1 _22369_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_12411_),
    .X(_12413_));
 sky130_fd_sc_hd__o2111a_2 _22370_ (.A1(net169),
    .A2(net268),
    .B1(_12411_),
    .C1(net319),
    .D1(net33),
    .X(_12414_));
 sky130_fd_sc_hd__o2111ai_4 _22371_ (.A1(net169),
    .A2(net268),
    .B1(_12411_),
    .C1(net319),
    .D1(net33),
    .Y(_12415_));
 sky130_fd_sc_hd__a21oi_1 _22372_ (.A1(_08878_),
    .A2(_12410_),
    .B1(net147),
    .Y(_12416_));
 sky130_fd_sc_hd__a22o_2 _22373_ (.A1(_08882_),
    .A2(_09298_),
    .B1(_12410_),
    .B2(_08878_),
    .X(_12418_));
 sky130_fd_sc_hd__o21ai_4 _22374_ (.A1(_12412_),
    .A2(_12414_),
    .B1(net147),
    .Y(_12419_));
 sky130_fd_sc_hd__o22ai_4 _22375_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_12412_),
    .B2(_12414_),
    .Y(_12420_));
 sky130_fd_sc_hd__nand3_2 _22376_ (.A(_12413_),
    .B(_12415_),
    .C(net147),
    .Y(_12421_));
 sky130_fd_sc_hd__a22oi_4 _22377_ (.A1(_12076_),
    .A2(_12079_),
    .B1(_12420_),
    .B2(_12421_),
    .Y(_12422_));
 sky130_fd_sc_hd__o211ai_4 _22378_ (.A1(net147),
    .A2(_12412_),
    .B1(_12408_),
    .C1(_12419_),
    .Y(_12423_));
 sky130_fd_sc_hd__a2bb2oi_4 _22379_ (.A1_N(_12074_),
    .A2_N(_12407_),
    .B1(_12418_),
    .B2(_12419_),
    .Y(_12424_));
 sky130_fd_sc_hd__nand4_4 _22380_ (.A(_12076_),
    .B(_12079_),
    .C(_12420_),
    .D(_12421_),
    .Y(_12425_));
 sky130_fd_sc_hd__o21ai_2 _22381_ (.A1(_12422_),
    .A2(_12424_),
    .B1(net133),
    .Y(_12426_));
 sky130_fd_sc_hd__o211ai_2 _22382_ (.A1(_10540_),
    .A2(net135),
    .B1(_12423_),
    .C1(_12425_),
    .Y(_12427_));
 sky130_fd_sc_hd__o21ai_2 _22383_ (.A1(_12422_),
    .A2(_12424_),
    .B1(_10546_),
    .Y(_12429_));
 sky130_fd_sc_hd__nand4_4 _22384_ (.A(net138),
    .B(net134),
    .C(_12423_),
    .D(_12425_),
    .Y(_12430_));
 sky130_fd_sc_hd__a32oi_4 _22385_ (.A1(_12077_),
    .A2(_12082_),
    .A3(_12079_),
    .B1(net138),
    .B2(net134),
    .Y(_12431_));
 sky130_fd_sc_hd__a32oi_4 _22386_ (.A1(_12080_),
    .A2(_12081_),
    .A3(_12083_),
    .B1(_12086_),
    .B2(_10546_),
    .Y(_12432_));
 sky130_fd_sc_hd__a21oi_2 _22387_ (.A1(_12429_),
    .A2(_12430_),
    .B1(_12432_),
    .Y(_12433_));
 sky130_fd_sc_hd__o211ai_4 _22388_ (.A1(_12084_),
    .A2(_12431_),
    .B1(_12427_),
    .C1(_12426_),
    .Y(_12434_));
 sky130_fd_sc_hd__nand3_4 _22389_ (.A(_12429_),
    .B(_12430_),
    .C(_12432_),
    .Y(_12435_));
 sky130_fd_sc_hd__a21oi_2 _22390_ (.A1(_12434_),
    .A2(_12435_),
    .B1(_12099_),
    .Y(_12436_));
 sky130_fd_sc_hd__a21o_1 _22391_ (.A1(_12434_),
    .A2(_12435_),
    .B1(_12099_),
    .X(_12437_));
 sky130_fd_sc_hd__o211ai_2 _22392_ (.A1(_11742_),
    .A2(_11042_),
    .B1(_12435_),
    .C1(_12434_),
    .Y(_12438_));
 sky130_fd_sc_hd__a22o_1 _22393_ (.A1(net142),
    .A2(_11743_),
    .B1(_12434_),
    .B2(_12435_),
    .X(_12440_));
 sky130_fd_sc_hd__o2111ai_4 _22394_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net142),
    .C1(_12434_),
    .D1(_12435_),
    .Y(_12441_));
 sky130_fd_sc_hd__nand2_1 _22395_ (.A(_12097_),
    .B(_12098_),
    .Y(_12442_));
 sky130_fd_sc_hd__a31oi_1 _22396_ (.A1(_12090_),
    .A2(_12091_),
    .A3(_12093_),
    .B1(_12098_),
    .Y(_12443_));
 sky130_fd_sc_hd__a22oi_2 _22397_ (.A1(_12095_),
    .A2(_12087_),
    .B1(_12094_),
    .B2(_12099_),
    .Y(_12444_));
 sky130_fd_sc_hd__nand3_4 _22398_ (.A(_12440_),
    .B(_12441_),
    .C(_12444_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand3_2 _22399_ (.A(_12094_),
    .B(_12438_),
    .C(_12442_),
    .Y(_12446_));
 sky130_fd_sc_hd__o211ai_2 _22400_ (.A1(_12096_),
    .A2(_12443_),
    .B1(_12438_),
    .C1(_12437_),
    .Y(_12447_));
 sky130_fd_sc_hd__o21ai_1 _22401_ (.A1(_12436_),
    .A2(_12446_),
    .B1(_12445_),
    .Y(_12448_));
 sky130_fd_sc_hd__a22oi_4 _22402_ (.A1(net25),
    .A2(_10335_),
    .B1(net159),
    .B2(net289),
    .Y(_12449_));
 sky130_fd_sc_hd__a22o_4 _22403_ (.A1(net25),
    .A2(_10335_),
    .B1(net159),
    .B2(net289),
    .X(_12451_));
 sky130_fd_sc_hd__nand2_1 _22404_ (.A(net289),
    .B(_08666_),
    .Y(_12452_));
 sky130_fd_sc_hd__o311a_4 _22405_ (.A1(net25),
    .A2(_08261_),
    .A3(net154),
    .B1(_12022_),
    .C1(_12018_),
    .X(_12453_));
 sky130_fd_sc_hd__o211ai_4 _22406_ (.A1(_08261_),
    .A2(net150),
    .B1(_12022_),
    .C1(_12018_),
    .Y(_12454_));
 sky130_fd_sc_hd__a21oi_1 _22407_ (.A1(_12449_),
    .A2(_12452_),
    .B1(_12454_),
    .Y(_12455_));
 sky130_fd_sc_hd__a21o_1 _22408_ (.A1(_12449_),
    .A2(_12452_),
    .B1(_12454_),
    .X(_12456_));
 sky130_fd_sc_hd__o311a_1 _22409_ (.A1(_04277_),
    .A2(_10324_),
    .A3(net162),
    .B1(_12449_),
    .C1(_12454_),
    .X(_12457_));
 sky130_fd_sc_hd__o221ai_4 _22410_ (.A1(_04277_),
    .A2(_10346_),
    .B1(_10324_),
    .B2(_08669_),
    .C1(_12454_),
    .Y(_12458_));
 sky130_fd_sc_hd__o2bb2ai_2 _22411_ (.A1_N(_12029_),
    .A2_N(_12033_),
    .B1(_12455_),
    .B2(_12457_),
    .Y(_12459_));
 sky130_fd_sc_hd__and4_1 _22412_ (.A(_12029_),
    .B(_12033_),
    .C(_12456_),
    .D(_12458_),
    .X(_12460_));
 sky130_fd_sc_hd__o2111ai_4 _22413_ (.A1(_12025_),
    .A2(_12026_),
    .B1(_12029_),
    .C1(_12456_),
    .D1(_12458_),
    .Y(_12462_));
 sky130_fd_sc_hd__o32a_2 _22414_ (.A1(_01304_),
    .A2(_07498_),
    .A3(_07502_),
    .B1(_01326_),
    .B2(_04223_),
    .X(_12463_));
 sky130_fd_sc_hd__a32o_1 _22415_ (.A1(_07499_),
    .A2(net167),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net21),
    .X(_12464_));
 sky130_fd_sc_hd__and3_1 _22416_ (.A(_07771_),
    .B(_12330_),
    .C(net165),
    .X(_12465_));
 sky130_fd_sc_hd__nor2_1 _22417_ (.A(_04245_),
    .B(_12363_),
    .Y(_12466_));
 sky130_fd_sc_hd__a31oi_4 _22418_ (.A1(_07771_),
    .A2(_12330_),
    .A3(net165),
    .B1(_12466_),
    .Y(_12467_));
 sky130_fd_sc_hd__o211ai_4 _22419_ (.A1(net168),
    .A2(net268),
    .B1(net252),
    .C1(net164),
    .Y(_12468_));
 sky130_fd_sc_hd__or3_2 _22420_ (.A(net35),
    .B(_04256_),
    .C(_03971_),
    .X(_12469_));
 sky130_fd_sc_hd__o21ai_1 _22421_ (.A1(_04256_),
    .A2(_11804_),
    .B1(_12468_),
    .Y(_12470_));
 sky130_fd_sc_hd__a21oi_4 _22422_ (.A1(_12468_),
    .A2(_12469_),
    .B1(_12467_),
    .Y(_12471_));
 sky130_fd_sc_hd__a21o_1 _22423_ (.A1(_12468_),
    .A2(_12469_),
    .B1(_12467_),
    .X(_12473_));
 sky130_fd_sc_hd__o311a_1 _22424_ (.A1(_03971_),
    .A2(net35),
    .A3(_04256_),
    .B1(_12468_),
    .C1(_12467_),
    .X(_12474_));
 sky130_fd_sc_hd__o221ai_2 _22425_ (.A1(_04256_),
    .A2(_11804_),
    .B1(_08209_),
    .B2(_11782_),
    .C1(_12467_),
    .Y(_12475_));
 sky130_fd_sc_hd__o21a_1 _22426_ (.A1(_12471_),
    .A2(_12474_),
    .B1(_12463_),
    .X(_12476_));
 sky130_fd_sc_hd__and3_1 _22427_ (.A(_12464_),
    .B(_12473_),
    .C(_12475_),
    .X(_12477_));
 sky130_fd_sc_hd__o21a_1 _22428_ (.A1(_12471_),
    .A2(_12474_),
    .B1(_12464_),
    .X(_12478_));
 sky130_fd_sc_hd__o21ai_1 _22429_ (.A1(_12471_),
    .A2(_12474_),
    .B1(_12464_),
    .Y(_12479_));
 sky130_fd_sc_hd__and3_1 _22430_ (.A(_12473_),
    .B(_12475_),
    .C(_12463_),
    .X(_12480_));
 sky130_fd_sc_hd__nand3_1 _22431_ (.A(_12473_),
    .B(_12475_),
    .C(_12463_),
    .Y(_12481_));
 sky130_fd_sc_hd__nand4_1 _22432_ (.A(_12459_),
    .B(_12462_),
    .C(_12479_),
    .D(_12481_),
    .Y(_12482_));
 sky130_fd_sc_hd__o2bb2ai_1 _22433_ (.A1_N(_12459_),
    .A2_N(_12462_),
    .B1(_12478_),
    .B2(_12480_),
    .Y(_12484_));
 sky130_fd_sc_hd__o211ai_2 _22434_ (.A1(_12478_),
    .A2(_12480_),
    .B1(_12459_),
    .C1(_12462_),
    .Y(_12485_));
 sky130_fd_sc_hd__o2bb2ai_1 _22435_ (.A1_N(_12459_),
    .A2_N(_12462_),
    .B1(_12476_),
    .B2(_12477_),
    .Y(_12486_));
 sky130_fd_sc_hd__nand3_4 _22436_ (.A(_12486_),
    .B(_11740_),
    .C(_12485_),
    .Y(_12487_));
 sky130_fd_sc_hd__o311a_2 _22437_ (.A1(_10297_),
    .A2(_10538_),
    .A3(_11735_),
    .B1(_12482_),
    .C1(_12484_),
    .X(_12488_));
 sky130_fd_sc_hd__o211ai_2 _22438_ (.A1(net134),
    .A2(_11735_),
    .B1(_12482_),
    .C1(_12484_),
    .Y(_12489_));
 sky130_fd_sc_hd__o31a_1 _22439_ (.A1(_11813_),
    .A2(_12032_),
    .A3(_12035_),
    .B1(_12057_),
    .X(_12490_));
 sky130_fd_sc_hd__a22o_2 _22440_ (.A1(_12038_),
    .A2(_12057_),
    .B1(_12487_),
    .B2(_12489_),
    .X(_12491_));
 sky130_fd_sc_hd__nand4_4 _22441_ (.A(_12038_),
    .B(_12057_),
    .C(_12487_),
    .D(_12489_),
    .Y(_12492_));
 sky130_fd_sc_hd__nand2_1 _22442_ (.A(_12491_),
    .B(_12492_),
    .Y(_12493_));
 sky130_fd_sc_hd__o2111a_1 _22443_ (.A1(_12436_),
    .A2(_12446_),
    .B1(_12491_),
    .C1(_12492_),
    .D1(_12445_),
    .X(_12495_));
 sky130_fd_sc_hd__o2111ai_4 _22444_ (.A1(_12436_),
    .A2(_12446_),
    .B1(_12491_),
    .C1(_12492_),
    .D1(_12445_),
    .Y(_12496_));
 sky130_fd_sc_hd__a22oi_2 _22445_ (.A1(_12445_),
    .A2(_12447_),
    .B1(_12491_),
    .B2(_12492_),
    .Y(_12497_));
 sky130_fd_sc_hd__nand2_1 _22446_ (.A(_12448_),
    .B(_12493_),
    .Y(_12498_));
 sky130_fd_sc_hd__nand4_4 _22447_ (.A(_12105_),
    .B(_12109_),
    .C(_12496_),
    .D(_12498_),
    .Y(_12499_));
 sky130_fd_sc_hd__o2bb2ai_4 _22448_ (.A1_N(_12105_),
    .A2_N(_12109_),
    .B1(_12495_),
    .B2(_12497_),
    .Y(_12500_));
 sky130_fd_sc_hd__o21ai_4 _22449_ (.A1(_12063_),
    .A2(_12060_),
    .B1(_12062_),
    .Y(_12501_));
 sky130_fd_sc_hd__o21ai_4 _22450_ (.A1(_12014_),
    .A2(_12059_),
    .B1(_12065_),
    .Y(_12502_));
 sky130_fd_sc_hd__o211ai_4 _22451_ (.A1(net174),
    .A2(_06759_),
    .B1(_03704_),
    .C1(net193),
    .Y(_12503_));
 sky130_fd_sc_hd__or3_1 _22452_ (.A(net39),
    .B(_04201_),
    .C(_04037_),
    .X(_12504_));
 sky130_fd_sc_hd__a221oi_1 _22453_ (.A1(net203),
    .A2(net272),
    .B1(net171),
    .B2(net20),
    .C1(_02869_),
    .Y(_12506_));
 sky130_fd_sc_hd__and3_1 _22454_ (.A(_04037_),
    .B(net20),
    .C(net37),
    .X(_12507_));
 sky130_fd_sc_hd__a31oi_2 _22455_ (.A1(_07072_),
    .A2(net168),
    .A3(_02858_),
    .B1(_12507_),
    .Y(_12508_));
 sky130_fd_sc_hd__o2bb2ai_2 _22456_ (.A1_N(_12503_),
    .A2_N(_12504_),
    .B1(_12506_),
    .B2(_12507_),
    .Y(_12509_));
 sky130_fd_sc_hd__inv_2 _22457_ (.A(_12509_),
    .Y(_12510_));
 sky130_fd_sc_hd__o211ai_4 _22458_ (.A1(_04201_),
    .A2(_03737_),
    .B1(_12503_),
    .C1(_12508_),
    .Y(_12511_));
 sky130_fd_sc_hd__o311a_1 _22459_ (.A1(net246),
    .A2(_05928_),
    .A3(_06451_),
    .B1(net281),
    .C1(net198),
    .X(_12512_));
 sky130_fd_sc_hd__nor2_1 _22460_ (.A(_04179_),
    .B(_04218_),
    .Y(_12513_));
 sky130_fd_sc_hd__a31o_1 _22461_ (.A1(net198),
    .A2(net172),
    .A3(net281),
    .B1(_12513_),
    .X(_12514_));
 sky130_fd_sc_hd__a21oi_1 _22462_ (.A1(_12509_),
    .A2(_12511_),
    .B1(_12514_),
    .Y(_12515_));
 sky130_fd_sc_hd__a21o_1 _22463_ (.A1(_12509_),
    .A2(_12511_),
    .B1(_12514_),
    .X(_12517_));
 sky130_fd_sc_hd__o211a_4 _22464_ (.A1(_12512_),
    .A2(_12513_),
    .B1(_12509_),
    .C1(_12511_),
    .X(_12518_));
 sky130_fd_sc_hd__o211ai_1 _22465_ (.A1(_12512_),
    .A2(_12513_),
    .B1(_12509_),
    .C1(_12511_),
    .Y(_12519_));
 sky130_fd_sc_hd__o2bb2ai_1 _22466_ (.A1_N(_12044_),
    .A2_N(_12048_),
    .B1(_12040_),
    .B2(_12041_),
    .Y(_12520_));
 sky130_fd_sc_hd__o21ai_2 _22467_ (.A1(_12044_),
    .A2(_12048_),
    .B1(_12520_),
    .Y(_12521_));
 sky130_fd_sc_hd__o21bai_4 _22468_ (.A1(_12515_),
    .A2(_12518_),
    .B1_N(_12521_),
    .Y(_12522_));
 sky130_fd_sc_hd__nand2_2 _22469_ (.A(_12517_),
    .B(_12521_),
    .Y(_12523_));
 sky130_fd_sc_hd__nand3_1 _22470_ (.A(_12517_),
    .B(_12519_),
    .C(_12521_),
    .Y(_12524_));
 sky130_fd_sc_hd__a21o_1 _22471_ (.A1(_12194_),
    .A2(_12195_),
    .B1(_12191_),
    .X(_12525_));
 sky130_fd_sc_hd__a21oi_1 _22472_ (.A1(_12522_),
    .A2(_12524_),
    .B1(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__a21o_2 _22473_ (.A1(_12522_),
    .A2(_12524_),
    .B1(_12525_),
    .X(_12528_));
 sky130_fd_sc_hd__o221a_1 _22474_ (.A1(_12191_),
    .A2(_12197_),
    .B1(_12518_),
    .B2(_12523_),
    .C1(_12522_),
    .X(_12529_));
 sky130_fd_sc_hd__o221ai_4 _22475_ (.A1(_12191_),
    .A2(_12197_),
    .B1(_12518_),
    .B2(_12523_),
    .C1(_12522_),
    .Y(_12530_));
 sky130_fd_sc_hd__o2bb2ai_4 _22476_ (.A1_N(_12185_),
    .A2_N(_12204_),
    .B1(_12205_),
    .B2(_12197_),
    .Y(_12531_));
 sky130_fd_sc_hd__nand3_4 _22477_ (.A(_12528_),
    .B(_12530_),
    .C(_12531_),
    .Y(_12532_));
 sky130_fd_sc_hd__o21bai_4 _22478_ (.A1(_12526_),
    .A2(_12529_),
    .B1_N(_12531_),
    .Y(_12533_));
 sky130_fd_sc_hd__a32o_1 _22479_ (.A1(net178),
    .A2(net177),
    .A3(_04895_),
    .B1(_04897_),
    .B2(net15),
    .X(_12534_));
 sky130_fd_sc_hd__o211ai_2 _22480_ (.A1(net231),
    .A2(_05927_),
    .B1(net279),
    .C1(_05933_),
    .Y(_12535_));
 sky130_fd_sc_hd__or3b_1 _22481_ (.A(net42),
    .B(_04157_),
    .C_N(net41),
    .X(_12536_));
 sky130_fd_sc_hd__a32oi_4 _22482_ (.A1(net202),
    .A2(net173),
    .A3(_04267_),
    .B1(_04269_),
    .B2(net17),
    .Y(_12537_));
 sky130_fd_sc_hd__a21oi_1 _22483_ (.A1(_12535_),
    .A2(_12536_),
    .B1(_12537_),
    .Y(_12539_));
 sky130_fd_sc_hd__a21o_1 _22484_ (.A1(_12535_),
    .A2(_12536_),
    .B1(_12537_),
    .X(_12540_));
 sky130_fd_sc_hd__o211a_1 _22485_ (.A1(_04157_),
    .A2(_04483_),
    .B1(_12535_),
    .C1(_12537_),
    .X(_12541_));
 sky130_fd_sc_hd__o211ai_2 _22486_ (.A1(_04157_),
    .A2(_04483_),
    .B1(_12535_),
    .C1(_12537_),
    .Y(_12542_));
 sky130_fd_sc_hd__o21bai_1 _22487_ (.A1(_12539_),
    .A2(_12541_),
    .B1_N(_12534_),
    .Y(_12543_));
 sky130_fd_sc_hd__nand3_1 _22488_ (.A(_12534_),
    .B(_12540_),
    .C(_12542_),
    .Y(_12544_));
 sky130_fd_sc_hd__o21ai_1 _22489_ (.A1(_12539_),
    .A2(_12541_),
    .B1(_12534_),
    .Y(_12545_));
 sky130_fd_sc_hd__nand3b_1 _22490_ (.A_N(_12534_),
    .B(_12540_),
    .C(_12542_),
    .Y(_12546_));
 sky130_fd_sc_hd__a22oi_2 _22491_ (.A1(_12136_),
    .A2(_12141_),
    .B1(_12543_),
    .B2(_12544_),
    .Y(_12547_));
 sky130_fd_sc_hd__nand3_2 _22492_ (.A(_12143_),
    .B(_12545_),
    .C(_12546_),
    .Y(_12548_));
 sky130_fd_sc_hd__a21oi_1 _22493_ (.A1(_12545_),
    .A2(_12546_),
    .B1(_12143_),
    .Y(_12550_));
 sky130_fd_sc_hd__nand4_2 _22494_ (.A(_12136_),
    .B(_12141_),
    .C(_12543_),
    .D(_12544_),
    .Y(_12551_));
 sky130_fd_sc_hd__a32o_1 _22495_ (.A1(net184),
    .A2(net213),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net11),
    .X(_12552_));
 sky130_fd_sc_hd__nand3_1 _22496_ (.A(net182),
    .B(net179),
    .C(net242),
    .Y(_12553_));
 sky130_fd_sc_hd__or3_1 _22497_ (.A(net45),
    .B(_04135_),
    .C(_04102_),
    .X(_12554_));
 sky130_fd_sc_hd__a32oi_4 _22498_ (.A1(net210),
    .A2(net183),
    .A3(net276),
    .B1(_05228_),
    .B2(net13),
    .Y(_12555_));
 sky130_fd_sc_hd__a21oi_1 _22499_ (.A1(_12553_),
    .A2(_12554_),
    .B1(_12555_),
    .Y(_12556_));
 sky130_fd_sc_hd__a21o_1 _22500_ (.A1(_12553_),
    .A2(_12554_),
    .B1(_12555_),
    .X(_12557_));
 sky130_fd_sc_hd__and3_1 _22501_ (.A(_12555_),
    .B(_12554_),
    .C(_12553_),
    .X(_12558_));
 sky130_fd_sc_hd__o211ai_2 _22502_ (.A1(_04135_),
    .A2(_04989_),
    .B1(_12553_),
    .C1(_12555_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand3b_2 _22503_ (.A_N(_12552_),
    .B(_12557_),
    .C(_12559_),
    .Y(_12561_));
 sky130_fd_sc_hd__o21ai_2 _22504_ (.A1(_12556_),
    .A2(_12558_),
    .B1(_12552_),
    .Y(_12562_));
 sky130_fd_sc_hd__nand2_1 _22505_ (.A(_12561_),
    .B(_12562_),
    .Y(_12563_));
 sky130_fd_sc_hd__and2_1 _22506_ (.A(_12561_),
    .B(_12562_),
    .X(_12564_));
 sky130_fd_sc_hd__and3_1 _22507_ (.A(_12563_),
    .B(_12551_),
    .C(_12548_),
    .X(_12565_));
 sky130_fd_sc_hd__o211a_1 _22508_ (.A1(_12547_),
    .A2(_12550_),
    .B1(_12561_),
    .C1(_12562_),
    .X(_12566_));
 sky130_fd_sc_hd__o21a_1 _22509_ (.A1(_12547_),
    .A2(_12550_),
    .B1(_12563_),
    .X(_12567_));
 sky130_fd_sc_hd__a22o_1 _22510_ (.A1(_12548_),
    .A2(_12551_),
    .B1(_12561_),
    .B2(_12562_),
    .X(_12568_));
 sky130_fd_sc_hd__and3_1 _22511_ (.A(_12548_),
    .B(_12551_),
    .C(_12564_),
    .X(_12569_));
 sky130_fd_sc_hd__nand4_1 _22512_ (.A(_12548_),
    .B(_12551_),
    .C(_12561_),
    .D(_12562_),
    .Y(_12570_));
 sky130_fd_sc_hd__nand2_1 _22513_ (.A(_12568_),
    .B(_12570_),
    .Y(_12572_));
 sky130_fd_sc_hd__o2bb2ai_2 _22514_ (.A1_N(_12532_),
    .A2_N(_12533_),
    .B1(_12567_),
    .B2(_12569_),
    .Y(_12573_));
 sky130_fd_sc_hd__o211ai_2 _22515_ (.A1(_12565_),
    .A2(_12566_),
    .B1(_12532_),
    .C1(_12533_),
    .Y(_12574_));
 sky130_fd_sc_hd__a32oi_4 _22516_ (.A1(_12528_),
    .A2(_12530_),
    .A3(_12531_),
    .B1(_12533_),
    .B2(_12572_),
    .Y(_12575_));
 sky130_fd_sc_hd__a32o_1 _22517_ (.A1(_12528_),
    .A2(_12530_),
    .A3(_12531_),
    .B1(_12533_),
    .B2(_12572_),
    .X(_12576_));
 sky130_fd_sc_hd__o2bb2ai_4 _22518_ (.A1_N(_12532_),
    .A2_N(_12533_),
    .B1(_12565_),
    .B2(_12566_),
    .Y(_12577_));
 sky130_fd_sc_hd__o211ai_4 _22519_ (.A1(_12567_),
    .A2(_12569_),
    .B1(_12532_),
    .C1(_12533_),
    .Y(_12578_));
 sky130_fd_sc_hd__a21oi_1 _22520_ (.A1(_12573_),
    .A2(_12574_),
    .B1(_12502_),
    .Y(_12579_));
 sky130_fd_sc_hd__nand3_4 _22521_ (.A(_12577_),
    .B(_12578_),
    .C(_12501_),
    .Y(_12580_));
 sky130_fd_sc_hd__a21oi_4 _22522_ (.A1(_12577_),
    .A2(_12578_),
    .B1(_12501_),
    .Y(_12581_));
 sky130_fd_sc_hd__nand3_4 _22523_ (.A(_12502_),
    .B(_12573_),
    .C(_12574_),
    .Y(_12583_));
 sky130_fd_sc_hd__a2bb2oi_1 _22524_ (.A1_N(_12213_),
    .A2_N(_12218_),
    .B1(_12580_),
    .B2(_12583_),
    .Y(_12584_));
 sky130_fd_sc_hd__o22ai_2 _22525_ (.A1(_12213_),
    .A2(_12218_),
    .B1(_12579_),
    .B2(_12581_),
    .Y(_12585_));
 sky130_fd_sc_hd__o211a_1 _22526_ (.A1(_12215_),
    .A2(_12217_),
    .B1(_12580_),
    .C1(_12583_),
    .X(_12586_));
 sky130_fd_sc_hd__o2111ai_4 _22527_ (.A1(_12182_),
    .A2(_12215_),
    .B1(_12580_),
    .C1(_12583_),
    .D1(_12214_),
    .Y(_12587_));
 sky130_fd_sc_hd__a21oi_1 _22528_ (.A1(_12580_),
    .A2(_12583_),
    .B1(_12219_),
    .Y(_12588_));
 sky130_fd_sc_hd__o22ai_2 _22529_ (.A1(_12215_),
    .A2(_12217_),
    .B1(_12579_),
    .B2(_12581_),
    .Y(_12589_));
 sky130_fd_sc_hd__and3_1 _22530_ (.A(_12580_),
    .B(_12583_),
    .C(_12219_),
    .X(_12590_));
 sky130_fd_sc_hd__o211ai_2 _22531_ (.A1(_12213_),
    .A2(_12218_),
    .B1(_12580_),
    .C1(_12583_),
    .Y(_12591_));
 sky130_fd_sc_hd__nand4_2 _22532_ (.A(_12499_),
    .B(_12500_),
    .C(_12589_),
    .D(_12591_),
    .Y(_12592_));
 sky130_fd_sc_hd__o2bb2ai_2 _22533_ (.A1_N(_12499_),
    .A2_N(_12500_),
    .B1(_12588_),
    .B2(_12590_),
    .Y(_12594_));
 sky130_fd_sc_hd__nand4_2 _22534_ (.A(_12499_),
    .B(_12500_),
    .C(_12585_),
    .D(_12587_),
    .Y(_12595_));
 sky130_fd_sc_hd__o2bb2ai_2 _22535_ (.A1_N(_12499_),
    .A2_N(_12500_),
    .B1(_12584_),
    .B2(_12586_),
    .Y(_12596_));
 sky130_fd_sc_hd__nand4_2 _22536_ (.A(_12115_),
    .B(_12242_),
    .C(_12595_),
    .D(_12596_),
    .Y(_12597_));
 sky130_fd_sc_hd__o2111a_1 _22537_ (.A1(_12114_),
    .A2(_12240_),
    .B1(_12592_),
    .C1(_12594_),
    .D1(_12116_),
    .X(_12598_));
 sky130_fd_sc_hd__o2111ai_4 _22538_ (.A1(_12114_),
    .A2(_12240_),
    .B1(_12592_),
    .C1(_12594_),
    .D1(_12116_),
    .Y(_12599_));
 sky130_fd_sc_hd__a21o_1 _22539_ (.A1(_12331_),
    .A2(_12295_),
    .B1(_12327_),
    .X(_12600_));
 sky130_fd_sc_hd__a21oi_1 _22540_ (.A1(_12331_),
    .A2(_12295_),
    .B1(_12327_),
    .Y(_12601_));
 sky130_fd_sc_hd__a21oi_1 _22541_ (.A1(_12299_),
    .A2(_12307_),
    .B1(_12304_),
    .Y(_12602_));
 sky130_fd_sc_hd__a32oi_4 _22542_ (.A1(net229),
    .A2(net227),
    .A3(net273),
    .B1(_06326_),
    .B2(net8),
    .Y(_12603_));
 sky130_fd_sc_hd__or3b_1 _22543_ (.A(_04080_),
    .B(net48),
    .C_N(net47),
    .X(_12605_));
 sky130_fd_sc_hd__o211ai_2 _22544_ (.A1(net233),
    .A2(_04557_),
    .B1(_05762_),
    .C1(net217),
    .Y(_12606_));
 sky130_fd_sc_hd__a32oi_4 _22545_ (.A1(net217),
    .A2(net186),
    .A3(_05762_),
    .B1(_05765_),
    .B2(net10),
    .Y(_12607_));
 sky130_fd_sc_hd__nand3_1 _22546_ (.A(_04409_),
    .B(net221),
    .C(net274),
    .Y(_12608_));
 sky130_fd_sc_hd__or3b_1 _22547_ (.A(_04069_),
    .B(net49),
    .C_N(net48),
    .X(_12609_));
 sky130_fd_sc_hd__a32oi_4 _22548_ (.A1(_04409_),
    .A2(net221),
    .A3(net274),
    .B1(_06029_),
    .B2(net9),
    .Y(_12610_));
 sky130_fd_sc_hd__a21oi_1 _22549_ (.A1(_12608_),
    .A2(_12609_),
    .B1(_12607_),
    .Y(_12611_));
 sky130_fd_sc_hd__a22o_1 _22550_ (.A1(_12605_),
    .A2(_12606_),
    .B1(_12608_),
    .B2(_12609_),
    .X(_12612_));
 sky130_fd_sc_hd__nand3_1 _22551_ (.A(_12603_),
    .B(_12607_),
    .C(_12610_),
    .Y(_12613_));
 sky130_fd_sc_hd__a21oi_1 _22552_ (.A1(_12607_),
    .A2(_12610_),
    .B1(_12603_),
    .Y(_12614_));
 sky130_fd_sc_hd__a41o_2 _22553_ (.A1(_12605_),
    .A2(_12606_),
    .A3(_12608_),
    .A4(_12609_),
    .B1(_12603_),
    .X(_12616_));
 sky130_fd_sc_hd__o21ai_1 _22554_ (.A1(_12607_),
    .A2(_12610_),
    .B1(_12616_),
    .Y(_12617_));
 sky130_fd_sc_hd__o211ai_4 _22555_ (.A1(_12607_),
    .A2(_12610_),
    .B1(_12613_),
    .C1(_12616_),
    .Y(_12618_));
 sky130_fd_sc_hd__a221o_2 _22556_ (.A1(_12605_),
    .A2(_12606_),
    .B1(_12608_),
    .B2(_12609_),
    .C1(_12603_),
    .X(_12619_));
 sky130_fd_sc_hd__o211a_1 _22557_ (.A1(_12612_),
    .A2(_12603_),
    .B1(_12167_),
    .C1(_12618_),
    .X(_12620_));
 sky130_fd_sc_hd__o211ai_2 _22558_ (.A1(_12612_),
    .A2(_12603_),
    .B1(_12167_),
    .C1(_12618_),
    .Y(_12621_));
 sky130_fd_sc_hd__a21oi_4 _22559_ (.A1(_12618_),
    .A2(_12619_),
    .B1(_12167_),
    .Y(_12622_));
 sky130_fd_sc_hd__a22o_1 _22560_ (.A1(_12163_),
    .A2(_12165_),
    .B1(_12618_),
    .B2(_12619_),
    .X(_12623_));
 sky130_fd_sc_hd__o21a_2 _22561_ (.A1(_12620_),
    .A2(_12622_),
    .B1(_12602_),
    .X(_12624_));
 sky130_fd_sc_hd__a31o_1 _22562_ (.A1(_12167_),
    .A2(_12618_),
    .A3(_12619_),
    .B1(_12602_),
    .X(_12625_));
 sky130_fd_sc_hd__o211a_1 _22563_ (.A1(_12304_),
    .A2(_12310_),
    .B1(_12621_),
    .C1(_12623_),
    .X(_12627_));
 sky130_fd_sc_hd__o22ai_2 _22564_ (.A1(_12304_),
    .A2(_12310_),
    .B1(_12620_),
    .B2(_12622_),
    .Y(_12628_));
 sky130_fd_sc_hd__nand3_1 _22565_ (.A(_12623_),
    .B(_12602_),
    .C(_12621_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand3_2 _22566_ (.A(_12176_),
    .B(_12628_),
    .C(_12629_),
    .Y(_12630_));
 sky130_fd_sc_hd__inv_2 _22567_ (.A(_12630_),
    .Y(_12631_));
 sky130_fd_sc_hd__o211ai_4 _22568_ (.A1(_12622_),
    .A2(_12625_),
    .B1(_12150_),
    .C1(_12174_),
    .Y(_12632_));
 sky130_fd_sc_hd__a21oi_1 _22569_ (.A1(_12628_),
    .A2(_12629_),
    .B1(_12176_),
    .Y(_12633_));
 sky130_fd_sc_hd__o21ai_1 _22570_ (.A1(_12624_),
    .A2(_12632_),
    .B1(_12630_),
    .Y(_12634_));
 sky130_fd_sc_hd__o31a_1 _22571_ (.A1(_11671_),
    .A2(_11676_),
    .A3(_12316_),
    .B1(_12320_),
    .X(_12635_));
 sky130_fd_sc_hd__o21ai_1 _22572_ (.A1(_12318_),
    .A2(_12324_),
    .B1(_12634_),
    .Y(_12636_));
 sky130_fd_sc_hd__o2111ai_4 _22573_ (.A1(_12624_),
    .A2(_12632_),
    .B1(_12630_),
    .C1(_12320_),
    .D1(_12325_),
    .Y(_12638_));
 sky130_fd_sc_hd__nand2_1 _22574_ (.A(_12634_),
    .B(_12635_),
    .Y(_12639_));
 sky130_fd_sc_hd__a31o_1 _22575_ (.A1(_12176_),
    .A2(_12628_),
    .A3(_12629_),
    .B1(_12635_),
    .X(_12640_));
 sky130_fd_sc_hd__o221a_2 _22576_ (.A1(_12318_),
    .A2(_12324_),
    .B1(_12624_),
    .B2(_12632_),
    .C1(_12630_),
    .X(_12641_));
 sky130_fd_sc_hd__nand3_4 _22577_ (.A(_12601_),
    .B(_12636_),
    .C(_12638_),
    .Y(_12642_));
 sky130_fd_sc_hd__inv_2 _22578_ (.A(_12642_),
    .Y(_12643_));
 sky130_fd_sc_hd__o2bb2ai_2 _22579_ (.A1_N(_12635_),
    .A2_N(_12634_),
    .B1(_12334_),
    .B2(_12327_),
    .Y(_12644_));
 sky130_fd_sc_hd__o211ai_4 _22580_ (.A1(_12633_),
    .A2(_12640_),
    .B1(_12639_),
    .C1(_12600_),
    .Y(_12645_));
 sky130_fd_sc_hd__a32o_1 _22581_ (.A1(_11354_),
    .A2(net253),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net3),
    .X(_12646_));
 sky130_fd_sc_hd__and3b_1 _22582_ (.A_N(net54),
    .B(net53),
    .C(net4),
    .X(_12647_));
 sky130_fd_sc_hd__o311a_2 _22583_ (.A1(net3),
    .A2(_09665_),
    .A3(_12988_),
    .B1(_07642_),
    .C1(net234),
    .X(_12649_));
 sky130_fd_sc_hd__a31o_1 _22584_ (.A1(net234),
    .A2(net251),
    .A3(_07642_),
    .B1(_12647_),
    .X(_12650_));
 sky130_fd_sc_hd__a32oi_4 _22585_ (.A1(_00625_),
    .A2(net250),
    .A3(net239),
    .B1(_07308_),
    .B2(net5),
    .Y(_12651_));
 sky130_fd_sc_hd__a32o_1 _22586_ (.A1(_00625_),
    .A2(net250),
    .A3(net239),
    .B1(_07308_),
    .B2(net5),
    .X(_12652_));
 sky130_fd_sc_hd__nand2_1 _22587_ (.A(net248),
    .B(net269),
    .Y(_12653_));
 sky130_fd_sc_hd__o211ai_1 _22588_ (.A1(net253),
    .A2(_02442_),
    .B1(net269),
    .C1(_02421_),
    .Y(_12654_));
 sky130_fd_sc_hd__or3b_1 _22589_ (.A(_04026_),
    .B(net52),
    .C_N(net51),
    .X(_12655_));
 sky130_fd_sc_hd__o21ai_1 _22590_ (.A1(_02410_),
    .A2(_12653_),
    .B1(_12655_),
    .Y(_12656_));
 sky130_fd_sc_hd__o2111ai_2 _22591_ (.A1(net253),
    .A2(_03954_),
    .B1(net51),
    .C1(_03952_),
    .D1(_04190_),
    .Y(_12657_));
 sky130_fd_sc_hd__or3_1 _22592_ (.A(net51),
    .B(_04190_),
    .C(_04048_),
    .X(_12658_));
 sky130_fd_sc_hd__o31ai_1 _22593_ (.A1(_06864_),
    .A2(_03957_),
    .A3(_03951_),
    .B1(_12658_),
    .Y(_12660_));
 sky130_fd_sc_hd__a22oi_1 _22594_ (.A1(_12654_),
    .A2(_12655_),
    .B1(_12657_),
    .B2(_12658_),
    .Y(_12661_));
 sky130_fd_sc_hd__a22o_2 _22595_ (.A1(_12654_),
    .A2(_12655_),
    .B1(_12657_),
    .B2(_12658_),
    .X(_12662_));
 sky130_fd_sc_hd__nor2_2 _22596_ (.A(_12656_),
    .B(_12660_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand3b_1 _22597_ (.A_N(_12656_),
    .B(_12657_),
    .C(_12658_),
    .Y(_12664_));
 sky130_fd_sc_hd__o21ai_1 _22598_ (.A1(_12661_),
    .A2(_12663_),
    .B1(_12652_),
    .Y(_12665_));
 sky130_fd_sc_hd__nand3_1 _22599_ (.A(_12662_),
    .B(_12664_),
    .C(_12651_),
    .Y(_12666_));
 sky130_fd_sc_hd__o21ai_1 _22600_ (.A1(_12661_),
    .A2(_12663_),
    .B1(_12651_),
    .Y(_12667_));
 sky130_fd_sc_hd__nand3_1 _22601_ (.A(_12652_),
    .B(_12662_),
    .C(_12664_),
    .Y(_12668_));
 sky130_fd_sc_hd__o21ai_1 _22602_ (.A1(_12259_),
    .A2(_12268_),
    .B1(_12267_),
    .Y(_12669_));
 sky130_fd_sc_hd__a21oi_1 _22603_ (.A1(_12260_),
    .A2(_12269_),
    .B1(_12266_),
    .Y(_12671_));
 sky130_fd_sc_hd__nand3_1 _22604_ (.A(_12665_),
    .B(_12666_),
    .C(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__nand3_2 _22605_ (.A(_12667_),
    .B(_12668_),
    .C(_12669_),
    .Y(_12673_));
 sky130_fd_sc_hd__a21o_1 _22606_ (.A1(_12672_),
    .A2(_12673_),
    .B1(_12650_),
    .X(_12674_));
 sky130_fd_sc_hd__o211ai_2 _22607_ (.A1(_12647_),
    .A2(_12649_),
    .B1(_12672_),
    .C1(_12673_),
    .Y(_12675_));
 sky130_fd_sc_hd__a31oi_1 _22608_ (.A1(_12271_),
    .A2(_12257_),
    .A3(_12270_),
    .B1(_12256_),
    .Y(_12676_));
 sky130_fd_sc_hd__a31o_1 _22609_ (.A1(_12271_),
    .A2(_12257_),
    .A3(_12270_),
    .B1(_12256_),
    .X(_12677_));
 sky130_fd_sc_hd__o2bb2ai_1 _22610_ (.A1_N(_12674_),
    .A2_N(_12675_),
    .B1(_12676_),
    .B2(_12274_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand4_4 _22611_ (.A(_12276_),
    .B(_12674_),
    .C(_12675_),
    .D(_12677_),
    .Y(_12679_));
 sky130_fd_sc_hd__a21oi_2 _22612_ (.A1(_12678_),
    .A2(_12679_),
    .B1(_12646_),
    .Y(_12680_));
 sky130_fd_sc_hd__and3_1 _22613_ (.A(_12646_),
    .B(_12678_),
    .C(_12679_),
    .X(_12682_));
 sky130_fd_sc_hd__inv_2 _22614_ (.A(_12682_),
    .Y(_12683_));
 sky130_fd_sc_hd__nor2_1 _22615_ (.A(_12680_),
    .B(_12682_),
    .Y(_12684_));
 sky130_fd_sc_hd__o211a_1 _22616_ (.A1(_12641_),
    .A2(_12644_),
    .B1(_12684_),
    .C1(_12642_),
    .X(_12685_));
 sky130_fd_sc_hd__o211ai_4 _22617_ (.A1(_12641_),
    .A2(_12644_),
    .B1(_12684_),
    .C1(_12642_),
    .Y(_12686_));
 sky130_fd_sc_hd__a21oi_1 _22618_ (.A1(_12642_),
    .A2(_12645_),
    .B1(_12684_),
    .Y(_12687_));
 sky130_fd_sc_hd__o2bb2ai_2 _22619_ (.A1_N(_12642_),
    .A2_N(_12645_),
    .B1(_12680_),
    .B2(_12682_),
    .Y(_12688_));
 sky130_fd_sc_hd__o2bb2ai_2 _22620_ (.A1_N(_12229_),
    .A2_N(_12237_),
    .B1(_12685_),
    .B2(_12687_),
    .Y(_12689_));
 sky130_fd_sc_hd__and3_1 _22621_ (.A(_12238_),
    .B(_12686_),
    .C(_12688_),
    .X(_12690_));
 sky130_fd_sc_hd__nand4_4 _22622_ (.A(_12229_),
    .B(_12237_),
    .C(_12686_),
    .D(_12688_),
    .Y(_12691_));
 sky130_fd_sc_hd__and3_1 _22623_ (.A(_12289_),
    .B(_12291_),
    .C(_12342_),
    .X(_12693_));
 sky130_fd_sc_hd__a31o_1 _22624_ (.A1(_12289_),
    .A2(_12291_),
    .A3(_12342_),
    .B1(_12344_),
    .X(_12694_));
 sky130_fd_sc_hd__and3_1 _22625_ (.A(_12689_),
    .B(_12691_),
    .C(_12694_),
    .X(_12695_));
 sky130_fd_sc_hd__a21oi_1 _22626_ (.A1(_12689_),
    .A2(_12691_),
    .B1(_12694_),
    .Y(_12696_));
 sky130_fd_sc_hd__o2bb2ai_2 _22627_ (.A1_N(_12689_),
    .A2_N(_12691_),
    .B1(_12693_),
    .B2(_12344_),
    .Y(_12697_));
 sky130_fd_sc_hd__o2111ai_4 _22628_ (.A1(_12293_),
    .A2(_12340_),
    .B1(_12345_),
    .C1(_12689_),
    .D1(_12691_),
    .Y(_12698_));
 sky130_fd_sc_hd__nand2_1 _22629_ (.A(_12697_),
    .B(_12698_),
    .Y(_12699_));
 sky130_fd_sc_hd__o2bb2ai_2 _22630_ (.A1_N(_12597_),
    .A2_N(_12599_),
    .B1(_12695_),
    .B2(_12696_),
    .Y(_12700_));
 sky130_fd_sc_hd__a32oi_4 _22631_ (.A1(_12405_),
    .A2(_12595_),
    .A3(_12596_),
    .B1(_12697_),
    .B2(_12698_),
    .Y(_12701_));
 sky130_fd_sc_hd__nand3_2 _22632_ (.A(_12699_),
    .B(_12599_),
    .C(_12597_),
    .Y(_12702_));
 sky130_fd_sc_hd__a21oi_2 _22633_ (.A1(_12700_),
    .A2(_12702_),
    .B1(_12404_),
    .Y(_12704_));
 sky130_fd_sc_hd__a21o_1 _22634_ (.A1(_12700_),
    .A2(_12702_),
    .B1(_12404_),
    .X(_12705_));
 sky130_fd_sc_hd__o211a_1 _22635_ (.A1(_12248_),
    .A2(_12361_),
    .B1(_12700_),
    .C1(_12702_),
    .X(_12706_));
 sky130_fd_sc_hd__o211ai_2 _22636_ (.A1(_12248_),
    .A2(_12361_),
    .B1(_12700_),
    .C1(_12702_),
    .Y(_12707_));
 sky130_fd_sc_hd__a21boi_2 _22637_ (.A1(_12351_),
    .A2(_12353_),
    .B1_N(_12350_),
    .Y(_12708_));
 sky130_fd_sc_hd__o21bai_1 _22638_ (.A1(_12704_),
    .A2(_12706_),
    .B1_N(_12708_),
    .Y(_12709_));
 sky130_fd_sc_hd__nand3_1 _22639_ (.A(_12705_),
    .B(_12707_),
    .C(_12708_),
    .Y(_12710_));
 sky130_fd_sc_hd__o21ai_1 _22640_ (.A1(_12704_),
    .A2(_12706_),
    .B1(_12708_),
    .Y(_12711_));
 sky130_fd_sc_hd__nand3b_1 _22641_ (.A_N(_12708_),
    .B(_12707_),
    .C(_12705_),
    .Y(_12712_));
 sky130_fd_sc_hd__nand3_1 _22642_ (.A(_12403_),
    .B(_12709_),
    .C(_12710_),
    .Y(_12713_));
 sky130_fd_sc_hd__nand3b_1 _22643_ (.A_N(_12403_),
    .B(_12711_),
    .C(_12712_),
    .Y(_12715_));
 sky130_fd_sc_hd__nor2_1 _22644_ (.A(_12254_),
    .B(_12285_),
    .Y(_12716_));
 sky130_fd_sc_hd__o21a_1 _22645_ (.A1(_12254_),
    .A2(_12285_),
    .B1(_12283_),
    .X(_12717_));
 sky130_fd_sc_hd__o2bb2ai_1 _22646_ (.A1_N(_12713_),
    .A2_N(_12715_),
    .B1(_12716_),
    .B2(_12284_),
    .Y(_12718_));
 sky130_fd_sc_hd__nand3_1 _22647_ (.A(_12713_),
    .B(_12715_),
    .C(_12717_),
    .Y(_12719_));
 sky130_fd_sc_hd__a21oi_1 _22648_ (.A1(_12377_),
    .A2(_12380_),
    .B1(_12378_),
    .Y(_12720_));
 sky130_fd_sc_hd__nand3_1 _22649_ (.A(_12718_),
    .B(_12719_),
    .C(_12720_),
    .Y(_12721_));
 sky130_fd_sc_hd__a22oi_2 _22650_ (.A1(_12379_),
    .A2(_12381_),
    .B1(_12718_),
    .B2(_12719_),
    .Y(_12722_));
 sky130_fd_sc_hd__a22o_1 _22651_ (.A1(_12379_),
    .A2(_12381_),
    .B1(_12718_),
    .B2(_12719_),
    .X(_12723_));
 sky130_fd_sc_hd__nand2_1 _22652_ (.A(_12721_),
    .B(_12723_),
    .Y(_12724_));
 sky130_fd_sc_hd__o22a_1 _22653_ (.A1(_12384_),
    .A2(_12387_),
    .B1(_12399_),
    .B2(_12401_),
    .X(_12726_));
 sky130_fd_sc_hd__a31o_1 _22654_ (.A1(_11990_),
    .A2(_12384_),
    .A3(_12386_),
    .B1(_12726_),
    .X(_12727_));
 sky130_fd_sc_hd__xnor2_1 _22655_ (.A(_12724_),
    .B(_12727_),
    .Y(net100));
 sky130_fd_sc_hd__a21boi_2 _22656_ (.A1(_12715_),
    .A2(_12717_),
    .B1_N(_12713_),
    .Y(_12728_));
 sky130_fd_sc_hd__nand2_1 _22657_ (.A(_12679_),
    .B(_12683_),
    .Y(_12729_));
 sky130_fd_sc_hd__a31o_1 _22658_ (.A1(_12238_),
    .A2(_12686_),
    .A3(_12688_),
    .B1(_12695_),
    .X(_12730_));
 sky130_fd_sc_hd__a21oi_1 _22659_ (.A1(_12699_),
    .A2(_12597_),
    .B1(_12598_),
    .Y(_12731_));
 sky130_fd_sc_hd__a31oi_2 _22660_ (.A1(_12501_),
    .A2(_12577_),
    .A3(_12578_),
    .B1(_12219_),
    .Y(_12732_));
 sky130_fd_sc_hd__a31o_1 _22661_ (.A1(_12501_),
    .A2(_12577_),
    .A3(_12578_),
    .B1(_12219_),
    .X(_12733_));
 sky130_fd_sc_hd__nand3_1 _22662_ (.A(net217),
    .B(net186),
    .C(net274),
    .Y(_12734_));
 sky130_fd_sc_hd__or3b_1 _22663_ (.A(_04080_),
    .B(net49),
    .C_N(net48),
    .X(_12736_));
 sky130_fd_sc_hd__o211ai_2 _22664_ (.A1(net233),
    .A2(_04787_),
    .B1(_05762_),
    .C1(net213),
    .Y(_12737_));
 sky130_fd_sc_hd__or3b_1 _22665_ (.A(_04091_),
    .B(net48),
    .C_N(net47),
    .X(_12738_));
 sky130_fd_sc_hd__a22o_1 _22666_ (.A1(_12734_),
    .A2(_12736_),
    .B1(_12737_),
    .B2(_12738_),
    .X(_12739_));
 sky130_fd_sc_hd__inv_2 _22667_ (.A(_12739_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand4_2 _22668_ (.A(_12734_),
    .B(_12736_),
    .C(_12737_),
    .D(_12738_),
    .Y(_12741_));
 sky130_fd_sc_hd__o311a_1 _22669_ (.A1(net7),
    .A2(net248),
    .A3(_04407_),
    .B1(net273),
    .C1(net221),
    .X(_12742_));
 sky130_fd_sc_hd__and3_1 _22670_ (.A(_04190_),
    .B(net49),
    .C(net9),
    .X(_12743_));
 sky130_fd_sc_hd__a31o_1 _22671_ (.A1(_04409_),
    .A2(net221),
    .A3(net273),
    .B1(_12743_),
    .X(_12744_));
 sky130_fd_sc_hd__a21oi_1 _22672_ (.A1(_12739_),
    .A2(_12741_),
    .B1(_12744_),
    .Y(_12745_));
 sky130_fd_sc_hd__a21o_1 _22673_ (.A1(_12739_),
    .A2(_12741_),
    .B1(_12744_),
    .X(_12747_));
 sky130_fd_sc_hd__o211a_2 _22674_ (.A1(_12742_),
    .A2(_12743_),
    .B1(_12739_),
    .C1(_12741_),
    .X(_12748_));
 sky130_fd_sc_hd__o211ai_2 _22675_ (.A1(_12742_),
    .A2(_12743_),
    .B1(_12739_),
    .C1(_12741_),
    .Y(_12749_));
 sky130_fd_sc_hd__a21o_1 _22676_ (.A1(_12552_),
    .A2(_12559_),
    .B1(_12556_),
    .X(_12750_));
 sky130_fd_sc_hd__a21oi_1 _22677_ (.A1(_12552_),
    .A2(_12559_),
    .B1(_12556_),
    .Y(_12751_));
 sky130_fd_sc_hd__a21oi_1 _22678_ (.A1(_12747_),
    .A2(_12749_),
    .B1(_12750_),
    .Y(_12752_));
 sky130_fd_sc_hd__o21ai_2 _22679_ (.A1(_12745_),
    .A2(_12748_),
    .B1(_12751_),
    .Y(_12753_));
 sky130_fd_sc_hd__nor3_2 _22680_ (.A(_12745_),
    .B(_12751_),
    .C(_12748_),
    .Y(_12754_));
 sky130_fd_sc_hd__nand3_2 _22681_ (.A(_12750_),
    .B(_12749_),
    .C(_12747_),
    .Y(_12755_));
 sky130_fd_sc_hd__a21o_1 _22682_ (.A1(_12753_),
    .A2(_12755_),
    .B1(_12617_),
    .X(_12756_));
 sky130_fd_sc_hd__o21ai_1 _22683_ (.A1(_12611_),
    .A2(_12614_),
    .B1(_12753_),
    .Y(_12758_));
 sky130_fd_sc_hd__o22ai_2 _22684_ (.A1(_12611_),
    .A2(_12614_),
    .B1(_12752_),
    .B2(_12754_),
    .Y(_12759_));
 sky130_fd_sc_hd__o2111ai_4 _22685_ (.A1(_12607_),
    .A2(_12610_),
    .B1(_12616_),
    .C1(_12753_),
    .D1(_12755_),
    .Y(_12760_));
 sky130_fd_sc_hd__a31oi_2 _22686_ (.A1(_12551_),
    .A2(_12561_),
    .A3(_12562_),
    .B1(_12547_),
    .Y(_12761_));
 sky130_fd_sc_hd__a21oi_2 _22687_ (.A1(_12563_),
    .A2(_12548_),
    .B1(_12550_),
    .Y(_12762_));
 sky130_fd_sc_hd__nand3_2 _22688_ (.A(_12759_),
    .B(_12760_),
    .C(_12762_),
    .Y(_12763_));
 sky130_fd_sc_hd__a21oi_2 _22689_ (.A1(_12759_),
    .A2(_12760_),
    .B1(_12762_),
    .Y(_12764_));
 sky130_fd_sc_hd__o211ai_4 _22690_ (.A1(_12754_),
    .A2(_12758_),
    .B1(_12761_),
    .C1(_12756_),
    .Y(_12765_));
 sky130_fd_sc_hd__and3_1 _22691_ (.A(_12305_),
    .B(_12311_),
    .C(_12623_),
    .X(_12766_));
 sky130_fd_sc_hd__o31a_1 _22692_ (.A1(_12304_),
    .A2(_12310_),
    .A3(_12622_),
    .B1(_12621_),
    .X(_12767_));
 sky130_fd_sc_hd__o2bb2ai_2 _22693_ (.A1_N(_12763_),
    .A2_N(_12765_),
    .B1(_12766_),
    .B2(_12620_),
    .Y(_12769_));
 sky130_fd_sc_hd__o21a_1 _22694_ (.A1(_12622_),
    .A2(_12627_),
    .B1(_12763_),
    .X(_12770_));
 sky130_fd_sc_hd__o211ai_4 _22695_ (.A1(_12622_),
    .A2(_12627_),
    .B1(_12763_),
    .C1(_12765_),
    .Y(_12771_));
 sky130_fd_sc_hd__o211a_1 _22696_ (.A1(_12624_),
    .A2(_12632_),
    .B1(_12320_),
    .C1(_12325_),
    .X(_12772_));
 sky130_fd_sc_hd__o21ai_1 _22697_ (.A1(_12624_),
    .A2(_12632_),
    .B1(_12640_),
    .Y(_12773_));
 sky130_fd_sc_hd__and3_1 _22698_ (.A(_12773_),
    .B(_12771_),
    .C(_12769_),
    .X(_12774_));
 sky130_fd_sc_hd__nand3_2 _22699_ (.A(_12773_),
    .B(_12771_),
    .C(_12769_),
    .Y(_12775_));
 sky130_fd_sc_hd__o2bb2a_1 _22700_ (.A1_N(_12769_),
    .A2_N(_12771_),
    .B1(_12772_),
    .B2(_12631_),
    .X(_12776_));
 sky130_fd_sc_hd__o2bb2ai_4 _22701_ (.A1_N(_12769_),
    .A2_N(_12771_),
    .B1(_12772_),
    .B2(_12631_),
    .Y(_12777_));
 sky130_fd_sc_hd__o21ai_2 _22702_ (.A1(_12647_),
    .A2(_12649_),
    .B1(_12672_),
    .Y(_12778_));
 sky130_fd_sc_hd__a32oi_2 _22703_ (.A1(_00625_),
    .A2(net250),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net5),
    .Y(_12780_));
 sky130_fd_sc_hd__a32o_1 _22704_ (.A1(_00625_),
    .A2(net250),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net5),
    .X(_12781_));
 sky130_fd_sc_hd__o21ai_1 _22705_ (.A1(_12651_),
    .A2(_12663_),
    .B1(_12662_),
    .Y(_12782_));
 sky130_fd_sc_hd__a22oi_2 _22706_ (.A1(_02464_),
    .A2(net239),
    .B1(_07308_),
    .B2(net6),
    .Y(_12783_));
 sky130_fd_sc_hd__a32o_1 _22707_ (.A1(_02421_),
    .A2(net248),
    .A3(net239),
    .B1(_07308_),
    .B2(net6),
    .X(_12784_));
 sky130_fd_sc_hd__a32oi_4 _22708_ (.A1(net229),
    .A2(net227),
    .A3(net240),
    .B1(_06865_),
    .B2(net8),
    .Y(_12785_));
 sky130_fd_sc_hd__a32o_1 _22709_ (.A1(net229),
    .A2(net227),
    .A3(net240),
    .B1(_06865_),
    .B2(net8),
    .X(_12786_));
 sky130_fd_sc_hd__nor2_1 _22710_ (.A(_04048_),
    .B(_07226_),
    .Y(_12787_));
 sky130_fd_sc_hd__a31oi_2 _22711_ (.A1(_03952_),
    .A2(net233),
    .A3(net269),
    .B1(_12787_),
    .Y(_12788_));
 sky130_fd_sc_hd__a31o_1 _22712_ (.A1(_03952_),
    .A2(net233),
    .A3(net269),
    .B1(_12787_),
    .X(_12789_));
 sky130_fd_sc_hd__nand2_1 _22713_ (.A(_12786_),
    .B(_12789_),
    .Y(_12791_));
 sky130_fd_sc_hd__o221a_1 _22714_ (.A1(_03961_),
    .A2(_07224_),
    .B1(_07226_),
    .B2(_04048_),
    .C1(_12785_),
    .X(_12792_));
 sky130_fd_sc_hd__nand2_2 _22715_ (.A(_12785_),
    .B(_12788_),
    .Y(_12793_));
 sky130_fd_sc_hd__a21o_1 _22716_ (.A1(_12791_),
    .A2(_12793_),
    .B1(_12784_),
    .X(_12794_));
 sky130_fd_sc_hd__o21ai_1 _22717_ (.A1(_12785_),
    .A2(_12788_),
    .B1(_12784_),
    .Y(_12795_));
 sky130_fd_sc_hd__nand3_1 _22718_ (.A(_12791_),
    .B(_12793_),
    .C(_12783_),
    .Y(_12796_));
 sky130_fd_sc_hd__a21o_1 _22719_ (.A1(_12791_),
    .A2(_12793_),
    .B1(_12783_),
    .X(_12797_));
 sky130_fd_sc_hd__o2111ai_4 _22720_ (.A1(_12651_),
    .A2(_12663_),
    .B1(_12796_),
    .C1(_12797_),
    .D1(_12662_),
    .Y(_12798_));
 sky130_fd_sc_hd__o211ai_2 _22721_ (.A1(_12792_),
    .A2(_12795_),
    .B1(_12782_),
    .C1(_12794_),
    .Y(_12799_));
 sky130_fd_sc_hd__a21o_1 _22722_ (.A1(_12798_),
    .A2(_12799_),
    .B1(_12780_),
    .X(_12800_));
 sky130_fd_sc_hd__nand3_2 _22723_ (.A(_12798_),
    .B(_12799_),
    .C(_12780_),
    .Y(_12802_));
 sky130_fd_sc_hd__nand4_4 _22724_ (.A(_12673_),
    .B(_12778_),
    .C(_12800_),
    .D(_12802_),
    .Y(_12803_));
 sky130_fd_sc_hd__inv_2 _22725_ (.A(_12803_),
    .Y(_12804_));
 sky130_fd_sc_hd__a22o_1 _22726_ (.A1(_12673_),
    .A2(_12778_),
    .B1(_12800_),
    .B2(_12802_),
    .X(_12805_));
 sky130_fd_sc_hd__inv_2 _22727_ (.A(_12805_),
    .Y(_12806_));
 sky130_fd_sc_hd__a32o_1 _22728_ (.A1(net234),
    .A2(net251),
    .A3(_08005_),
    .B1(_08006_),
    .B2(net4),
    .X(_12807_));
 sky130_fd_sc_hd__a21oi_1 _22729_ (.A1(_12803_),
    .A2(_12805_),
    .B1(_12807_),
    .Y(_12808_));
 sky130_fd_sc_hd__a21o_1 _22730_ (.A1(_12803_),
    .A2(_12805_),
    .B1(_12807_),
    .X(_12809_));
 sky130_fd_sc_hd__and3_1 _22731_ (.A(_12803_),
    .B(_12805_),
    .C(_12807_),
    .X(_12810_));
 sky130_fd_sc_hd__nand3_1 _22732_ (.A(_12803_),
    .B(_12805_),
    .C(_12807_),
    .Y(_12811_));
 sky130_fd_sc_hd__nand2_1 _22733_ (.A(_12809_),
    .B(_12811_),
    .Y(_12813_));
 sky130_fd_sc_hd__o211ai_2 _22734_ (.A1(_12808_),
    .A2(_12810_),
    .B1(_12775_),
    .C1(_12777_),
    .Y(_12814_));
 sky130_fd_sc_hd__a21o_1 _22735_ (.A1(_12775_),
    .A2(_12777_),
    .B1(_12813_),
    .X(_12815_));
 sky130_fd_sc_hd__o2bb2ai_1 _22736_ (.A1_N(_12775_),
    .A2_N(_12777_),
    .B1(_12808_),
    .B2(_12810_),
    .Y(_12816_));
 sky130_fd_sc_hd__and3_1 _22737_ (.A(_12777_),
    .B(_12809_),
    .C(_12811_),
    .X(_12817_));
 sky130_fd_sc_hd__nand4_2 _22738_ (.A(_12775_),
    .B(_12777_),
    .C(_12809_),
    .D(_12811_),
    .Y(_12818_));
 sky130_fd_sc_hd__nand4_4 _22739_ (.A(_12583_),
    .B(_12733_),
    .C(_12816_),
    .D(_12818_),
    .Y(_12819_));
 sky130_fd_sc_hd__inv_2 _22740_ (.A(_12819_),
    .Y(_12820_));
 sky130_fd_sc_hd__o211a_1 _22741_ (.A1(_12581_),
    .A2(_12732_),
    .B1(_12814_),
    .C1(_12815_),
    .X(_12821_));
 sky130_fd_sc_hd__o211ai_2 _22742_ (.A1(_12581_),
    .A2(_12732_),
    .B1(_12814_),
    .C1(_12815_),
    .Y(_12822_));
 sky130_fd_sc_hd__o22a_1 _22743_ (.A1(_12680_),
    .A2(_12682_),
    .B1(_12641_),
    .B2(_12644_),
    .X(_12824_));
 sky130_fd_sc_hd__o2bb2a_1 _22744_ (.A1_N(_12684_),
    .A2_N(_12642_),
    .B1(_12641_),
    .B2(_12644_),
    .X(_12825_));
 sky130_fd_sc_hd__a21oi_1 _22745_ (.A1(_12819_),
    .A2(_12822_),
    .B1(_12825_),
    .Y(_12826_));
 sky130_fd_sc_hd__and3_1 _22746_ (.A(_12819_),
    .B(_12822_),
    .C(_12825_),
    .X(_12827_));
 sky130_fd_sc_hd__o2bb2ai_1 _22747_ (.A1_N(_12819_),
    .A2_N(_12822_),
    .B1(_12824_),
    .B2(_12643_),
    .Y(_12828_));
 sky130_fd_sc_hd__nand3b_1 _22748_ (.A_N(_12825_),
    .B(_12822_),
    .C(_12819_),
    .Y(_12829_));
 sky130_fd_sc_hd__nand2_1 _22749_ (.A(_12828_),
    .B(_12829_),
    .Y(_12830_));
 sky130_fd_sc_hd__nand3_2 _22750_ (.A(_12500_),
    .B(_12585_),
    .C(_12587_),
    .Y(_12831_));
 sky130_fd_sc_hd__nand3_1 _22751_ (.A(_12499_),
    .B(_12589_),
    .C(_12591_),
    .Y(_12832_));
 sky130_fd_sc_hd__o311a_1 _22752_ (.A1(_11813_),
    .A2(_12032_),
    .A3(_12035_),
    .B1(_12057_),
    .C1(_12487_),
    .X(_12833_));
 sky130_fd_sc_hd__o21ai_4 _22753_ (.A1(_12490_),
    .A2(_12488_),
    .B1(_12487_),
    .Y(_12835_));
 sky130_fd_sc_hd__a31o_2 _22754_ (.A1(_12038_),
    .A2(_12057_),
    .A3(_12487_),
    .B1(_12488_),
    .X(_12836_));
 sky130_fd_sc_hd__o22a_1 _22755_ (.A1(_05077_),
    .A2(_05463_),
    .B1(_05465_),
    .B2(_04113_),
    .X(_12837_));
 sky130_fd_sc_hd__nand3_2 _22756_ (.A(net182),
    .B(net179),
    .C(_05225_),
    .Y(_12838_));
 sky130_fd_sc_hd__or3_2 _22757_ (.A(net46),
    .B(_04135_),
    .C(_04124_),
    .X(_12839_));
 sky130_fd_sc_hd__or3_1 _22758_ (.A(net45),
    .B(_04146_),
    .C(_04102_),
    .X(_12840_));
 sky130_fd_sc_hd__o211ai_4 _22759_ (.A1(net184),
    .A2(_05551_),
    .B1(net242),
    .C1(net178),
    .Y(_12841_));
 sky130_fd_sc_hd__o2111a_1 _22760_ (.A1(_04146_),
    .A2(_04989_),
    .B1(_12838_),
    .C1(_12839_),
    .D1(_12841_),
    .X(_12842_));
 sky130_fd_sc_hd__o2111ai_4 _22761_ (.A1(_04146_),
    .A2(_04989_),
    .B1(_12838_),
    .C1(_12839_),
    .D1(_12841_),
    .Y(_12843_));
 sky130_fd_sc_hd__a22oi_1 _22762_ (.A1(_12838_),
    .A2(_12839_),
    .B1(_12840_),
    .B2(_12841_),
    .Y(_12844_));
 sky130_fd_sc_hd__a22o_1 _22763_ (.A1(_12838_),
    .A2(_12839_),
    .B1(_12840_),
    .B2(_12841_),
    .X(_12846_));
 sky130_fd_sc_hd__nand2_1 _22764_ (.A(_12846_),
    .B(_12837_),
    .Y(_12847_));
 sky130_fd_sc_hd__nand3b_1 _22765_ (.A_N(_12837_),
    .B(_12843_),
    .C(_12846_),
    .Y(_12848_));
 sky130_fd_sc_hd__o21ai_2 _22766_ (.A1(_12837_),
    .A2(_12842_),
    .B1(_12846_),
    .Y(_12849_));
 sky130_fd_sc_hd__o21ai_1 _22767_ (.A1(_12842_),
    .A2(_12844_),
    .B1(_12837_),
    .Y(_12850_));
 sky130_fd_sc_hd__nand2_1 _22768_ (.A(_12848_),
    .B(_12850_),
    .Y(_12851_));
 sky130_fd_sc_hd__a21o_1 _22769_ (.A1(_12534_),
    .A2(_12542_),
    .B1(_12539_),
    .X(_12852_));
 sky130_fd_sc_hd__a32o_1 _22770_ (.A1(_05933_),
    .A2(_04895_),
    .A3(net174),
    .B1(_04897_),
    .B2(net16),
    .X(_12853_));
 sky130_fd_sc_hd__o211ai_2 _22771_ (.A1(net174),
    .A2(_06451_),
    .B1(_04267_),
    .C1(net198),
    .Y(_12854_));
 sky130_fd_sc_hd__or3b_1 _22772_ (.A(net41),
    .B(_04179_),
    .C_N(net40),
    .X(_12855_));
 sky130_fd_sc_hd__a32oi_4 _22773_ (.A1(net202),
    .A2(net173),
    .A3(net279),
    .B1(_04482_),
    .B2(net17),
    .Y(_12857_));
 sky130_fd_sc_hd__a21oi_2 _22774_ (.A1(_12854_),
    .A2(_12855_),
    .B1(_12857_),
    .Y(_12858_));
 sky130_fd_sc_hd__a21o_1 _22775_ (.A1(_12854_),
    .A2(_12855_),
    .B1(_12857_),
    .X(_12859_));
 sky130_fd_sc_hd__o211a_1 _22776_ (.A1(_04179_),
    .A2(_04270_),
    .B1(_12854_),
    .C1(_12857_),
    .X(_12860_));
 sky130_fd_sc_hd__o221ai_4 _22777_ (.A1(_04179_),
    .A2(_04270_),
    .B1(_06454_),
    .B2(_04268_),
    .C1(_12857_),
    .Y(_12861_));
 sky130_fd_sc_hd__nand3_2 _22778_ (.A(_12853_),
    .B(_12859_),
    .C(_12861_),
    .Y(_12862_));
 sky130_fd_sc_hd__inv_2 _22779_ (.A(_12862_),
    .Y(_12863_));
 sky130_fd_sc_hd__o21bai_2 _22780_ (.A1(_12858_),
    .A2(_12860_),
    .B1_N(_12853_),
    .Y(_12864_));
 sky130_fd_sc_hd__nand2_1 _22781_ (.A(_12852_),
    .B(_12864_),
    .Y(_12865_));
 sky130_fd_sc_hd__and3_2 _22782_ (.A(_12864_),
    .B(_12852_),
    .C(_12862_),
    .X(_12866_));
 sky130_fd_sc_hd__a21oi_2 _22783_ (.A1(_12862_),
    .A2(_12864_),
    .B1(_12852_),
    .Y(_12868_));
 sky130_fd_sc_hd__a21o_1 _22784_ (.A1(_12862_),
    .A2(_12864_),
    .B1(_12852_),
    .X(_12869_));
 sky130_fd_sc_hd__nand3_2 _22785_ (.A(_12848_),
    .B(_12850_),
    .C(_12869_),
    .Y(_12870_));
 sky130_fd_sc_hd__nor2_1 _22786_ (.A(_12866_),
    .B(_12870_),
    .Y(_12871_));
 sky130_fd_sc_hd__o21ai_2 _22787_ (.A1(_12866_),
    .A2(_12868_),
    .B1(_12851_),
    .Y(_12872_));
 sky130_fd_sc_hd__inv_2 _22788_ (.A(_12872_),
    .Y(_12873_));
 sky130_fd_sc_hd__o21ai_1 _22789_ (.A1(_12866_),
    .A2(_12870_),
    .B1(_12872_),
    .Y(_12874_));
 sky130_fd_sc_hd__o2bb2ai_4 _22790_ (.A1_N(_12522_),
    .A2_N(_12525_),
    .B1(_12523_),
    .B2(_12518_),
    .Y(_12875_));
 sky130_fd_sc_hd__a21oi_4 _22791_ (.A1(_12511_),
    .A2(_12514_),
    .B1(_12510_),
    .Y(_12876_));
 sky130_fd_sc_hd__a32o_1 _22792_ (.A1(net194),
    .A2(net171),
    .A3(net281),
    .B1(_04217_),
    .B2(net19),
    .X(_12877_));
 sky130_fd_sc_hd__or3b_2 _22793_ (.A(net38),
    .B(_04223_),
    .C_N(net37),
    .X(_12879_));
 sky130_fd_sc_hd__nand3_4 _22794_ (.A(_07499_),
    .B(net167),
    .C(_02858_),
    .Y(_12880_));
 sky130_fd_sc_hd__o211ai_4 _22795_ (.A1(net174),
    .A2(_07074_),
    .B1(_03704_),
    .C1(_07072_),
    .Y(_12881_));
 sky130_fd_sc_hd__or3_4 _22796_ (.A(net39),
    .B(_04212_),
    .C(_04037_),
    .X(_12882_));
 sky130_fd_sc_hd__o2111a_1 _22797_ (.A1(_04223_),
    .A2(_02891_),
    .B1(_12880_),
    .C1(_12881_),
    .D1(_12882_),
    .X(_12883_));
 sky130_fd_sc_hd__o2111ai_4 _22798_ (.A1(_04223_),
    .A2(_02891_),
    .B1(_12880_),
    .C1(_12881_),
    .D1(_12882_),
    .Y(_12884_));
 sky130_fd_sc_hd__a22oi_4 _22799_ (.A1(_12879_),
    .A2(_12880_),
    .B1(_12881_),
    .B2(_12882_),
    .Y(_12885_));
 sky130_fd_sc_hd__a22o_1 _22800_ (.A1(_12879_),
    .A2(_12880_),
    .B1(_12881_),
    .B2(_12882_),
    .X(_12886_));
 sky130_fd_sc_hd__o21bai_4 _22801_ (.A1(_12883_),
    .A2(_12885_),
    .B1_N(_12877_),
    .Y(_12887_));
 sky130_fd_sc_hd__and3_2 _22802_ (.A(_12877_),
    .B(_12884_),
    .C(_12886_),
    .X(_12888_));
 sky130_fd_sc_hd__nand3_4 _22803_ (.A(_12877_),
    .B(_12884_),
    .C(_12886_),
    .Y(_12890_));
 sky130_fd_sc_hd__nor2_1 _22804_ (.A(_12464_),
    .B(_12471_),
    .Y(_12891_));
 sky130_fd_sc_hd__a31oi_4 _22805_ (.A1(_12467_),
    .A2(_12468_),
    .A3(_12469_),
    .B1(_12463_),
    .Y(_12892_));
 sky130_fd_sc_hd__o32a_1 _22806_ (.A1(_12465_),
    .A2(_12466_),
    .A3(_12470_),
    .B1(_12464_),
    .B2(_12471_),
    .X(_12893_));
 sky130_fd_sc_hd__a21oi_4 _22807_ (.A1(_12887_),
    .A2(_12890_),
    .B1(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__o2bb2ai_2 _22808_ (.A1_N(_12887_),
    .A2_N(_12890_),
    .B1(_12891_),
    .B2(_12474_),
    .Y(_12895_));
 sky130_fd_sc_hd__o21ai_2 _22809_ (.A1(_12471_),
    .A2(_12892_),
    .B1(_12887_),
    .Y(_12896_));
 sky130_fd_sc_hd__o211a_1 _22810_ (.A1(_12471_),
    .A2(_12892_),
    .B1(_12890_),
    .C1(_12887_),
    .X(_12897_));
 sky130_fd_sc_hd__o211ai_2 _22811_ (.A1(_12471_),
    .A2(_12892_),
    .B1(_12890_),
    .C1(_12887_),
    .Y(_12898_));
 sky130_fd_sc_hd__a31o_1 _22812_ (.A1(_12887_),
    .A2(_12890_),
    .A3(_12893_),
    .B1(_12876_),
    .X(_12899_));
 sky130_fd_sc_hd__o221a_1 _22813_ (.A1(_12510_),
    .A2(_12518_),
    .B1(_12888_),
    .B2(_12896_),
    .C1(_12895_),
    .X(_12901_));
 sky130_fd_sc_hd__o221ai_4 _22814_ (.A1(_12510_),
    .A2(_12518_),
    .B1(_12888_),
    .B2(_12896_),
    .C1(_12895_),
    .Y(_12902_));
 sky130_fd_sc_hd__a21boi_1 _22815_ (.A1(_12895_),
    .A2(_12898_),
    .B1_N(_12876_),
    .Y(_12903_));
 sky130_fd_sc_hd__o21ai_4 _22816_ (.A1(_12894_),
    .A2(_12897_),
    .B1(_12876_),
    .Y(_12904_));
 sky130_fd_sc_hd__o211a_2 _22817_ (.A1(_12899_),
    .A2(_12894_),
    .B1(_12875_),
    .C1(_12904_),
    .X(_12905_));
 sky130_fd_sc_hd__o211ai_4 _22818_ (.A1(_12894_),
    .A2(_12899_),
    .B1(_12904_),
    .C1(_12875_),
    .Y(_12906_));
 sky130_fd_sc_hd__a21oi_4 _22819_ (.A1(_12902_),
    .A2(_12904_),
    .B1(_12875_),
    .Y(_12907_));
 sky130_fd_sc_hd__o21bai_4 _22820_ (.A1(_12901_),
    .A2(_12903_),
    .B1_N(_12875_),
    .Y(_12908_));
 sky130_fd_sc_hd__o21bai_2 _22821_ (.A1(_12905_),
    .A2(_12907_),
    .B1_N(_12874_),
    .Y(_12909_));
 sky130_fd_sc_hd__nand2_1 _22822_ (.A(_12874_),
    .B(_12906_),
    .Y(_12910_));
 sky130_fd_sc_hd__o211ai_2 _22823_ (.A1(_12871_),
    .A2(_12873_),
    .B1(_12906_),
    .C1(_12908_),
    .Y(_12912_));
 sky130_fd_sc_hd__o211a_1 _22824_ (.A1(_12866_),
    .A2(_12870_),
    .B1(_12872_),
    .C1(_12908_),
    .X(_12913_));
 sky130_fd_sc_hd__o2111ai_4 _22825_ (.A1(_12866_),
    .A2(_12870_),
    .B1(_12872_),
    .C1(_12906_),
    .D1(_12908_),
    .Y(_12914_));
 sky130_fd_sc_hd__o22ai_4 _22826_ (.A1(_12871_),
    .A2(_12873_),
    .B1(_12905_),
    .B2(_12907_),
    .Y(_12915_));
 sky130_fd_sc_hd__and3_1 _22827_ (.A(_12915_),
    .B(_12835_),
    .C(_12914_),
    .X(_12916_));
 sky130_fd_sc_hd__nand3_4 _22828_ (.A(_12915_),
    .B(_12835_),
    .C(_12914_),
    .Y(_12917_));
 sky130_fd_sc_hd__a2bb2oi_1 _22829_ (.A1_N(_12488_),
    .A2_N(_12833_),
    .B1(_12914_),
    .B2(_12915_),
    .Y(_12918_));
 sky130_fd_sc_hd__o211ai_1 _22830_ (.A1(_12910_),
    .A2(_12907_),
    .B1(_12836_),
    .C1(_12909_),
    .Y(_12919_));
 sky130_fd_sc_hd__a31oi_4 _22831_ (.A1(_12836_),
    .A2(_12909_),
    .A3(_12912_),
    .B1(_12575_),
    .Y(_12920_));
 sky130_fd_sc_hd__nand2_2 _22832_ (.A(_12920_),
    .B(_12917_),
    .Y(_12921_));
 sky130_fd_sc_hd__a21o_1 _22833_ (.A1(_12917_),
    .A2(_12919_),
    .B1(_12576_),
    .X(_12923_));
 sky130_fd_sc_hd__a211o_1 _22834_ (.A1(_12909_),
    .A2(_12912_),
    .B1(_12575_),
    .C1(_12836_),
    .X(_12924_));
 sky130_fd_sc_hd__o2111ai_1 _22835_ (.A1(_12910_),
    .A2(_12907_),
    .B1(_12836_),
    .C1(_12575_),
    .D1(_12909_),
    .Y(_12925_));
 sky130_fd_sc_hd__a31oi_1 _22836_ (.A1(_12915_),
    .A2(_12835_),
    .A3(_12914_),
    .B1(_12576_),
    .Y(_12926_));
 sky130_fd_sc_hd__a21oi_1 _22837_ (.A1(_12576_),
    .A2(_12919_),
    .B1(_12916_),
    .Y(_12927_));
 sky130_fd_sc_hd__o21ai_2 _22838_ (.A1(_12918_),
    .A2(_12926_),
    .B1(_12925_),
    .Y(_12928_));
 sky130_fd_sc_hd__nand3_2 _22839_ (.A(_12447_),
    .B(_12491_),
    .C(_12492_),
    .Y(_12929_));
 sky130_fd_sc_hd__nand2_1 _22840_ (.A(_12445_),
    .B(_12929_),
    .Y(_12930_));
 sky130_fd_sc_hd__a31oi_2 _22841_ (.A1(_12429_),
    .A2(_12430_),
    .A3(_12432_),
    .B1(_12099_),
    .Y(_12931_));
 sky130_fd_sc_hd__o21ai_2 _22842_ (.A1(_12098_),
    .A2(_12433_),
    .B1(_12435_),
    .Y(_12932_));
 sky130_fd_sc_hd__a32oi_4 _22843_ (.A1(_12419_),
    .A2(_12408_),
    .A3(_12418_),
    .B1(net134),
    .B2(net138),
    .Y(_12934_));
 sky130_fd_sc_hd__o21ai_2 _22844_ (.A1(_10546_),
    .A2(_12424_),
    .B1(_12423_),
    .Y(_12935_));
 sky130_fd_sc_hd__a21oi_1 _22845_ (.A1(net133),
    .A2(_12425_),
    .B1(_12422_),
    .Y(_12936_));
 sky130_fd_sc_hd__o21ai_2 _22846_ (.A1(_12410_),
    .A2(_08878_),
    .B1(net147),
    .Y(_12937_));
 sky130_fd_sc_hd__a31o_1 _22847_ (.A1(net307),
    .A2(net296),
    .A3(net287),
    .B1(_08658_),
    .X(_12938_));
 sky130_fd_sc_hd__o22ai_4 _22848_ (.A1(_03982_),
    .A2(_08660_),
    .B1(_11343_),
    .B2(_12938_),
    .Y(_12939_));
 sky130_fd_sc_hd__o2111a_2 _22849_ (.A1(net169),
    .A2(net268),
    .B1(net33),
    .C1(_12939_),
    .D1(net319),
    .X(_12940_));
 sky130_fd_sc_hd__o2111ai_4 _22850_ (.A1(net169),
    .A2(net268),
    .B1(net33),
    .C1(_12939_),
    .D1(net319),
    .Y(_12941_));
 sky130_fd_sc_hd__a31oi_4 _22851_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_12939_),
    .Y(_12942_));
 sky130_fd_sc_hd__a31o_1 _22852_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_12939_),
    .X(_12943_));
 sky130_fd_sc_hd__nand3_2 _22853_ (.A(_12943_),
    .B(net147),
    .C(_12941_),
    .Y(_12945_));
 sky130_fd_sc_hd__o22ai_4 _22854_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_12940_),
    .B2(_12942_),
    .Y(_12946_));
 sky130_fd_sc_hd__o21ai_4 _22855_ (.A1(_12940_),
    .A2(_12942_),
    .B1(net146),
    .Y(_12947_));
 sky130_fd_sc_hd__a21oi_1 _22856_ (.A1(_08882_),
    .A2(_09298_),
    .B1(_12942_),
    .Y(_12948_));
 sky130_fd_sc_hd__o21ai_4 _22857_ (.A1(_12939_),
    .A2(net156),
    .B1(_09300_),
    .Y(_12949_));
 sky130_fd_sc_hd__o221a_1 _22858_ (.A1(net156),
    .A2(_12411_),
    .B1(_12942_),
    .B2(net146),
    .C1(_12937_),
    .X(_12950_));
 sky130_fd_sc_hd__a2bb2oi_2 _22859_ (.A1_N(_12414_),
    .A2_N(_12416_),
    .B1(_12945_),
    .B2(_12946_),
    .Y(_12951_));
 sky130_fd_sc_hd__nand2_1 _22860_ (.A(_12950_),
    .B(_12947_),
    .Y(_12952_));
 sky130_fd_sc_hd__a22oi_4 _22861_ (.A1(_12413_),
    .A2(_12937_),
    .B1(_12947_),
    .B2(_12949_),
    .Y(_12953_));
 sky130_fd_sc_hd__nand4_4 _22862_ (.A(_12415_),
    .B(_12418_),
    .C(_12945_),
    .D(_12946_),
    .Y(_12954_));
 sky130_fd_sc_hd__nand3_1 _22863_ (.A(net133),
    .B(_12952_),
    .C(_12954_),
    .Y(_12956_));
 sky130_fd_sc_hd__o22ai_2 _22864_ (.A1(_10540_),
    .A2(net135),
    .B1(_12951_),
    .B2(_12953_),
    .Y(_12957_));
 sky130_fd_sc_hd__o211ai_4 _22865_ (.A1(_10540_),
    .A2(net135),
    .B1(_12952_),
    .C1(_12954_),
    .Y(_12958_));
 sky130_fd_sc_hd__o21ai_4 _22866_ (.A1(_12951_),
    .A2(_12953_),
    .B1(net133),
    .Y(_12959_));
 sky130_fd_sc_hd__and3_2 _22867_ (.A(_12935_),
    .B(_12956_),
    .C(_12957_),
    .X(_12960_));
 sky130_fd_sc_hd__nand3_2 _22868_ (.A(_12935_),
    .B(_12956_),
    .C(_12957_),
    .Y(_12961_));
 sky130_fd_sc_hd__o211a_1 _22869_ (.A1(_12424_),
    .A2(_12934_),
    .B1(_12958_),
    .C1(_12959_),
    .X(_12962_));
 sky130_fd_sc_hd__o211ai_4 _22870_ (.A1(_12424_),
    .A2(_12934_),
    .B1(_12958_),
    .C1(_12959_),
    .Y(_12963_));
 sky130_fd_sc_hd__o2bb2ai_1 _22871_ (.A1_N(_12961_),
    .A2_N(_12963_),
    .B1(_11042_),
    .B2(_11742_),
    .Y(_12964_));
 sky130_fd_sc_hd__o2111ai_4 _22872_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net142),
    .C1(_12961_),
    .D1(_12963_),
    .Y(_12965_));
 sky130_fd_sc_hd__a21o_1 _22873_ (.A1(_12961_),
    .A2(_12963_),
    .B1(_12099_),
    .X(_12967_));
 sky130_fd_sc_hd__a31oi_2 _22874_ (.A1(_12936_),
    .A2(_12958_),
    .A3(_12959_),
    .B1(_12098_),
    .Y(_12968_));
 sky130_fd_sc_hd__a31o_1 _22875_ (.A1(_12936_),
    .A2(_12958_),
    .A3(_12959_),
    .B1(net132),
    .X(_12969_));
 sky130_fd_sc_hd__o211ai_4 _22876_ (.A1(_12433_),
    .A2(_12931_),
    .B1(_12964_),
    .C1(_12965_),
    .Y(_12970_));
 sky130_fd_sc_hd__o211ai_4 _22877_ (.A1(_12960_),
    .A2(_12969_),
    .B1(_12932_),
    .C1(_12967_),
    .Y(_12971_));
 sky130_fd_sc_hd__nor2_2 _22878_ (.A(_04245_),
    .B(_01326_),
    .Y(_12972_));
 sky130_fd_sc_hd__o311a_1 _22879_ (.A1(_03958_),
    .A2(_05927_),
    .A3(_07767_),
    .B1(_07771_),
    .C1(_01293_),
    .X(_12973_));
 sky130_fd_sc_hd__a31oi_2 _22880_ (.A1(_07771_),
    .A2(_01293_),
    .A3(net165),
    .B1(_12972_),
    .Y(_12974_));
 sky130_fd_sc_hd__a31o_1 _22881_ (.A1(_07771_),
    .A2(_01293_),
    .A3(net165),
    .B1(_12972_),
    .X(_12975_));
 sky130_fd_sc_hd__a211oi_2 _22882_ (.A1(_07075_),
    .A2(_08205_),
    .B1(_12341_),
    .C1(_08203_),
    .Y(_12976_));
 sky130_fd_sc_hd__nor2_2 _22883_ (.A(_04256_),
    .B(_12363_),
    .Y(_12978_));
 sky130_fd_sc_hd__a31oi_4 _22884_ (.A1(net164),
    .A2(net161),
    .A3(_12330_),
    .B1(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__and3_2 _22885_ (.A(_03993_),
    .B(net25),
    .C(net34),
    .X(_12980_));
 sky130_fd_sc_hd__or3_1 _22886_ (.A(net35),
    .B(net319),
    .C(_03971_),
    .X(_12981_));
 sky130_fd_sc_hd__a21oi_1 _22887_ (.A1(net150),
    .A2(_08668_),
    .B1(_11782_),
    .Y(_12982_));
 sky130_fd_sc_hd__o21ai_2 _22888_ (.A1(net159),
    .A2(_08666_),
    .B1(net252),
    .Y(_12983_));
 sky130_fd_sc_hd__o311a_1 _22889_ (.A1(_03971_),
    .A2(net35),
    .A3(net319),
    .B1(_12979_),
    .C1(_12983_),
    .X(_12984_));
 sky130_fd_sc_hd__o211ai_4 _22890_ (.A1(net319),
    .A2(_11804_),
    .B1(_12979_),
    .C1(_12983_),
    .Y(_12985_));
 sky130_fd_sc_hd__o22a_2 _22891_ (.A1(_12976_),
    .A2(_12978_),
    .B1(_12980_),
    .B2(_12982_),
    .X(_12986_));
 sky130_fd_sc_hd__o22ai_2 _22892_ (.A1(_12976_),
    .A2(_12978_),
    .B1(_12980_),
    .B2(_12982_),
    .Y(_12987_));
 sky130_fd_sc_hd__o211ai_2 _22893_ (.A1(_12972_),
    .A2(_12973_),
    .B1(_12985_),
    .C1(_12987_),
    .Y(_12989_));
 sky130_fd_sc_hd__o21ai_1 _22894_ (.A1(_12984_),
    .A2(_12986_),
    .B1(_12974_),
    .Y(_12990_));
 sky130_fd_sc_hd__o22ai_2 _22895_ (.A1(_12972_),
    .A2(_12973_),
    .B1(_12984_),
    .B2(_12986_),
    .Y(_12991_));
 sky130_fd_sc_hd__nand3_1 _22896_ (.A(_12987_),
    .B(_12974_),
    .C(_12985_),
    .Y(_12992_));
 sky130_fd_sc_hd__o211ai_4 _22897_ (.A1(_12451_),
    .A2(_12457_),
    .B1(_12989_),
    .C1(_12990_),
    .Y(_12993_));
 sky130_fd_sc_hd__nand4_4 _22898_ (.A(_12991_),
    .B(_12449_),
    .C(_12458_),
    .D(_12992_),
    .Y(_12994_));
 sky130_fd_sc_hd__a21oi_4 _22899_ (.A1(_12993_),
    .A2(_12994_),
    .B1(_11740_),
    .Y(_12995_));
 sky130_fd_sc_hd__a22o_1 _22900_ (.A1(net137),
    .A2(_11736_),
    .B1(_12993_),
    .B2(_12994_),
    .X(_12996_));
 sky130_fd_sc_hd__and3_1 _22901_ (.A(_12993_),
    .B(_12994_),
    .C(_11740_),
    .X(_12997_));
 sky130_fd_sc_hd__o2111ai_4 _22902_ (.A1(_11527_),
    .A2(_11732_),
    .B1(_12994_),
    .C1(net137),
    .D1(_12993_),
    .Y(_12998_));
 sky130_fd_sc_hd__a31o_2 _22903_ (.A1(_12459_),
    .A2(_12479_),
    .A3(_12481_),
    .B1(_12460_),
    .X(_13000_));
 sky130_fd_sc_hd__a21oi_1 _22904_ (.A1(_12996_),
    .A2(_12998_),
    .B1(_13000_),
    .Y(_13001_));
 sky130_fd_sc_hd__and3_1 _22905_ (.A(_12996_),
    .B(_12998_),
    .C(_13000_),
    .X(_13002_));
 sky130_fd_sc_hd__a21boi_1 _22906_ (.A1(_12996_),
    .A2(_12998_),
    .B1_N(_13000_),
    .Y(_13003_));
 sky130_fd_sc_hd__o21ai_1 _22907_ (.A1(_12995_),
    .A2(_12997_),
    .B1(_13000_),
    .Y(_13004_));
 sky130_fd_sc_hd__a311oi_2 _22908_ (.A1(_11740_),
    .A2(_12993_),
    .A3(_12994_),
    .B1(_13000_),
    .C1(_12995_),
    .Y(_13005_));
 sky130_fd_sc_hd__nand3b_1 _22909_ (.A_N(_13000_),
    .B(_12998_),
    .C(_12996_),
    .Y(_13006_));
 sky130_fd_sc_hd__o211ai_2 _22910_ (.A1(_13003_),
    .A2(_13005_),
    .B1(_12970_),
    .C1(_12971_),
    .Y(_13007_));
 sky130_fd_sc_hd__o2bb2ai_1 _22911_ (.A1_N(_12970_),
    .A2_N(_12971_),
    .B1(_13001_),
    .B2(_13002_),
    .Y(_13008_));
 sky130_fd_sc_hd__o2bb2ai_2 _22912_ (.A1_N(_12970_),
    .A2_N(_12971_),
    .B1(_13003_),
    .B2(_13005_),
    .Y(_13009_));
 sky130_fd_sc_hd__nand3_1 _22913_ (.A(_12970_),
    .B(_13004_),
    .C(_13006_),
    .Y(_13011_));
 sky130_fd_sc_hd__nand4_2 _22914_ (.A(_12970_),
    .B(_12971_),
    .C(_13004_),
    .D(_13006_),
    .Y(_13012_));
 sky130_fd_sc_hd__a22oi_4 _22915_ (.A1(_12445_),
    .A2(_12929_),
    .B1(_13009_),
    .B2(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__a22o_2 _22916_ (.A1(_12445_),
    .A2(_12929_),
    .B1(_13009_),
    .B2(_13012_),
    .X(_13014_));
 sky130_fd_sc_hd__a21oi_2 _22917_ (.A1(_13007_),
    .A2(_13008_),
    .B1(_12930_),
    .Y(_13015_));
 sky130_fd_sc_hd__a21o_2 _22918_ (.A1(_13007_),
    .A2(_13008_),
    .B1(_12930_),
    .X(_13016_));
 sky130_fd_sc_hd__o2111ai_1 _22919_ (.A1(_12917_),
    .A2(_12575_),
    .B1(_13014_),
    .C1(_12928_),
    .D1(_13016_),
    .Y(_13017_));
 sky130_fd_sc_hd__o211ai_1 _22920_ (.A1(_13013_),
    .A2(_13015_),
    .B1(_12921_),
    .C1(_12923_),
    .Y(_13018_));
 sky130_fd_sc_hd__and4_1 _22921_ (.A(_12921_),
    .B(_12923_),
    .C(_13014_),
    .D(_13016_),
    .X(_13019_));
 sky130_fd_sc_hd__nand4_4 _22922_ (.A(_12921_),
    .B(_12923_),
    .C(_13014_),
    .D(_13016_),
    .Y(_13020_));
 sky130_fd_sc_hd__o221ai_4 _22923_ (.A1(_12575_),
    .A2(_12917_),
    .B1(_13013_),
    .B2(_13015_),
    .C1(_12928_),
    .Y(_13022_));
 sky130_fd_sc_hd__nand3_1 _22924_ (.A(_12499_),
    .B(_12831_),
    .C(_13022_),
    .Y(_13023_));
 sky130_fd_sc_hd__a22oi_2 _22925_ (.A1(_12500_),
    .A2(_12832_),
    .B1(_13017_),
    .B2(_13018_),
    .Y(_13024_));
 sky130_fd_sc_hd__nand4_1 _22926_ (.A(_12499_),
    .B(_12831_),
    .C(_13020_),
    .D(_13022_),
    .Y(_13025_));
 sky130_fd_sc_hd__a22oi_4 _22927_ (.A1(_12499_),
    .A2(_12831_),
    .B1(_13020_),
    .B2(_13022_),
    .Y(_13026_));
 sky130_fd_sc_hd__a22o_1 _22928_ (.A1(_12499_),
    .A2(_12831_),
    .B1(_13020_),
    .B2(_13022_),
    .X(_13027_));
 sky130_fd_sc_hd__o211ai_1 _22929_ (.A1(_13019_),
    .A2(_13023_),
    .B1(_12830_),
    .C1(_13027_),
    .Y(_13028_));
 sky130_fd_sc_hd__o22ai_1 _22930_ (.A1(_12826_),
    .A2(_12827_),
    .B1(_13024_),
    .B2(_13026_),
    .Y(_13029_));
 sky130_fd_sc_hd__o211ai_2 _22931_ (.A1(_12826_),
    .A2(_12827_),
    .B1(_13025_),
    .C1(_13027_),
    .Y(_13030_));
 sky130_fd_sc_hd__o2bb2ai_1 _22932_ (.A1_N(_12828_),
    .A2_N(_12829_),
    .B1(_13024_),
    .B2(_13026_),
    .Y(_13031_));
 sky130_fd_sc_hd__o211a_1 _22933_ (.A1(_12598_),
    .A2(_12701_),
    .B1(_13030_),
    .C1(_13031_),
    .X(_13033_));
 sky130_fd_sc_hd__o211ai_2 _22934_ (.A1(_12598_),
    .A2(_12701_),
    .B1(_13030_),
    .C1(_13031_),
    .Y(_13034_));
 sky130_fd_sc_hd__nand3_2 _22935_ (.A(_12731_),
    .B(_13028_),
    .C(_13029_),
    .Y(_13035_));
 sky130_fd_sc_hd__o21ai_1 _22936_ (.A1(_12690_),
    .A2(_12695_),
    .B1(_13035_),
    .Y(_13036_));
 sky130_fd_sc_hd__o211a_1 _22937_ (.A1(_12690_),
    .A2(_12695_),
    .B1(_13034_),
    .C1(_13035_),
    .X(_13037_));
 sky130_fd_sc_hd__a21oi_1 _22938_ (.A1(_13034_),
    .A2(_13035_),
    .B1(_12730_),
    .Y(_13038_));
 sky130_fd_sc_hd__a21o_1 _22939_ (.A1(_13034_),
    .A2(_13035_),
    .B1(_12730_),
    .X(_13039_));
 sky130_fd_sc_hd__o21ai_2 _22940_ (.A1(_12708_),
    .A2(_12704_),
    .B1(_12707_),
    .Y(_13040_));
 sky130_fd_sc_hd__o21a_1 _22941_ (.A1(_12708_),
    .A2(_12704_),
    .B1(_12707_),
    .X(_13041_));
 sky130_fd_sc_hd__o21a_1 _22942_ (.A1(_13037_),
    .A2(_13038_),
    .B1(_13041_),
    .X(_13042_));
 sky130_fd_sc_hd__o21ai_2 _22943_ (.A1(_13037_),
    .A2(_13038_),
    .B1(_13041_),
    .Y(_13044_));
 sky130_fd_sc_hd__o211ai_4 _22944_ (.A1(_13033_),
    .A2(_13036_),
    .B1(_13040_),
    .C1(_13039_),
    .Y(_13045_));
 sky130_fd_sc_hd__a22o_1 _22945_ (.A1(_12679_),
    .A2(_12683_),
    .B1(_13044_),
    .B2(_13045_),
    .X(_13046_));
 sky130_fd_sc_hd__nand4_1 _22946_ (.A(_12679_),
    .B(_12683_),
    .C(_13044_),
    .D(_13045_),
    .Y(_13047_));
 sky130_fd_sc_hd__a21o_1 _22947_ (.A1(_13044_),
    .A2(_13045_),
    .B1(_12729_),
    .X(_13048_));
 sky130_fd_sc_hd__nand2_1 _22948_ (.A(_13044_),
    .B(_12729_),
    .Y(_13049_));
 sky130_fd_sc_hd__nand3_2 _22949_ (.A(_13044_),
    .B(_13045_),
    .C(_12729_),
    .Y(_13050_));
 sky130_fd_sc_hd__nand3b_2 _22950_ (.A_N(_12728_),
    .B(_13046_),
    .C(_13047_),
    .Y(_13051_));
 sky130_fd_sc_hd__nand3_2 _22951_ (.A(_12728_),
    .B(_13048_),
    .C(_13050_),
    .Y(_13052_));
 sky130_fd_sc_hd__nand2_1 _22952_ (.A(_13051_),
    .B(_13052_),
    .Y(_13053_));
 sky130_fd_sc_hd__a31o_1 _22953_ (.A1(_11990_),
    .A2(_12384_),
    .A3(_12386_),
    .B1(_12722_),
    .X(_13055_));
 sky130_fd_sc_hd__o21ai_1 _22954_ (.A1(_13055_),
    .A2(_12726_),
    .B1(_12721_),
    .Y(_13056_));
 sky130_fd_sc_hd__xor2_1 _22955_ (.A(_13053_),
    .B(_13056_),
    .X(net101));
 sky130_fd_sc_hd__a31oi_4 _22956_ (.A1(_12679_),
    .A2(_12683_),
    .A3(_13045_),
    .B1(_13042_),
    .Y(_13057_));
 sky130_fd_sc_hd__a21oi_1 _22957_ (.A1(_12730_),
    .A2(_13035_),
    .B1(_13033_),
    .Y(_13058_));
 sky130_fd_sc_hd__a21o_1 _22958_ (.A1(_12730_),
    .A2(_13035_),
    .B1(_13033_),
    .X(_13059_));
 sky130_fd_sc_hd__o22ai_2 _22959_ (.A1(_13019_),
    .A2(_13023_),
    .B1(_13026_),
    .B2(_12830_),
    .Y(_13060_));
 sky130_fd_sc_hd__o22a_1 _22960_ (.A1(_13019_),
    .A2(_13023_),
    .B1(_13026_),
    .B2(_12830_),
    .X(_13061_));
 sky130_fd_sc_hd__o31a_1 _22961_ (.A1(_10324_),
    .A2(_08668_),
    .A3(_12453_),
    .B1(_12993_),
    .X(_13062_));
 sky130_fd_sc_hd__o21ai_2 _22962_ (.A1(_12452_),
    .A2(_12453_),
    .B1(_12993_),
    .Y(_13063_));
 sky130_fd_sc_hd__o221a_4 _22963_ (.A1(net319),
    .A2(_10346_),
    .B1(net150),
    .B2(_10324_),
    .C1(_12453_),
    .X(_13065_));
 sky130_fd_sc_hd__nand2_8 _22964_ (.A(_12449_),
    .B(_12453_),
    .Y(_13066_));
 sky130_fd_sc_hd__o32a_4 _22965_ (.A1(_01304_),
    .A2(_08203_),
    .A3(net154),
    .B1(_01326_),
    .B2(_04256_),
    .X(_13067_));
 sky130_fd_sc_hd__a32o_1 _22966_ (.A1(net164),
    .A2(net161),
    .A3(_01293_),
    .B1(_01315_),
    .B2(net24),
    .X(_13068_));
 sky130_fd_sc_hd__o21ai_4 _22967_ (.A1(net159),
    .A2(_08666_),
    .B1(_12330_),
    .Y(_13069_));
 sky130_fd_sc_hd__or3_4 _22968_ (.A(net36),
    .B(net319),
    .C(_03993_),
    .X(_13070_));
 sky130_fd_sc_hd__o21ai_1 _22969_ (.A1(net319),
    .A2(_12363_),
    .B1(_13069_),
    .Y(_13071_));
 sky130_fd_sc_hd__and3_1 _22970_ (.A(_03971_),
    .B(net319),
    .C(net35),
    .X(_13072_));
 sky130_fd_sc_hd__a21oi_4 _22971_ (.A1(net161),
    .A2(_13072_),
    .B1(_12980_),
    .Y(_13073_));
 sky130_fd_sc_hd__a31o_1 _22972_ (.A1(net319),
    .A2(net161),
    .A3(net252),
    .B1(_12980_),
    .X(_13074_));
 sky130_fd_sc_hd__a21oi_4 _22973_ (.A1(_13069_),
    .A2(_13070_),
    .B1(_13073_),
    .Y(_13076_));
 sky130_fd_sc_hd__a21o_1 _22974_ (.A1(_13069_),
    .A2(_13070_),
    .B1(_13073_),
    .X(_13077_));
 sky130_fd_sc_hd__o311a_4 _22975_ (.A1(_03993_),
    .A2(net36),
    .A3(net319),
    .B1(_13073_),
    .C1(_13069_),
    .X(_13078_));
 sky130_fd_sc_hd__o21a_1 _22976_ (.A1(_13076_),
    .A2(_13078_),
    .B1(_13067_),
    .X(_13079_));
 sky130_fd_sc_hd__o21ai_4 _22977_ (.A1(_13076_),
    .A2(_13078_),
    .B1(_13067_),
    .Y(_13080_));
 sky130_fd_sc_hd__a31oi_2 _22978_ (.A1(_13069_),
    .A2(_13070_),
    .A3(_13073_),
    .B1(_13067_),
    .Y(_13081_));
 sky130_fd_sc_hd__a31o_1 _22979_ (.A1(_13069_),
    .A2(_13070_),
    .A3(_13073_),
    .B1(_13067_),
    .X(_13082_));
 sky130_fd_sc_hd__a21oi_1 _22980_ (.A1(_13080_),
    .A2(_13082_),
    .B1(_13066_),
    .Y(_13083_));
 sky130_fd_sc_hd__a21o_1 _22981_ (.A1(_13080_),
    .A2(_13082_),
    .B1(_13066_),
    .X(_13084_));
 sky130_fd_sc_hd__o221a_1 _22982_ (.A1(_12451_),
    .A2(_12454_),
    .B1(_13067_),
    .B2(_13078_),
    .C1(_13080_),
    .X(_13085_));
 sky130_fd_sc_hd__o221ai_4 _22983_ (.A1(_12451_),
    .A2(_12454_),
    .B1(_13067_),
    .B2(_13078_),
    .C1(_13080_),
    .Y(_13087_));
 sky130_fd_sc_hd__o32a_2 _22984_ (.A1(_10297_),
    .A2(_10538_),
    .A3(_11735_),
    .B1(_13083_),
    .B2(_13085_),
    .X(_13088_));
 sky130_fd_sc_hd__o21ai_2 _22985_ (.A1(_13083_),
    .A2(_13085_),
    .B1(_11741_),
    .Y(_13089_));
 sky130_fd_sc_hd__and3_1 _22986_ (.A(_13084_),
    .B(_13087_),
    .C(_11740_),
    .X(_13090_));
 sky130_fd_sc_hd__o2111ai_4 _22987_ (.A1(_11527_),
    .A2(_11732_),
    .B1(_13087_),
    .C1(net137),
    .D1(_13084_),
    .Y(_13091_));
 sky130_fd_sc_hd__a21o_2 _22988_ (.A1(_13089_),
    .A2(_13091_),
    .B1(_13063_),
    .X(_13092_));
 sky130_fd_sc_hd__nor2_1 _22989_ (.A(_13062_),
    .B(_13088_),
    .Y(_13093_));
 sky130_fd_sc_hd__nand3_4 _22990_ (.A(_13063_),
    .B(_13089_),
    .C(_13091_),
    .Y(_13094_));
 sky130_fd_sc_hd__a31oi_2 _22991_ (.A1(_12935_),
    .A2(_12956_),
    .A3(_12957_),
    .B1(_12099_),
    .Y(_13095_));
 sky130_fd_sc_hd__o21ai_1 _22992_ (.A1(net132),
    .A2(_12962_),
    .B1(_12961_),
    .Y(_13096_));
 sky130_fd_sc_hd__o311a_1 _22993_ (.A1(_03286_),
    .A2(net44),
    .A3(net319),
    .B1(_09298_),
    .C1(_12941_),
    .X(_13098_));
 sky130_fd_sc_hd__nor2_1 _22994_ (.A(_04004_),
    .B(_08660_),
    .Y(_13099_));
 sky130_fd_sc_hd__a31o_2 _22995_ (.A1(_12977_),
    .A2(_12999_),
    .A3(_08657_),
    .B1(_13099_),
    .X(_13100_));
 sky130_fd_sc_hd__a31oi_4 _22996_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_13100_),
    .Y(_13101_));
 sky130_fd_sc_hd__a31o_1 _22997_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_13100_),
    .X(_13102_));
 sky130_fd_sc_hd__o2111a_1 _22998_ (.A1(net24),
    .A2(net166),
    .B1(net33),
    .C1(_13100_),
    .D1(net319),
    .X(_13103_));
 sky130_fd_sc_hd__o2111ai_4 _22999_ (.A1(net24),
    .A2(net166),
    .B1(net33),
    .C1(_13100_),
    .D1(net319),
    .Y(_13104_));
 sky130_fd_sc_hd__o21ai_1 _23000_ (.A1(_13100_),
    .A2(net156),
    .B1(_09300_),
    .Y(_13105_));
 sky130_fd_sc_hd__o21ai_2 _23001_ (.A1(_13101_),
    .A2(_13103_),
    .B1(net146),
    .Y(_13106_));
 sky130_fd_sc_hd__o22ai_4 _23002_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_13101_),
    .B2(_13103_),
    .Y(_13107_));
 sky130_fd_sc_hd__nand3_2 _23003_ (.A(_13102_),
    .B(_13104_),
    .C(net146),
    .Y(_13109_));
 sky130_fd_sc_hd__a22oi_2 _23004_ (.A1(_12941_),
    .A2(_12949_),
    .B1(_13107_),
    .B2(_13109_),
    .Y(_13110_));
 sky130_fd_sc_hd__o221ai_4 _23005_ (.A1(_12940_),
    .A2(_12948_),
    .B1(_13101_),
    .B2(net146),
    .C1(_13106_),
    .Y(_13111_));
 sky130_fd_sc_hd__a2bb2oi_2 _23006_ (.A1_N(_12942_),
    .A2_N(_13098_),
    .B1(_13105_),
    .B2(_13106_),
    .Y(_13112_));
 sky130_fd_sc_hd__nand4_4 _23007_ (.A(_12941_),
    .B(_12949_),
    .C(_13107_),
    .D(_13109_),
    .Y(_13113_));
 sky130_fd_sc_hd__a21oi_1 _23008_ (.A1(net138),
    .A2(net134),
    .B1(_13110_),
    .Y(_13114_));
 sky130_fd_sc_hd__o21ai_1 _23009_ (.A1(_10546_),
    .A2(_13112_),
    .B1(_13111_),
    .Y(_13115_));
 sky130_fd_sc_hd__o211ai_4 _23010_ (.A1(_10540_),
    .A2(net135),
    .B1(_13111_),
    .C1(_13113_),
    .Y(_13116_));
 sky130_fd_sc_hd__o21ai_2 _23011_ (.A1(_13110_),
    .A2(_13112_),
    .B1(net133),
    .Y(_13117_));
 sky130_fd_sc_hd__a22o_1 _23012_ (.A1(net138),
    .A2(net134),
    .B1(_13111_),
    .B2(_13113_),
    .X(_13118_));
 sky130_fd_sc_hd__nand4_2 _23013_ (.A(net138),
    .B(net134),
    .C(_13111_),
    .D(_13113_),
    .Y(_13120_));
 sky130_fd_sc_hd__o21ai_1 _23014_ (.A1(_10546_),
    .A2(_12953_),
    .B1(_12952_),
    .Y(_13121_));
 sky130_fd_sc_hd__a22oi_4 _23015_ (.A1(_12947_),
    .A2(_12950_),
    .B1(net133),
    .B2(_12954_),
    .Y(_13122_));
 sky130_fd_sc_hd__nand3_4 _23016_ (.A(_13116_),
    .B(_13117_),
    .C(_13122_),
    .Y(_13123_));
 sky130_fd_sc_hd__nand3_4 _23017_ (.A(_13118_),
    .B(_13120_),
    .C(_13121_),
    .Y(_13124_));
 sky130_fd_sc_hd__o2111ai_4 _23018_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net142),
    .C1(_13123_),
    .D1(_13124_),
    .Y(_13125_));
 sky130_fd_sc_hd__o2bb2ai_4 _23019_ (.A1_N(_13123_),
    .A2_N(_13124_),
    .B1(_11042_),
    .B2(_11742_),
    .Y(_13126_));
 sky130_fd_sc_hd__a21o_1 _23020_ (.A1(_13123_),
    .A2(_13124_),
    .B1(_12099_),
    .X(_13127_));
 sky130_fd_sc_hd__o211ai_1 _23021_ (.A1(_11042_),
    .A2(_11742_),
    .B1(_13123_),
    .C1(_13124_),
    .Y(_13128_));
 sky130_fd_sc_hd__a2bb2oi_4 _23022_ (.A1_N(_12960_),
    .A2_N(_12968_),
    .B1(_13125_),
    .B2(_13126_),
    .Y(_13129_));
 sky130_fd_sc_hd__nand3_1 _23023_ (.A(_13127_),
    .B(_13128_),
    .C(_13096_),
    .Y(_13131_));
 sky130_fd_sc_hd__o211a_1 _23024_ (.A1(_12962_),
    .A2(_13095_),
    .B1(_13125_),
    .C1(_13126_),
    .X(_13132_));
 sky130_fd_sc_hd__o211ai_4 _23025_ (.A1(_12962_),
    .A2(_13095_),
    .B1(_13125_),
    .C1(_13126_),
    .Y(_13133_));
 sky130_fd_sc_hd__o2bb2ai_2 _23026_ (.A1_N(_13092_),
    .A2_N(_13094_),
    .B1(_13129_),
    .B2(_13132_),
    .Y(_13134_));
 sky130_fd_sc_hd__nand3_2 _23027_ (.A(_13092_),
    .B(_13094_),
    .C(_13133_),
    .Y(_13135_));
 sky130_fd_sc_hd__nand4_1 _23028_ (.A(_13092_),
    .B(_13094_),
    .C(_13131_),
    .D(_13133_),
    .Y(_13136_));
 sky130_fd_sc_hd__nand2_2 _23029_ (.A(_12971_),
    .B(_13011_),
    .Y(_13137_));
 sky130_fd_sc_hd__a21oi_2 _23030_ (.A1(_13134_),
    .A2(_13136_),
    .B1(_13137_),
    .Y(_13138_));
 sky130_fd_sc_hd__a21o_2 _23031_ (.A1(_13134_),
    .A2(_13136_),
    .B1(_13137_),
    .X(_13139_));
 sky130_fd_sc_hd__o211a_2 _23032_ (.A1(_13129_),
    .A2(_13135_),
    .B1(_13137_),
    .C1(_13134_),
    .X(_13140_));
 sky130_fd_sc_hd__o211ai_4 _23033_ (.A1(_13129_),
    .A2(_13135_),
    .B1(_13137_),
    .C1(_13134_),
    .Y(_13142_));
 sky130_fd_sc_hd__and2_1 _23034_ (.A(_12998_),
    .B(_13000_),
    .X(_13143_));
 sky130_fd_sc_hd__o21ai_2 _23035_ (.A1(_13000_),
    .A2(_12995_),
    .B1(_12998_),
    .Y(_13144_));
 sky130_fd_sc_hd__o21ai_2 _23036_ (.A1(_12876_),
    .A2(_12894_),
    .B1(_12898_),
    .Y(_13145_));
 sky130_fd_sc_hd__o311a_1 _23037_ (.A1(net246),
    .A2(_05928_),
    .A3(_07074_),
    .B1(net281),
    .C1(_07072_),
    .X(_13146_));
 sky130_fd_sc_hd__nor2_1 _23038_ (.A(_04212_),
    .B(_04218_),
    .Y(_13147_));
 sky130_fd_sc_hd__o22a_1 _23039_ (.A1(_04212_),
    .A2(_04218_),
    .B1(_07079_),
    .B2(_04216_),
    .X(_13148_));
 sky130_fd_sc_hd__a31o_1 _23040_ (.A1(_07072_),
    .A2(net168),
    .A3(net281),
    .B1(_13147_),
    .X(_13149_));
 sky130_fd_sc_hd__nor2_1 _23041_ (.A(_04223_),
    .B(_03737_),
    .Y(_13150_));
 sky130_fd_sc_hd__a211oi_2 _23042_ (.A1(net203),
    .A2(_07500_),
    .B1(_03714_),
    .C1(_07498_),
    .Y(_13151_));
 sky130_fd_sc_hd__a31oi_2 _23043_ (.A1(_07499_),
    .A2(net167),
    .A3(_03704_),
    .B1(_13150_),
    .Y(_13153_));
 sky130_fd_sc_hd__and3_1 _23044_ (.A(_04037_),
    .B(net22),
    .C(net37),
    .X(_13154_));
 sky130_fd_sc_hd__a31oi_1 _23045_ (.A1(_07771_),
    .A2(_02858_),
    .A3(net165),
    .B1(_13154_),
    .Y(_13155_));
 sky130_fd_sc_hd__a31o_1 _23046_ (.A1(_07771_),
    .A2(_02858_),
    .A3(net165),
    .B1(_13154_),
    .X(_13156_));
 sky130_fd_sc_hd__o21ai_4 _23047_ (.A1(_13150_),
    .A2(_13151_),
    .B1(_13156_),
    .Y(_13157_));
 sky130_fd_sc_hd__o221a_2 _23048_ (.A1(_04245_),
    .A2(_02891_),
    .B1(_07772_),
    .B2(_02869_),
    .C1(_13153_),
    .X(_13158_));
 sky130_fd_sc_hd__nand2_2 _23049_ (.A(_13153_),
    .B(_13155_),
    .Y(_13159_));
 sky130_fd_sc_hd__nand2_1 _23050_ (.A(_13157_),
    .B(_13159_),
    .Y(_13160_));
 sky130_fd_sc_hd__a21oi_2 _23051_ (.A1(_13157_),
    .A2(_13159_),
    .B1(_13149_),
    .Y(_13161_));
 sky130_fd_sc_hd__a21o_1 _23052_ (.A1(_13157_),
    .A2(_13159_),
    .B1(_13149_),
    .X(_13162_));
 sky130_fd_sc_hd__o211a_2 _23053_ (.A1(_13146_),
    .A2(_13147_),
    .B1(_13157_),
    .C1(_13159_),
    .X(_13164_));
 sky130_fd_sc_hd__o211ai_1 _23054_ (.A1(_13146_),
    .A2(_13147_),
    .B1(_13157_),
    .C1(_13159_),
    .Y(_13165_));
 sky130_fd_sc_hd__a31oi_2 _23055_ (.A1(_12983_),
    .A2(_12979_),
    .A3(_12981_),
    .B1(_12974_),
    .Y(_13166_));
 sky130_fd_sc_hd__a21oi_2 _23056_ (.A1(_12975_),
    .A2(_12985_),
    .B1(_12986_),
    .Y(_13167_));
 sky130_fd_sc_hd__o21ai_4 _23057_ (.A1(_13161_),
    .A2(_13164_),
    .B1(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__inv_2 _23058_ (.A(_13168_),
    .Y(_13169_));
 sky130_fd_sc_hd__o2bb2ai_2 _23059_ (.A1_N(_13160_),
    .A2_N(_13148_),
    .B1(_12986_),
    .B2(_13166_),
    .Y(_13170_));
 sky130_fd_sc_hd__o211ai_2 _23060_ (.A1(_12986_),
    .A2(_13166_),
    .B1(_13165_),
    .C1(_13162_),
    .Y(_13171_));
 sky130_fd_sc_hd__a21o_1 _23061_ (.A1(_12877_),
    .A2(_12884_),
    .B1(_12885_),
    .X(_13172_));
 sky130_fd_sc_hd__o221a_1 _23062_ (.A1(_12885_),
    .A2(_12888_),
    .B1(_13164_),
    .B2(_13170_),
    .C1(_13168_),
    .X(_13173_));
 sky130_fd_sc_hd__o221ai_4 _23063_ (.A1(_12885_),
    .A2(_12888_),
    .B1(_13164_),
    .B2(_13170_),
    .C1(_13168_),
    .Y(_13175_));
 sky130_fd_sc_hd__a21oi_2 _23064_ (.A1(_13168_),
    .A2(_13171_),
    .B1(_13172_),
    .Y(_13176_));
 sky130_fd_sc_hd__a21o_1 _23065_ (.A1(_13168_),
    .A2(_13171_),
    .B1(_13172_),
    .X(_13177_));
 sky130_fd_sc_hd__o221a_2 _23066_ (.A1(_12876_),
    .A2(_12894_),
    .B1(_13173_),
    .B2(_13176_),
    .C1(_12898_),
    .X(_13178_));
 sky130_fd_sc_hd__o21bai_4 _23067_ (.A1(_13173_),
    .A2(_13176_),
    .B1_N(_13145_),
    .Y(_13179_));
 sky130_fd_sc_hd__nand3_4 _23068_ (.A(_13145_),
    .B(_13175_),
    .C(_13177_),
    .Y(_13180_));
 sky130_fd_sc_hd__inv_2 _23069_ (.A(_13180_),
    .Y(_13181_));
 sky130_fd_sc_hd__a32oi_4 _23070_ (.A1(net182),
    .A2(net179),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net14),
    .Y(_13182_));
 sky130_fd_sc_hd__a32o_1 _23071_ (.A1(net182),
    .A2(net179),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net14),
    .X(_13183_));
 sky130_fd_sc_hd__and3_1 _23072_ (.A(_04124_),
    .B(net16),
    .C(net43),
    .X(_13184_));
 sky130_fd_sc_hd__a31oi_4 _23073_ (.A1(_05933_),
    .A2(net242),
    .A3(net174),
    .B1(_13184_),
    .Y(_13186_));
 sky130_fd_sc_hd__a31o_1 _23074_ (.A1(_05933_),
    .A2(net242),
    .A3(net174),
    .B1(_13184_),
    .X(_13187_));
 sky130_fd_sc_hd__nor2_1 _23075_ (.A(_04146_),
    .B(_05229_),
    .Y(_13188_));
 sky130_fd_sc_hd__a31oi_4 _23076_ (.A1(net178),
    .A2(net177),
    .A3(_05225_),
    .B1(_13188_),
    .Y(_13189_));
 sky130_fd_sc_hd__a31o_1 _23077_ (.A1(net178),
    .A2(net177),
    .A3(_05225_),
    .B1(_13188_),
    .X(_13190_));
 sky130_fd_sc_hd__nor2_2 _23078_ (.A(_13186_),
    .B(_13189_),
    .Y(_13191_));
 sky130_fd_sc_hd__o221a_4 _23079_ (.A1(_04157_),
    .A2(_04989_),
    .B1(_05935_),
    .B2(_04986_),
    .C1(_13189_),
    .X(_13192_));
 sky130_fd_sc_hd__o21ai_4 _23080_ (.A1(_13191_),
    .A2(_13192_),
    .B1(_13182_),
    .Y(_13193_));
 sky130_fd_sc_hd__o21ai_2 _23081_ (.A1(_13186_),
    .A2(_13189_),
    .B1(_13183_),
    .Y(_13194_));
 sky130_fd_sc_hd__a21o_1 _23082_ (.A1(_13186_),
    .A2(_13189_),
    .B1(_13194_),
    .X(_13195_));
 sky130_fd_sc_hd__o21a_1 _23083_ (.A1(_13192_),
    .A2(_13194_),
    .B1(_13193_),
    .X(_13197_));
 sky130_fd_sc_hd__o21ai_1 _23084_ (.A1(_13192_),
    .A2(_13194_),
    .B1(_13193_),
    .Y(_13198_));
 sky130_fd_sc_hd__a21o_2 _23085_ (.A1(_12853_),
    .A2(_12861_),
    .B1(_12858_),
    .X(_13199_));
 sky130_fd_sc_hd__a32o_1 _23086_ (.A1(net202),
    .A2(net173),
    .A3(_04895_),
    .B1(_04897_),
    .B2(net17),
    .X(_13200_));
 sky130_fd_sc_hd__nor2_1 _23087_ (.A(_04179_),
    .B(_04483_),
    .Y(_13201_));
 sky130_fd_sc_hd__a31oi_4 _23088_ (.A1(net198),
    .A2(net172),
    .A3(net279),
    .B1(_13201_),
    .Y(_13202_));
 sky130_fd_sc_hd__or3b_1 _23089_ (.A(net41),
    .B(_04201_),
    .C_N(net40),
    .X(_13203_));
 sky130_fd_sc_hd__o211ai_2 _23090_ (.A1(net174),
    .A2(_06759_),
    .B1(_04267_),
    .C1(net193),
    .Y(_13204_));
 sky130_fd_sc_hd__o311a_1 _23091_ (.A1(_04268_),
    .A2(_06756_),
    .A3(net189),
    .B1(_13203_),
    .C1(_13202_),
    .X(_13205_));
 sky130_fd_sc_hd__o211ai_2 _23092_ (.A1(_04201_),
    .A2(_04270_),
    .B1(_13204_),
    .C1(_13202_),
    .Y(_13206_));
 sky130_fd_sc_hd__a21oi_2 _23093_ (.A1(_13203_),
    .A2(_13204_),
    .B1(_13202_),
    .Y(_13208_));
 sky130_fd_sc_hd__a21o_2 _23094_ (.A1(_13203_),
    .A2(_13204_),
    .B1(_13202_),
    .X(_13209_));
 sky130_fd_sc_hd__nand3_4 _23095_ (.A(_13200_),
    .B(_13206_),
    .C(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__o21bai_4 _23096_ (.A1(_13205_),
    .A2(_13208_),
    .B1_N(_13200_),
    .Y(_13211_));
 sky130_fd_sc_hd__and3_2 _23097_ (.A(_13199_),
    .B(_13210_),
    .C(_13211_),
    .X(_13212_));
 sky130_fd_sc_hd__o211ai_2 _23098_ (.A1(_12858_),
    .A2(_12863_),
    .B1(_13210_),
    .C1(_13211_),
    .Y(_13213_));
 sky130_fd_sc_hd__a21oi_4 _23099_ (.A1(_13210_),
    .A2(_13211_),
    .B1(_13199_),
    .Y(_13214_));
 sky130_fd_sc_hd__a221o_2 _23100_ (.A1(_12853_),
    .A2(_12861_),
    .B1(_13210_),
    .B2(_13211_),
    .C1(_12858_),
    .X(_13215_));
 sky130_fd_sc_hd__o221a_1 _23101_ (.A1(_13194_),
    .A2(_13192_),
    .B1(_13214_),
    .B2(_13212_),
    .C1(_13193_),
    .X(_13216_));
 sky130_fd_sc_hd__o21ai_1 _23102_ (.A1(_13212_),
    .A2(_13214_),
    .B1(_13197_),
    .Y(_13217_));
 sky130_fd_sc_hd__and3_1 _23103_ (.A(_13198_),
    .B(_13213_),
    .C(_13215_),
    .X(_13219_));
 sky130_fd_sc_hd__a211o_1 _23104_ (.A1(_13193_),
    .A2(_13195_),
    .B1(_13212_),
    .C1(_13214_),
    .X(_13220_));
 sky130_fd_sc_hd__nand2_2 _23105_ (.A(_13215_),
    .B(_13197_),
    .Y(_13221_));
 sky130_fd_sc_hd__and3_1 _23106_ (.A(_13215_),
    .B(_13197_),
    .C(_13213_),
    .X(_13222_));
 sky130_fd_sc_hd__o2bb2a_1 _23107_ (.A1_N(_13193_),
    .A2_N(_13195_),
    .B1(_13212_),
    .B2(_13214_),
    .X(_13223_));
 sky130_fd_sc_hd__a22o_1 _23108_ (.A1(_13193_),
    .A2(_13195_),
    .B1(_13213_),
    .B2(_13215_),
    .X(_13224_));
 sky130_fd_sc_hd__o21ai_2 _23109_ (.A1(_13212_),
    .A2(_13221_),
    .B1(_13224_),
    .Y(_13225_));
 sky130_fd_sc_hd__nand4_2 _23110_ (.A(_13179_),
    .B(_13180_),
    .C(_13217_),
    .D(_13220_),
    .Y(_13226_));
 sky130_fd_sc_hd__o2bb2ai_1 _23111_ (.A1_N(_13179_),
    .A2_N(_13180_),
    .B1(_13216_),
    .B2(_13219_),
    .Y(_13227_));
 sky130_fd_sc_hd__o2bb2ai_2 _23112_ (.A1_N(_13179_),
    .A2_N(_13180_),
    .B1(_13222_),
    .B2(_13223_),
    .Y(_13228_));
 sky130_fd_sc_hd__o211a_1 _23113_ (.A1(_13212_),
    .A2(_13221_),
    .B1(_13224_),
    .C1(_13179_),
    .X(_13230_));
 sky130_fd_sc_hd__o2111ai_4 _23114_ (.A1(_13212_),
    .A2(_13221_),
    .B1(_13224_),
    .C1(_13180_),
    .D1(_13179_),
    .Y(_13231_));
 sky130_fd_sc_hd__inv_2 _23115_ (.A(_13231_),
    .Y(_13232_));
 sky130_fd_sc_hd__o211ai_4 _23116_ (.A1(_12995_),
    .A2(_13143_),
    .B1(_13226_),
    .C1(_13227_),
    .Y(_13233_));
 sky130_fd_sc_hd__nand2_1 _23117_ (.A(_13228_),
    .B(_13144_),
    .Y(_13234_));
 sky130_fd_sc_hd__nand3_2 _23118_ (.A(_13228_),
    .B(_13231_),
    .C(_13144_),
    .Y(_13235_));
 sky130_fd_sc_hd__o21ai_2 _23119_ (.A1(_12874_),
    .A2(_12907_),
    .B1(_12906_),
    .Y(_13236_));
 sky130_fd_sc_hd__a22oi_2 _23120_ (.A1(_12908_),
    .A2(_12910_),
    .B1(_13233_),
    .B2(_13235_),
    .Y(_13237_));
 sky130_fd_sc_hd__a22o_2 _23121_ (.A1(_12908_),
    .A2(_12910_),
    .B1(_13233_),
    .B2(_13235_),
    .X(_13238_));
 sky130_fd_sc_hd__o211a_1 _23122_ (.A1(_12905_),
    .A2(_12913_),
    .B1(_13233_),
    .C1(_13235_),
    .X(_13239_));
 sky130_fd_sc_hd__o211ai_4 _23123_ (.A1(_12905_),
    .A2(_12913_),
    .B1(_13233_),
    .C1(_13235_),
    .Y(_13241_));
 sky130_fd_sc_hd__o211ai_2 _23124_ (.A1(_13138_),
    .A2(_13140_),
    .B1(_13238_),
    .C1(_13241_),
    .Y(_13242_));
 sky130_fd_sc_hd__o211ai_2 _23125_ (.A1(_13237_),
    .A2(_13239_),
    .B1(_13139_),
    .C1(_13142_),
    .Y(_13243_));
 sky130_fd_sc_hd__o22a_1 _23126_ (.A1(_13138_),
    .A2(_13140_),
    .B1(_13237_),
    .B2(_13239_),
    .X(_13244_));
 sky130_fd_sc_hd__o22ai_2 _23127_ (.A1(_13138_),
    .A2(_13140_),
    .B1(_13237_),
    .B2(_13239_),
    .Y(_13245_));
 sky130_fd_sc_hd__and4_1 _23128_ (.A(_13139_),
    .B(_13142_),
    .C(_13238_),
    .D(_13241_),
    .X(_13246_));
 sky130_fd_sc_hd__nand4_2 _23129_ (.A(_13139_),
    .B(_13142_),
    .C(_13238_),
    .D(_13241_),
    .Y(_13247_));
 sky130_fd_sc_hd__and3_1 _23130_ (.A(_12924_),
    .B(_12928_),
    .C(_13016_),
    .X(_13248_));
 sky130_fd_sc_hd__o211ai_2 _23131_ (.A1(_12917_),
    .A2(_12575_),
    .B1(_13016_),
    .C1(_12928_),
    .Y(_13249_));
 sky130_fd_sc_hd__nand3_1 _23132_ (.A(_12921_),
    .B(_12923_),
    .C(_13014_),
    .Y(_13250_));
 sky130_fd_sc_hd__nand4_4 _23133_ (.A(_13014_),
    .B(_13245_),
    .C(_13247_),
    .D(_13249_),
    .Y(_13252_));
 sky130_fd_sc_hd__nand4_4 _23134_ (.A(_13016_),
    .B(_13242_),
    .C(_13243_),
    .D(_13250_),
    .Y(_13253_));
 sky130_fd_sc_hd__a21oi_1 _23135_ (.A1(_12763_),
    .A2(_12767_),
    .B1(_12764_),
    .Y(_13254_));
 sky130_fd_sc_hd__a21o_1 _23136_ (.A1(_12741_),
    .A2(_12744_),
    .B1(_12740_),
    .X(_13255_));
 sky130_fd_sc_hd__o211ai_2 _23137_ (.A1(_04787_),
    .A2(net208),
    .B1(_05762_),
    .C1(net209),
    .Y(_13256_));
 sky130_fd_sc_hd__or3b_2 _23138_ (.A(_04113_),
    .B(net48),
    .C_N(net47),
    .X(_13257_));
 sky130_fd_sc_hd__o211ai_2 _23139_ (.A1(net233),
    .A2(_04787_),
    .B1(net274),
    .C1(net213),
    .Y(_13258_));
 sky130_fd_sc_hd__or3b_2 _23140_ (.A(_04091_),
    .B(net49),
    .C_N(net48),
    .X(_13259_));
 sky130_fd_sc_hd__a22oi_2 _23141_ (.A1(_13256_),
    .A2(_13257_),
    .B1(_13258_),
    .B2(_13259_),
    .Y(_13260_));
 sky130_fd_sc_hd__a22o_1 _23142_ (.A1(_13256_),
    .A2(_13257_),
    .B1(_13258_),
    .B2(_13259_),
    .X(_13261_));
 sky130_fd_sc_hd__nand4_2 _23143_ (.A(_13256_),
    .B(_13257_),
    .C(_13258_),
    .D(_13259_),
    .Y(_13263_));
 sky130_fd_sc_hd__a32o_1 _23144_ (.A1(net217),
    .A2(net186),
    .A3(net273),
    .B1(_06326_),
    .B2(net10),
    .X(_13264_));
 sky130_fd_sc_hd__a21oi_1 _23145_ (.A1(_13261_),
    .A2(_13263_),
    .B1(_13264_),
    .Y(_13265_));
 sky130_fd_sc_hd__a21o_1 _23146_ (.A1(_13261_),
    .A2(_13263_),
    .B1(_13264_),
    .X(_13266_));
 sky130_fd_sc_hd__and3_1 _23147_ (.A(_13261_),
    .B(_13263_),
    .C(_13264_),
    .X(_13267_));
 sky130_fd_sc_hd__nand3_1 _23148_ (.A(_13261_),
    .B(_13263_),
    .C(_13264_),
    .Y(_13268_));
 sky130_fd_sc_hd__o2bb2ai_2 _23149_ (.A1_N(_12843_),
    .A2_N(_12847_),
    .B1(_13265_),
    .B2(_13267_),
    .Y(_13269_));
 sky130_fd_sc_hd__nand3_4 _23150_ (.A(_13266_),
    .B(_13268_),
    .C(_12849_),
    .Y(_13270_));
 sky130_fd_sc_hd__a21oi_1 _23151_ (.A1(_13269_),
    .A2(_13270_),
    .B1(_13255_),
    .Y(_13271_));
 sky130_fd_sc_hd__a21o_1 _23152_ (.A1(_13269_),
    .A2(_13270_),
    .B1(_13255_),
    .X(_13272_));
 sky130_fd_sc_hd__o211a_2 _23153_ (.A1(_12740_),
    .A2(_12748_),
    .B1(_13269_),
    .C1(_13270_),
    .X(_13274_));
 sky130_fd_sc_hd__o211ai_4 _23154_ (.A1(_12740_),
    .A2(_12748_),
    .B1(_13269_),
    .C1(_13270_),
    .Y(_13275_));
 sky130_fd_sc_hd__o22ai_4 _23155_ (.A1(_12865_),
    .A2(_12863_),
    .B1(_12851_),
    .B2(_12868_),
    .Y(_13276_));
 sky130_fd_sc_hd__o21bai_4 _23156_ (.A1(_13271_),
    .A2(_13274_),
    .B1_N(_13276_),
    .Y(_13277_));
 sky130_fd_sc_hd__nand2_1 _23157_ (.A(_13272_),
    .B(_13276_),
    .Y(_13278_));
 sky130_fd_sc_hd__nand3_1 _23158_ (.A(_13272_),
    .B(_13275_),
    .C(_13276_),
    .Y(_13279_));
 sky130_fd_sc_hd__and3_1 _23159_ (.A(_12612_),
    .B(_12616_),
    .C(_12755_),
    .X(_13280_));
 sky130_fd_sc_hd__o31a_2 _23160_ (.A1(_12611_),
    .A2(_12614_),
    .A3(_12754_),
    .B1(_12753_),
    .X(_13281_));
 sky130_fd_sc_hd__o211ai_4 _23161_ (.A1(_13274_),
    .A2(_13278_),
    .B1(_13281_),
    .C1(_13277_),
    .Y(_13282_));
 sky130_fd_sc_hd__o2bb2ai_2 _23162_ (.A1_N(_13277_),
    .A2_N(_13279_),
    .B1(_13280_),
    .B2(_12752_),
    .Y(_13283_));
 sky130_fd_sc_hd__o211a_1 _23163_ (.A1(_12764_),
    .A2(_12770_),
    .B1(_13282_),
    .C1(_13283_),
    .X(_13285_));
 sky130_fd_sc_hd__o211ai_4 _23164_ (.A1(_12764_),
    .A2(_12770_),
    .B1(_13282_),
    .C1(_13283_),
    .Y(_13286_));
 sky130_fd_sc_hd__a32oi_4 _23165_ (.A1(_00625_),
    .A2(net250),
    .A3(net238),
    .B1(_08006_),
    .B2(net5),
    .Y(_13287_));
 sky130_fd_sc_hd__a32oi_4 _23166_ (.A1(net229),
    .A2(net227),
    .A3(net269),
    .B1(_07225_),
    .B2(net8),
    .Y(_13288_));
 sky130_fd_sc_hd__nand4_2 _23167_ (.A(_04190_),
    .B(net225),
    .C(net51),
    .D(_04409_),
    .Y(_13289_));
 sky130_fd_sc_hd__or3_1 _23168_ (.A(net51),
    .B(_04190_),
    .C(_04069_),
    .X(_13290_));
 sky130_fd_sc_hd__a21oi_1 _23169_ (.A1(_13289_),
    .A2(_13290_),
    .B1(_13288_),
    .Y(_13291_));
 sky130_fd_sc_hd__a21o_1 _23170_ (.A1(_13289_),
    .A2(_13290_),
    .B1(_13288_),
    .X(_13292_));
 sky130_fd_sc_hd__and3_1 _23171_ (.A(_13288_),
    .B(_13289_),
    .C(_13290_),
    .X(_13293_));
 sky130_fd_sc_hd__o211ai_2 _23172_ (.A1(_04069_),
    .A2(_06866_),
    .B1(_13289_),
    .C1(_13288_),
    .Y(_13294_));
 sky130_fd_sc_hd__a32o_1 _23173_ (.A1(_03952_),
    .A2(net233),
    .A3(net239),
    .B1(_07308_),
    .B2(net7),
    .X(_13296_));
 sky130_fd_sc_hd__o21bai_2 _23174_ (.A1(_13291_),
    .A2(_13293_),
    .B1_N(_13296_),
    .Y(_13297_));
 sky130_fd_sc_hd__nand3_4 _23175_ (.A(_13292_),
    .B(_13294_),
    .C(_13296_),
    .Y(_13298_));
 sky130_fd_sc_hd__a21oi_1 _23176_ (.A1(_12786_),
    .A2(_12789_),
    .B1(_12784_),
    .Y(_13299_));
 sky130_fd_sc_hd__o21ai_1 _23177_ (.A1(_12785_),
    .A2(_12788_),
    .B1(_12783_),
    .Y(_13300_));
 sky130_fd_sc_hd__o2bb2ai_2 _23178_ (.A1_N(_13297_),
    .A2_N(_13298_),
    .B1(_13299_),
    .B2(_12792_),
    .Y(_13301_));
 sky130_fd_sc_hd__nand4_4 _23179_ (.A(_12793_),
    .B(_13297_),
    .C(_13298_),
    .D(_13300_),
    .Y(_13302_));
 sky130_fd_sc_hd__a32o_1 _23180_ (.A1(_02421_),
    .A2(net248),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net6),
    .X(_13303_));
 sky130_fd_sc_hd__a21o_1 _23181_ (.A1(_13301_),
    .A2(_13302_),
    .B1(_13303_),
    .X(_13304_));
 sky130_fd_sc_hd__nand3_4 _23182_ (.A(_13301_),
    .B(_13302_),
    .C(_13303_),
    .Y(_13305_));
 sky130_fd_sc_hd__a21bo_1 _23183_ (.A1(_12781_),
    .A2(_12798_),
    .B1_N(_12799_),
    .X(_13307_));
 sky130_fd_sc_hd__and3_1 _23184_ (.A(_13304_),
    .B(_13307_),
    .C(_13305_),
    .X(_13308_));
 sky130_fd_sc_hd__a21oi_4 _23185_ (.A1(_13304_),
    .A2(_13305_),
    .B1(_13307_),
    .Y(_13309_));
 sky130_fd_sc_hd__o21ai_2 _23186_ (.A1(_13308_),
    .A2(_13309_),
    .B1(_13287_),
    .Y(_13310_));
 sky130_fd_sc_hd__a31o_1 _23187_ (.A1(_13304_),
    .A2(_13307_),
    .A3(_13305_),
    .B1(_13287_),
    .X(_13311_));
 sky130_fd_sc_hd__o21ai_2 _23188_ (.A1(_13309_),
    .A2(_13311_),
    .B1(_13310_),
    .Y(_13312_));
 sky130_fd_sc_hd__a21boi_1 _23189_ (.A1(_13282_),
    .A2(_13283_),
    .B1_N(_13254_),
    .Y(_13313_));
 sky130_fd_sc_hd__a21bo_1 _23190_ (.A1(_13282_),
    .A2(_13283_),
    .B1_N(_13254_),
    .X(_13314_));
 sky130_fd_sc_hd__o2111ai_4 _23191_ (.A1(_13311_),
    .A2(_13309_),
    .B1(_13286_),
    .C1(_13310_),
    .D1(_13314_),
    .Y(_13315_));
 sky130_fd_sc_hd__o21ai_1 _23192_ (.A1(_13285_),
    .A2(_13313_),
    .B1(_13312_),
    .Y(_13316_));
 sky130_fd_sc_hd__nand3_1 _23193_ (.A(_13286_),
    .B(_13312_),
    .C(_13314_),
    .Y(_13318_));
 sky130_fd_sc_hd__o21bai_1 _23194_ (.A1(_13285_),
    .A2(_13313_),
    .B1_N(_13312_),
    .Y(_13319_));
 sky130_fd_sc_hd__nand3_2 _23195_ (.A(_12927_),
    .B(_13318_),
    .C(_13319_),
    .Y(_13320_));
 sky130_fd_sc_hd__o211ai_4 _23196_ (.A1(_12916_),
    .A2(_12920_),
    .B1(_13315_),
    .C1(_13316_),
    .Y(_13321_));
 sky130_fd_sc_hd__inv_2 _23197_ (.A(_13321_),
    .Y(_13322_));
 sky130_fd_sc_hd__o21a_1 _23198_ (.A1(_12808_),
    .A2(_12810_),
    .B1(_12775_),
    .X(_13323_));
 sky130_fd_sc_hd__a31o_1 _23199_ (.A1(_12777_),
    .A2(_12809_),
    .A3(_12811_),
    .B1(_12774_),
    .X(_13324_));
 sky130_fd_sc_hd__a21oi_2 _23200_ (.A1(_13320_),
    .A2(_13321_),
    .B1(_13324_),
    .Y(_13325_));
 sky130_fd_sc_hd__o2bb2ai_1 _23201_ (.A1_N(_13320_),
    .A2_N(_13321_),
    .B1(_13323_),
    .B2(_12776_),
    .Y(_13326_));
 sky130_fd_sc_hd__o211a_2 _23202_ (.A1(_12774_),
    .A2(_12817_),
    .B1(_13320_),
    .C1(_13321_),
    .X(_13327_));
 sky130_fd_sc_hd__o211ai_2 _23203_ (.A1(_12774_),
    .A2(_12817_),
    .B1(_13320_),
    .C1(_13321_),
    .Y(_13329_));
 sky130_fd_sc_hd__nor2_1 _23204_ (.A(_13325_),
    .B(_13327_),
    .Y(_13330_));
 sky130_fd_sc_hd__nand3_2 _23205_ (.A(_13253_),
    .B(_13326_),
    .C(_13329_),
    .Y(_13331_));
 sky130_fd_sc_hd__nand2_1 _23206_ (.A(_13252_),
    .B(_13253_),
    .Y(_13332_));
 sky130_fd_sc_hd__nand4_1 _23207_ (.A(_13252_),
    .B(_13253_),
    .C(_13326_),
    .D(_13329_),
    .Y(_13333_));
 sky130_fd_sc_hd__o2bb2ai_1 _23208_ (.A1_N(_13252_),
    .A2_N(_13253_),
    .B1(_13325_),
    .B2(_13327_),
    .Y(_13334_));
 sky130_fd_sc_hd__o211ai_4 _23209_ (.A1(_13325_),
    .A2(_13327_),
    .B1(_13252_),
    .C1(_13253_),
    .Y(_13335_));
 sky130_fd_sc_hd__nand2_1 _23210_ (.A(_13330_),
    .B(_13332_),
    .Y(_13336_));
 sky130_fd_sc_hd__and3_1 _23211_ (.A(_13334_),
    .B(_13060_),
    .C(_13333_),
    .X(_13337_));
 sky130_fd_sc_hd__nand3_2 _23212_ (.A(_13334_),
    .B(_13060_),
    .C(_13333_),
    .Y(_13338_));
 sky130_fd_sc_hd__nand3_2 _23213_ (.A(_13061_),
    .B(_13335_),
    .C(_13336_),
    .Y(_13340_));
 sky130_fd_sc_hd__and3_1 _23214_ (.A(_12645_),
    .B(_12686_),
    .C(_12819_),
    .X(_13341_));
 sky130_fd_sc_hd__a21oi_1 _23215_ (.A1(_12645_),
    .A2(_12686_),
    .B1(_12821_),
    .Y(_13342_));
 sky130_fd_sc_hd__a31o_1 _23216_ (.A1(_12645_),
    .A2(_12686_),
    .A3(_12819_),
    .B1(_12821_),
    .X(_13343_));
 sky130_fd_sc_hd__o2bb2ai_1 _23217_ (.A1_N(_13338_),
    .A2_N(_13340_),
    .B1(_13342_),
    .B2(_12820_),
    .Y(_13344_));
 sky130_fd_sc_hd__o2111ai_1 _23218_ (.A1(_12821_),
    .A2(_12825_),
    .B1(_13338_),
    .C1(_13340_),
    .D1(_12819_),
    .Y(_13345_));
 sky130_fd_sc_hd__o2bb2ai_1 _23219_ (.A1_N(_13338_),
    .A2_N(_13340_),
    .B1(_13341_),
    .B2(_12821_),
    .Y(_13346_));
 sky130_fd_sc_hd__a31oi_4 _23220_ (.A1(_13061_),
    .A2(_13335_),
    .A3(_13336_),
    .B1(_13343_),
    .Y(_13347_));
 sky130_fd_sc_hd__o211ai_1 _23221_ (.A1(_12820_),
    .A2(_13342_),
    .B1(_13340_),
    .C1(_13338_),
    .Y(_13348_));
 sky130_fd_sc_hd__nand3_2 _23222_ (.A(_13344_),
    .B(_13345_),
    .C(_13058_),
    .Y(_13349_));
 sky130_fd_sc_hd__and3_2 _23223_ (.A(_13059_),
    .B(_13346_),
    .C(_13348_),
    .X(_13351_));
 sky130_fd_sc_hd__nand3_2 _23224_ (.A(_13059_),
    .B(_13346_),
    .C(_13348_),
    .Y(_13352_));
 sky130_fd_sc_hd__nor2_1 _23225_ (.A(_12807_),
    .B(_12806_),
    .Y(_13353_));
 sky130_fd_sc_hd__and2_1 _23226_ (.A(_12803_),
    .B(_12807_),
    .X(_13354_));
 sky130_fd_sc_hd__o21a_1 _23227_ (.A1(_12806_),
    .A2(_13354_),
    .B1(_13349_),
    .X(_13355_));
 sky130_fd_sc_hd__o21ai_2 _23228_ (.A1(_12806_),
    .A2(_13354_),
    .B1(_13349_),
    .Y(_13356_));
 sky130_fd_sc_hd__o2bb2ai_1 _23229_ (.A1_N(_13349_),
    .A2_N(_13352_),
    .B1(_13353_),
    .B2(_12804_),
    .Y(_13357_));
 sky130_fd_sc_hd__o2bb2ai_1 _23230_ (.A1_N(_13349_),
    .A2_N(_13352_),
    .B1(_13354_),
    .B2(_12806_),
    .Y(_13358_));
 sky130_fd_sc_hd__o211ai_2 _23231_ (.A1(_12804_),
    .A2(_13353_),
    .B1(_13352_),
    .C1(_13349_),
    .Y(_13359_));
 sky130_fd_sc_hd__nand2_1 _23232_ (.A(_13358_),
    .B(_13359_),
    .Y(_13360_));
 sky130_fd_sc_hd__and4_1 _23233_ (.A(_13045_),
    .B(_13049_),
    .C(_13358_),
    .D(_13359_),
    .X(_13362_));
 sky130_fd_sc_hd__nand4_2 _23234_ (.A(_13045_),
    .B(_13049_),
    .C(_13358_),
    .D(_13359_),
    .Y(_13363_));
 sky130_fd_sc_hd__o211ai_2 _23235_ (.A1(_13351_),
    .A2(_13356_),
    .B1(_13357_),
    .C1(_13057_),
    .Y(_13364_));
 sky130_fd_sc_hd__nand2_1 _23236_ (.A(_13363_),
    .B(_13364_),
    .Y(_13365_));
 sky130_fd_sc_hd__a21boi_1 _23237_ (.A1(_13052_),
    .A2(_13056_),
    .B1_N(_13051_),
    .Y(_13366_));
 sky130_fd_sc_hd__xnor2_1 _23238_ (.A(_13365_),
    .B(_13366_),
    .Y(net102));
 sky130_fd_sc_hd__o21bai_2 _23239_ (.A1(_13287_),
    .A2(_13309_),
    .B1_N(_13308_),
    .Y(_13367_));
 sky130_fd_sc_hd__inv_2 _23240_ (.A(_13367_),
    .Y(_13368_));
 sky130_fd_sc_hd__a21oi_2 _23241_ (.A1(_13320_),
    .A2(_13324_),
    .B1(_13322_),
    .Y(_13369_));
 sky130_fd_sc_hd__o41a_1 _23242_ (.A1(_13013_),
    .A2(_13244_),
    .A3(_13246_),
    .A4(_13248_),
    .B1(_13331_),
    .X(_13370_));
 sky130_fd_sc_hd__o41ai_4 _23243_ (.A1(_13013_),
    .A2(_13244_),
    .A3(_13246_),
    .A4(_13248_),
    .B1(_13331_),
    .Y(_13372_));
 sky130_fd_sc_hd__nand3_1 _23244_ (.A(_13139_),
    .B(_13238_),
    .C(_13241_),
    .Y(_13373_));
 sky130_fd_sc_hd__a31o_1 _23245_ (.A1(_13139_),
    .A2(_13238_),
    .A3(_13241_),
    .B1(_13140_),
    .X(_13374_));
 sky130_fd_sc_hd__a31oi_2 _23246_ (.A1(_13139_),
    .A2(_13238_),
    .A3(_13241_),
    .B1(_13140_),
    .Y(_13375_));
 sky130_fd_sc_hd__a41o_1 _23247_ (.A1(net307),
    .A2(net293),
    .A3(net288),
    .A4(_00635_),
    .B1(_08658_),
    .X(_13376_));
 sky130_fd_sc_hd__o22ai_4 _23248_ (.A1(_04015_),
    .A2(_08660_),
    .B1(_00614_),
    .B2(_13376_),
    .Y(_13377_));
 sky130_fd_sc_hd__o2111a_1 _23249_ (.A1(net169),
    .A2(net268),
    .B1(net33),
    .C1(_13377_),
    .D1(net319),
    .X(_13378_));
 sky130_fd_sc_hd__o2111ai_4 _23250_ (.A1(net169),
    .A2(net268),
    .B1(net33),
    .C1(_13377_),
    .D1(net319),
    .Y(_13379_));
 sky130_fd_sc_hd__a31oi_4 _23251_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_13377_),
    .Y(_13380_));
 sky130_fd_sc_hd__a31o_1 _23252_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_13377_),
    .X(_13381_));
 sky130_fd_sc_hd__a21oi_2 _23253_ (.A1(_13379_),
    .A2(_13381_),
    .B1(_09300_),
    .Y(_00001_));
 sky130_fd_sc_hd__o21ai_1 _23254_ (.A1(_13378_),
    .A2(_13380_),
    .B1(net146),
    .Y(_00002_));
 sky130_fd_sc_hd__o22ai_2 _23255_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_13378_),
    .B2(_13380_),
    .Y(_00003_));
 sky130_fd_sc_hd__o2111ai_4 _23256_ (.A1(_04495_),
    .A2(net150),
    .B1(_08882_),
    .C1(_13379_),
    .D1(_13381_),
    .Y(_00004_));
 sky130_fd_sc_hd__a21oi_2 _23257_ (.A1(net156),
    .A2(_13100_),
    .B1(_09300_),
    .Y(_00005_));
 sky130_fd_sc_hd__nand2_1 _23258_ (.A(_13104_),
    .B(net146),
    .Y(_00006_));
 sky130_fd_sc_hd__o21ai_1 _23259_ (.A1(net146),
    .A2(_13101_),
    .B1(_13104_),
    .Y(_00007_));
 sky130_fd_sc_hd__o211a_1 _23260_ (.A1(_13101_),
    .A2(_00005_),
    .B1(_00004_),
    .C1(_00003_),
    .X(_00008_));
 sky130_fd_sc_hd__o211ai_4 _23261_ (.A1(_13101_),
    .A2(_00005_),
    .B1(_00004_),
    .C1(_00003_),
    .Y(_00009_));
 sky130_fd_sc_hd__o211ai_4 _23262_ (.A1(net146),
    .A2(_13380_),
    .B1(_00006_),
    .C1(_13102_),
    .Y(_00010_));
 sky130_fd_sc_hd__o211ai_1 _23263_ (.A1(net146),
    .A2(_13380_),
    .B1(_00007_),
    .C1(_00002_),
    .Y(_00012_));
 sky130_fd_sc_hd__o21ai_1 _23264_ (.A1(_00001_),
    .A2(_00010_),
    .B1(_00009_),
    .Y(_00013_));
 sky130_fd_sc_hd__a2bb2oi_1 _23265_ (.A1_N(_10540_),
    .A2_N(net135),
    .B1(_00009_),
    .B2(_00012_),
    .Y(_00014_));
 sky130_fd_sc_hd__o21ai_1 _23266_ (.A1(_10540_),
    .A2(net135),
    .B1(_00013_),
    .Y(_00015_));
 sky130_fd_sc_hd__o2111a_4 _23267_ (.A1(_00010_),
    .A2(_00001_),
    .B1(net134),
    .C1(net138),
    .D1(_00009_),
    .X(_00016_));
 sky130_fd_sc_hd__o2111ai_1 _23268_ (.A1(_00010_),
    .A2(_00001_),
    .B1(net134),
    .C1(net138),
    .D1(_00009_),
    .Y(_00017_));
 sky130_fd_sc_hd__o22ai_4 _23269_ (.A1(_13112_),
    .A2(_13114_),
    .B1(_00014_),
    .B2(_00016_),
    .Y(_00018_));
 sky130_fd_sc_hd__nand2_2 _23270_ (.A(_00015_),
    .B(_13115_),
    .Y(_00019_));
 sky130_fd_sc_hd__nand3_1 _23271_ (.A(_00015_),
    .B(_00017_),
    .C(_13115_),
    .Y(_00020_));
 sky130_fd_sc_hd__a21oi_1 _23272_ (.A1(_00018_),
    .A2(_00020_),
    .B1(_12099_),
    .Y(_00021_));
 sky130_fd_sc_hd__a21o_1 _23273_ (.A1(_00018_),
    .A2(_00020_),
    .B1(_12099_),
    .X(_00023_));
 sky130_fd_sc_hd__o311a_1 _23274_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_00018_),
    .C1(_00020_),
    .X(_00024_));
 sky130_fd_sc_hd__o221ai_4 _23275_ (.A1(_11042_),
    .A2(_11742_),
    .B1(_00016_),
    .B2(_00019_),
    .C1(_00018_),
    .Y(_00025_));
 sky130_fd_sc_hd__a32oi_4 _23276_ (.A1(_13116_),
    .A2(_13117_),
    .A3(_13122_),
    .B1(_13124_),
    .B2(net132),
    .Y(_00026_));
 sky130_fd_sc_hd__o21bai_4 _23277_ (.A1(_00021_),
    .A2(_00024_),
    .B1_N(_00026_),
    .Y(_00027_));
 sky130_fd_sc_hd__and3_1 _23278_ (.A(_00023_),
    .B(_00025_),
    .C(_00026_),
    .X(_00028_));
 sky130_fd_sc_hd__nand3_2 _23279_ (.A(_00023_),
    .B(_00025_),
    .C(_00026_),
    .Y(_00029_));
 sky130_fd_sc_hd__a21oi_2 _23280_ (.A1(net150),
    .A2(_08668_),
    .B1(_01304_),
    .Y(_00030_));
 sky130_fd_sc_hd__nor2_2 _23281_ (.A(net319),
    .B(_01326_),
    .Y(_00031_));
 sky130_fd_sc_hd__or3b_1 _23282_ (.A(net37),
    .B(net319),
    .C_N(net36),
    .X(_00032_));
 sky130_fd_sc_hd__o22a_1 _23283_ (.A1(net319),
    .A2(_01326_),
    .B1(_01304_),
    .B2(_08669_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _23284_ (.A1(net25),
    .A2(_01315_),
    .B1(_08670_),
    .B2(_01293_),
    .X(_00035_));
 sky130_fd_sc_hd__a22oi_4 _23285_ (.A1(net25),
    .A2(_12352_),
    .B1(net159),
    .B2(_12330_),
    .Y(_00036_));
 sky130_fd_sc_hd__o311a_4 _23286_ (.A1(net25),
    .A2(_12341_),
    .A3(net154),
    .B1(_13070_),
    .C1(_13073_),
    .X(_00037_));
 sky130_fd_sc_hd__a221o_2 _23287_ (.A1(net25),
    .A2(_12352_),
    .B1(net159),
    .B2(_12330_),
    .C1(_13074_),
    .X(_00038_));
 sky130_fd_sc_hd__o2bb2ai_4 _23288_ (.A1_N(_13073_),
    .A2_N(_00036_),
    .B1(_00031_),
    .B2(_00030_),
    .Y(_00039_));
 sky130_fd_sc_hd__nand4b_4 _23289_ (.A_N(_00030_),
    .B(_00032_),
    .C(_00036_),
    .D(_13073_),
    .Y(_00040_));
 sky130_fd_sc_hd__o211ai_4 _23290_ (.A1(_12451_),
    .A2(_12454_),
    .B1(_00039_),
    .C1(_00040_),
    .Y(_00041_));
 sky130_fd_sc_hd__a21o_1 _23291_ (.A1(_00039_),
    .A2(_00040_),
    .B1(_13066_),
    .X(_00042_));
 sky130_fd_sc_hd__o2bb2ai_2 _23292_ (.A1_N(_00041_),
    .A2_N(_00042_),
    .B1(net134),
    .B2(_11735_),
    .Y(_00043_));
 sky130_fd_sc_hd__o2111ai_4 _23293_ (.A1(_11527_),
    .A2(_11732_),
    .B1(net135),
    .C1(_00041_),
    .D1(_00042_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand2_1 _23294_ (.A(_00043_),
    .B(_00045_),
    .Y(_00046_));
 sky130_fd_sc_hd__o2111a_1 _23295_ (.A1(_12451_),
    .A2(_12454_),
    .B1(_13080_),
    .C1(_13082_),
    .D1(_00046_),
    .X(_00047_));
 sky130_fd_sc_hd__a21o_1 _23296_ (.A1(_00043_),
    .A2(_00045_),
    .B1(_13087_),
    .X(_00048_));
 sky130_fd_sc_hd__o311a_1 _23297_ (.A1(_13065_),
    .A2(_13079_),
    .A3(_13081_),
    .B1(_00043_),
    .C1(_00045_),
    .X(_00049_));
 sky130_fd_sc_hd__a31o_1 _23298_ (.A1(_13066_),
    .A2(_13080_),
    .A3(_13082_),
    .B1(_00046_),
    .X(_00050_));
 sky130_fd_sc_hd__nand2_1 _23299_ (.A(_00048_),
    .B(_00050_),
    .Y(_00051_));
 sky130_fd_sc_hd__o2bb2ai_1 _23300_ (.A1_N(_00027_),
    .A2_N(_00029_),
    .B1(_00047_),
    .B2(_00049_),
    .Y(_00052_));
 sky130_fd_sc_hd__nand4_2 _23301_ (.A(_00027_),
    .B(_00029_),
    .C(_00048_),
    .D(_00050_),
    .Y(_00053_));
 sky130_fd_sc_hd__a21o_1 _23302_ (.A1(_00027_),
    .A2(_00029_),
    .B1(_00051_),
    .X(_00054_));
 sky130_fd_sc_hd__o21a_1 _23303_ (.A1(_00047_),
    .A2(_00049_),
    .B1(_00027_),
    .X(_00056_));
 sky130_fd_sc_hd__o211ai_2 _23304_ (.A1(_00047_),
    .A2(_00049_),
    .B1(_00027_),
    .C1(_00029_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand2_2 _23305_ (.A(_00054_),
    .B(_00057_),
    .Y(_00058_));
 sky130_fd_sc_hd__a31o_1 _23306_ (.A1(_13092_),
    .A2(_13094_),
    .A3(_13133_),
    .B1(_13129_),
    .X(_00059_));
 sky130_fd_sc_hd__a31oi_4 _23307_ (.A1(_13092_),
    .A2(_13094_),
    .A3(_13133_),
    .B1(_13129_),
    .Y(_00060_));
 sky130_fd_sc_hd__nand3_2 _23308_ (.A(_00054_),
    .B(_00057_),
    .C(_00059_),
    .Y(_00061_));
 sky130_fd_sc_hd__nand3_4 _23309_ (.A(_00052_),
    .B(_00053_),
    .C(_00060_),
    .Y(_00062_));
 sky130_fd_sc_hd__nand2_1 _23310_ (.A(_00061_),
    .B(_00062_),
    .Y(_00063_));
 sky130_fd_sc_hd__a32o_2 _23311_ (.A1(_07499_),
    .A2(net167),
    .A3(net281),
    .B1(_04217_),
    .B2(net21),
    .X(_00064_));
 sky130_fd_sc_hd__nor2_1 _23312_ (.A(_04245_),
    .B(_03737_),
    .Y(_00065_));
 sky130_fd_sc_hd__a31oi_4 _23313_ (.A1(_07771_),
    .A2(_03704_),
    .A3(net165),
    .B1(_00065_),
    .Y(_00067_));
 sky130_fd_sc_hd__or3b_2 _23314_ (.A(net38),
    .B(_04256_),
    .C_N(net37),
    .X(_00068_));
 sky130_fd_sc_hd__o211ai_2 _23315_ (.A1(net168),
    .A2(net268),
    .B1(_02858_),
    .C1(net164),
    .Y(_00069_));
 sky130_fd_sc_hd__o311a_1 _23316_ (.A1(_02869_),
    .A2(_08203_),
    .A3(net154),
    .B1(_00068_),
    .C1(_00067_),
    .X(_00070_));
 sky130_fd_sc_hd__o221ai_4 _23317_ (.A1(_04256_),
    .A2(_02891_),
    .B1(_08209_),
    .B2(_02869_),
    .C1(_00067_),
    .Y(_00071_));
 sky130_fd_sc_hd__a21oi_4 _23318_ (.A1(_00068_),
    .A2(_00069_),
    .B1(_00067_),
    .Y(_00072_));
 sky130_fd_sc_hd__a21o_1 _23319_ (.A1(_00068_),
    .A2(_00069_),
    .B1(_00067_),
    .X(_00073_));
 sky130_fd_sc_hd__nand3_4 _23320_ (.A(_00064_),
    .B(_00071_),
    .C(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_2 _23321_ (.A(_00074_),
    .Y(_00075_));
 sky130_fd_sc_hd__o21bai_4 _23322_ (.A1(_00070_),
    .A2(_00072_),
    .B1_N(_00064_),
    .Y(_00076_));
 sky130_fd_sc_hd__a21oi_2 _23323_ (.A1(_13071_),
    .A2(_13074_),
    .B1(_13068_),
    .Y(_00078_));
 sky130_fd_sc_hd__o21ai_1 _23324_ (.A1(_13067_),
    .A2(_13078_),
    .B1(_13077_),
    .Y(_00079_));
 sky130_fd_sc_hd__a21oi_2 _23325_ (.A1(_00074_),
    .A2(_00076_),
    .B1(_00079_),
    .Y(_00080_));
 sky130_fd_sc_hd__o2bb2ai_4 _23326_ (.A1_N(_00074_),
    .A2_N(_00076_),
    .B1(_00078_),
    .B2(_13078_),
    .Y(_00081_));
 sky130_fd_sc_hd__o211ai_4 _23327_ (.A1(_13076_),
    .A2(_13081_),
    .B1(_00074_),
    .C1(_00076_),
    .Y(_00082_));
 sky130_fd_sc_hd__inv_2 _23328_ (.A(_00082_),
    .Y(_00083_));
 sky130_fd_sc_hd__o221a_2 _23329_ (.A1(_04212_),
    .A2(_04218_),
    .B1(_07079_),
    .B2(_04216_),
    .C1(_13157_),
    .X(_00084_));
 sky130_fd_sc_hd__o21a_1 _23330_ (.A1(_13148_),
    .A2(_13158_),
    .B1(_13157_),
    .X(_00085_));
 sky130_fd_sc_hd__nand3b_4 _23331_ (.A_N(_00085_),
    .B(_00082_),
    .C(_00081_),
    .Y(_00086_));
 sky130_fd_sc_hd__o2bb2ai_4 _23332_ (.A1_N(_00081_),
    .A2_N(_00082_),
    .B1(_00084_),
    .B2(_13158_),
    .Y(_00087_));
 sky130_fd_sc_hd__o311a_1 _23333_ (.A1(_13161_),
    .A2(_13164_),
    .A3(_13167_),
    .B1(_12890_),
    .C1(_12886_),
    .X(_00089_));
 sky130_fd_sc_hd__a2bb2o_2 _23334_ (.A1_N(_13164_),
    .A2_N(_13170_),
    .B1(_13172_),
    .B2(_13168_),
    .X(_00090_));
 sky130_fd_sc_hd__a21oi_2 _23335_ (.A1(_00086_),
    .A2(_00087_),
    .B1(_00090_),
    .Y(_00091_));
 sky130_fd_sc_hd__o2bb2ai_4 _23336_ (.A1_N(_00086_),
    .A2_N(_00087_),
    .B1(_00089_),
    .B2(_13169_),
    .Y(_00092_));
 sky130_fd_sc_hd__and3_1 _23337_ (.A(_00090_),
    .B(_00087_),
    .C(_00086_),
    .X(_00093_));
 sky130_fd_sc_hd__nand3_4 _23338_ (.A(_00090_),
    .B(_00087_),
    .C(_00086_),
    .Y(_00094_));
 sky130_fd_sc_hd__a32o_1 _23339_ (.A1(net178),
    .A2(net177),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net15),
    .X(_00095_));
 sky130_fd_sc_hd__a32oi_4 _23340_ (.A1(net202),
    .A2(net173),
    .A3(net242),
    .B1(_04988_),
    .B2(net17),
    .Y(_00096_));
 sky130_fd_sc_hd__a211o_1 _23341_ (.A1(net177),
    .A2(net16),
    .B1(_05226_),
    .C1(net203),
    .X(_00097_));
 sky130_fd_sc_hd__or3_1 _23342_ (.A(net46),
    .B(_04157_),
    .C(_04124_),
    .X(_00098_));
 sky130_fd_sc_hd__o221a_1 _23343_ (.A1(_04157_),
    .A2(_05229_),
    .B1(_05935_),
    .B2(_05226_),
    .C1(_00096_),
    .X(_00100_));
 sky130_fd_sc_hd__o221ai_4 _23344_ (.A1(_04157_),
    .A2(_05229_),
    .B1(_05935_),
    .B2(_05226_),
    .C1(_00096_),
    .Y(_00101_));
 sky130_fd_sc_hd__a21oi_1 _23345_ (.A1(_00097_),
    .A2(_00098_),
    .B1(_00096_),
    .Y(_00102_));
 sky130_fd_sc_hd__nor2_1 _23346_ (.A(_00095_),
    .B(_00102_),
    .Y(_00103_));
 sky130_fd_sc_hd__a21o_1 _23347_ (.A1(_00095_),
    .A2(_00101_),
    .B1(_00102_),
    .X(_00104_));
 sky130_fd_sc_hd__nand2_1 _23348_ (.A(_00102_),
    .B(_00095_),
    .Y(_00105_));
 sky130_fd_sc_hd__a2bb2oi_2 _23349_ (.A1_N(_00095_),
    .A2_N(_00101_),
    .B1(_00105_),
    .B2(_00104_),
    .Y(_00106_));
 sky130_fd_sc_hd__a21oi_1 _23350_ (.A1(_13200_),
    .A2(_13206_),
    .B1(_13208_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3_1 _23351_ (.A(_04102_),
    .B(net18),
    .C(net42),
    .X(_00108_));
 sky130_fd_sc_hd__o311a_1 _23352_ (.A1(net246),
    .A2(_05928_),
    .A3(_06451_),
    .B1(_04895_),
    .C1(net197),
    .X(_00109_));
 sky130_fd_sc_hd__a31o_1 _23353_ (.A1(net197),
    .A2(net172),
    .A3(_04895_),
    .B1(_00108_),
    .X(_00111_));
 sky130_fd_sc_hd__or3b_1 _23354_ (.A(net42),
    .B(_04201_),
    .C_N(net41),
    .X(_00112_));
 sky130_fd_sc_hd__o211ai_4 _23355_ (.A1(net174),
    .A2(_06759_),
    .B1(_04480_),
    .C1(net194),
    .Y(_00113_));
 sky130_fd_sc_hd__a221oi_4 _23356_ (.A1(net203),
    .A2(net272),
    .B1(net171),
    .B2(net20),
    .C1(_04268_),
    .Y(_00114_));
 sky130_fd_sc_hd__nor2_2 _23357_ (.A(_04212_),
    .B(_04270_),
    .Y(_00115_));
 sky130_fd_sc_hd__a31oi_2 _23358_ (.A1(_07072_),
    .A2(net168),
    .A3(_04267_),
    .B1(_00115_),
    .Y(_00116_));
 sky130_fd_sc_hd__o221ai_4 _23359_ (.A1(_04212_),
    .A2(_04270_),
    .B1(_04483_),
    .B2(_04201_),
    .C1(_00113_),
    .Y(_00117_));
 sky130_fd_sc_hd__o221ai_4 _23360_ (.A1(_04201_),
    .A2(_04483_),
    .B1(_06764_),
    .B2(_04481_),
    .C1(_00116_),
    .Y(_00118_));
 sky130_fd_sc_hd__o2bb2a_1 _23361_ (.A1_N(_00112_),
    .A2_N(_00113_),
    .B1(_00114_),
    .B2(_00115_),
    .X(_00119_));
 sky130_fd_sc_hd__o2bb2ai_4 _23362_ (.A1_N(_00112_),
    .A2_N(_00113_),
    .B1(_00114_),
    .B2(_00115_),
    .Y(_00120_));
 sky130_fd_sc_hd__o21a_1 _23363_ (.A1(_00114_),
    .A2(_00117_),
    .B1(_00120_),
    .X(_00122_));
 sky130_fd_sc_hd__o221a_2 _23364_ (.A1(_00108_),
    .A2(_00109_),
    .B1(_00114_),
    .B2(_00117_),
    .C1(_00120_),
    .X(_00123_));
 sky130_fd_sc_hd__o221ai_2 _23365_ (.A1(_00108_),
    .A2(_00109_),
    .B1(_00114_),
    .B2(_00117_),
    .C1(_00120_),
    .Y(_00124_));
 sky130_fd_sc_hd__a21oi_2 _23366_ (.A1(_00118_),
    .A2(_00120_),
    .B1(_00111_),
    .Y(_00125_));
 sky130_fd_sc_hd__o21bai_1 _23367_ (.A1(_00111_),
    .A2(_00122_),
    .B1_N(_00107_),
    .Y(_00126_));
 sky130_fd_sc_hd__a211oi_4 _23368_ (.A1(_13209_),
    .A2(_13210_),
    .B1(_00123_),
    .C1(_00125_),
    .Y(_00127_));
 sky130_fd_sc_hd__o211a_1 _23369_ (.A1(_00123_),
    .A2(_00125_),
    .B1(_13209_),
    .C1(_13210_),
    .X(_00128_));
 sky130_fd_sc_hd__o21ai_2 _23370_ (.A1(_00123_),
    .A2(_00125_),
    .B1(_00107_),
    .Y(_00129_));
 sky130_fd_sc_hd__nand2_2 _23371_ (.A(_00129_),
    .B(_00106_),
    .Y(_00130_));
 sky130_fd_sc_hd__o211a_1 _23372_ (.A1(_00123_),
    .A2(_00126_),
    .B1(_00129_),
    .C1(_00106_),
    .X(_00131_));
 sky130_fd_sc_hd__o21bai_4 _23373_ (.A1(_00127_),
    .A2(_00128_),
    .B1_N(_00106_),
    .Y(_00133_));
 sky130_fd_sc_hd__inv_2 _23374_ (.A(_00133_),
    .Y(_00134_));
 sky130_fd_sc_hd__o21ai_2 _23375_ (.A1(_00127_),
    .A2(_00130_),
    .B1(_00133_),
    .Y(_00135_));
 sky130_fd_sc_hd__o2111ai_4 _23376_ (.A1(_00127_),
    .A2(_00130_),
    .B1(_00133_),
    .C1(_00094_),
    .D1(_00092_),
    .Y(_00136_));
 sky130_fd_sc_hd__o2bb2ai_4 _23377_ (.A1_N(_00092_),
    .A2_N(_00094_),
    .B1(_00131_),
    .B2(_00134_),
    .Y(_00137_));
 sky130_fd_sc_hd__o311a_1 _23378_ (.A1(_10324_),
    .A2(_08668_),
    .A3(_12453_),
    .B1(_12993_),
    .C1(_13091_),
    .X(_00138_));
 sky130_fd_sc_hd__o21ai_2 _23379_ (.A1(_13062_),
    .A2(_13088_),
    .B1(_13091_),
    .Y(_00139_));
 sky130_fd_sc_hd__a21oi_4 _23380_ (.A1(_00136_),
    .A2(_00137_),
    .B1(_00139_),
    .Y(_00140_));
 sky130_fd_sc_hd__o2bb2ai_4 _23381_ (.A1_N(_00136_),
    .A2_N(_00137_),
    .B1(_00138_),
    .B2(_13088_),
    .Y(_00141_));
 sky130_fd_sc_hd__o211a_1 _23382_ (.A1(_13090_),
    .A2(_13093_),
    .B1(_00136_),
    .C1(_00137_),
    .X(_00142_));
 sky130_fd_sc_hd__o211ai_4 _23383_ (.A1(_13090_),
    .A2(_13093_),
    .B1(_00136_),
    .C1(_00137_),
    .Y(_00144_));
 sky130_fd_sc_hd__and3_1 _23384_ (.A(_13180_),
    .B(_13217_),
    .C(_13220_),
    .X(_00145_));
 sky130_fd_sc_hd__o21ai_2 _23385_ (.A1(_13178_),
    .A2(_13225_),
    .B1(_13180_),
    .Y(_00146_));
 sky130_fd_sc_hd__o2bb2ai_2 _23386_ (.A1_N(_00141_),
    .A2_N(_00144_),
    .B1(_00145_),
    .B2(_13178_),
    .Y(_00147_));
 sky130_fd_sc_hd__o211ai_2 _23387_ (.A1(_13181_),
    .A2(_13230_),
    .B1(_00141_),
    .C1(_00144_),
    .Y(_00148_));
 sky130_fd_sc_hd__o22ai_4 _23388_ (.A1(_13181_),
    .A2(_13230_),
    .B1(_00140_),
    .B2(_00142_),
    .Y(_00149_));
 sky130_fd_sc_hd__o2111ai_4 _23389_ (.A1(_13178_),
    .A2(_13225_),
    .B1(_00141_),
    .C1(_00144_),
    .D1(_13180_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand3_1 _23390_ (.A(_00063_),
    .B(_00149_),
    .C(_00150_),
    .Y(_00151_));
 sky130_fd_sc_hd__nand3_2 _23391_ (.A(_00062_),
    .B(_00147_),
    .C(_00148_),
    .Y(_00152_));
 sky130_fd_sc_hd__nand4_1 _23392_ (.A(_00061_),
    .B(_00062_),
    .C(_00147_),
    .D(_00148_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand4_4 _23393_ (.A(_00061_),
    .B(_00062_),
    .C(_00149_),
    .D(_00150_),
    .Y(_00155_));
 sky130_fd_sc_hd__nand3_2 _23394_ (.A(_00063_),
    .B(_00147_),
    .C(_00148_),
    .Y(_00156_));
 sky130_fd_sc_hd__nand2_1 _23395_ (.A(_00151_),
    .B(_00153_),
    .Y(_00157_));
 sky130_fd_sc_hd__a22oi_4 _23396_ (.A1(_13142_),
    .A2(_13373_),
    .B1(_00155_),
    .B2(_00156_),
    .Y(_00158_));
 sky130_fd_sc_hd__nand3_1 _23397_ (.A(_13374_),
    .B(_00151_),
    .C(_00153_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand3_2 _23398_ (.A(_13375_),
    .B(_00155_),
    .C(_00156_),
    .Y(_00160_));
 sky130_fd_sc_hd__a21boi_1 _23399_ (.A1(_13277_),
    .A2(_13281_),
    .B1_N(_13279_),
    .Y(_00161_));
 sky130_fd_sc_hd__o2bb2ai_2 _23400_ (.A1_N(_13281_),
    .A2_N(_13277_),
    .B1(_13274_),
    .B2(_13278_),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _23401_ (.A(_13270_),
    .B(_13275_),
    .Y(_00163_));
 sky130_fd_sc_hd__a32oi_4 _23402_ (.A1(_13199_),
    .A2(_13210_),
    .A3(_13211_),
    .B1(_13195_),
    .B2(_13193_),
    .Y(_00164_));
 sky130_fd_sc_hd__a32o_1 _23403_ (.A1(_13199_),
    .A2(_13210_),
    .A3(_13211_),
    .B1(_13195_),
    .B2(_13193_),
    .X(_00166_));
 sky130_fd_sc_hd__a21o_1 _23404_ (.A1(_13263_),
    .A2(_13264_),
    .B1(_13260_),
    .X(_00167_));
 sky130_fd_sc_hd__a21oi_2 _23405_ (.A1(_13187_),
    .A2(_13190_),
    .B1(_13183_),
    .Y(_00168_));
 sky130_fd_sc_hd__a21oi_2 _23406_ (.A1(_13186_),
    .A2(_13189_),
    .B1(_13182_),
    .Y(_00169_));
 sky130_fd_sc_hd__o311a_1 _23407_ (.A1(net7),
    .A2(net248),
    .A3(_04787_),
    .B1(net273),
    .C1(net213),
    .X(_00170_));
 sky130_fd_sc_hd__and3_1 _23408_ (.A(_04190_),
    .B(net49),
    .C(net11),
    .X(_00171_));
 sky130_fd_sc_hd__a21oi_1 _23409_ (.A1(_04792_),
    .A2(net273),
    .B1(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__a31o_1 _23410_ (.A1(net184),
    .A2(net213),
    .A3(net273),
    .B1(_00171_),
    .X(_00173_));
 sky130_fd_sc_hd__nand3_2 _23411_ (.A(_05290_),
    .B(_05292_),
    .C(_05762_),
    .Y(_00174_));
 sky130_fd_sc_hd__or3b_2 _23412_ (.A(_04135_),
    .B(net48),
    .C_N(net47),
    .X(_00175_));
 sky130_fd_sc_hd__nor2_2 _23413_ (.A(_04113_),
    .B(_06030_),
    .Y(_00177_));
 sky130_fd_sc_hd__o311a_1 _23414_ (.A1(net11),
    .A2(_04557_),
    .A3(net208),
    .B1(net274),
    .C1(net209),
    .X(_00178_));
 sky130_fd_sc_hd__o211ai_1 _23415_ (.A1(_04787_),
    .A2(net208),
    .B1(net274),
    .C1(net209),
    .Y(_00179_));
 sky130_fd_sc_hd__a31oi_1 _23416_ (.A1(net209),
    .A2(_05074_),
    .A3(net274),
    .B1(_00177_),
    .Y(_00180_));
 sky130_fd_sc_hd__nand3_2 _23417_ (.A(_00174_),
    .B(_00175_),
    .C(_00179_),
    .Y(_00181_));
 sky130_fd_sc_hd__o211ai_2 _23418_ (.A1(_04135_),
    .A2(_05766_),
    .B1(_00174_),
    .C1(_00180_),
    .Y(_00182_));
 sky130_fd_sc_hd__o2bb2a_1 _23419_ (.A1_N(_00174_),
    .A2_N(_00175_),
    .B1(_00177_),
    .B2(_00178_),
    .X(_00183_));
 sky130_fd_sc_hd__o2bb2ai_4 _23420_ (.A1_N(_00174_),
    .A2_N(_00175_),
    .B1(_00177_),
    .B2(_00178_),
    .Y(_00184_));
 sky130_fd_sc_hd__o21ai_1 _23421_ (.A1(_00177_),
    .A2(_00181_),
    .B1(_00184_),
    .Y(_00185_));
 sky130_fd_sc_hd__o221a_2 _23422_ (.A1(_00170_),
    .A2(_00171_),
    .B1(_00177_),
    .B2(_00181_),
    .C1(_00184_),
    .X(_00186_));
 sky130_fd_sc_hd__o221ai_4 _23423_ (.A1(_00170_),
    .A2(_00171_),
    .B1(_00177_),
    .B2(_00181_),
    .C1(_00184_),
    .Y(_00188_));
 sky130_fd_sc_hd__a21oi_1 _23424_ (.A1(_00182_),
    .A2(_00184_),
    .B1(_00173_),
    .Y(_00189_));
 sky130_fd_sc_hd__a21o_1 _23425_ (.A1(_00182_),
    .A2(_00184_),
    .B1(_00173_),
    .X(_00190_));
 sky130_fd_sc_hd__o2bb2ai_1 _23426_ (.A1_N(_00172_),
    .A2_N(_00185_),
    .B1(_13191_),
    .B2(_00169_),
    .Y(_00191_));
 sky130_fd_sc_hd__o211a_2 _23427_ (.A1(_13191_),
    .A2(_00169_),
    .B1(_00188_),
    .C1(_00190_),
    .X(_00192_));
 sky130_fd_sc_hd__o211ai_2 _23428_ (.A1(_13191_),
    .A2(_00169_),
    .B1(_00188_),
    .C1(_00190_),
    .Y(_00193_));
 sky130_fd_sc_hd__o22ai_4 _23429_ (.A1(_13192_),
    .A2(_00168_),
    .B1(_00186_),
    .B2(_00189_),
    .Y(_00194_));
 sky130_fd_sc_hd__o21ai_2 _23430_ (.A1(_13260_),
    .A2(_13267_),
    .B1(_00194_),
    .Y(_00195_));
 sky130_fd_sc_hd__inv_2 _23431_ (.A(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__o221a_1 _23432_ (.A1(_13260_),
    .A2(_13267_),
    .B1(_00186_),
    .B2(_00191_),
    .C1(_00194_),
    .X(_00197_));
 sky130_fd_sc_hd__a21oi_2 _23433_ (.A1(_00193_),
    .A2(_00194_),
    .B1(_00167_),
    .Y(_00199_));
 sky130_fd_sc_hd__a21o_1 _23434_ (.A1(_00193_),
    .A2(_00194_),
    .B1(_00167_),
    .X(_00200_));
 sky130_fd_sc_hd__o2111a_1 _23435_ (.A1(_00195_),
    .A2(_00192_),
    .B1(_00166_),
    .C1(_13215_),
    .D1(_00200_),
    .X(_00201_));
 sky130_fd_sc_hd__o2111ai_4 _23436_ (.A1(_00195_),
    .A2(_00192_),
    .B1(_00166_),
    .C1(_13215_),
    .D1(_00200_),
    .Y(_00202_));
 sky130_fd_sc_hd__o221a_1 _23437_ (.A1(_13198_),
    .A2(_13214_),
    .B1(_00197_),
    .B2(_00199_),
    .C1(_13213_),
    .X(_00203_));
 sky130_fd_sc_hd__o22ai_4 _23438_ (.A1(_13214_),
    .A2(_00164_),
    .B1(_00197_),
    .B2(_00199_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _23439_ (.A(_00163_),
    .B(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__a21o_1 _23440_ (.A1(_00202_),
    .A2(_00204_),
    .B1(_00163_),
    .X(_00206_));
 sky130_fd_sc_hd__nand4_2 _23441_ (.A(_13270_),
    .B(_13275_),
    .C(_00202_),
    .D(_00204_),
    .Y(_00207_));
 sky130_fd_sc_hd__a22o_1 _23442_ (.A1(_13270_),
    .A2(_13275_),
    .B1(_00202_),
    .B2(_00204_),
    .X(_00208_));
 sky130_fd_sc_hd__nand3_4 _23443_ (.A(_00208_),
    .B(_00161_),
    .C(_00207_),
    .Y(_00210_));
 sky130_fd_sc_hd__o211ai_4 _23444_ (.A1(_00205_),
    .A2(_00201_),
    .B1(_00162_),
    .C1(_00206_),
    .Y(_00211_));
 sky130_fd_sc_hd__o311a_1 _23445_ (.A1(net259),
    .A2(_11387_),
    .A3(_02442_),
    .B1(net238),
    .C1(_02421_),
    .X(_00212_));
 sky130_fd_sc_hd__and3_1 _23446_ (.A(_04266_),
    .B(net54),
    .C(net6),
    .X(_00213_));
 sky130_fd_sc_hd__o2bb2a_1 _23447_ (.A1_N(_02464_),
    .A2_N(net238),
    .B1(_08007_),
    .B2(_04026_),
    .X(_00214_));
 sky130_fd_sc_hd__a31o_1 _23448_ (.A1(_02421_),
    .A2(net248),
    .A3(net238),
    .B1(_00213_),
    .X(_00215_));
 sky130_fd_sc_hd__nand2_1 _23449_ (.A(_13302_),
    .B(_13305_),
    .Y(_00216_));
 sky130_fd_sc_hd__a22oi_2 _23450_ (.A1(_03959_),
    .A2(_07642_),
    .B1(_07643_),
    .B2(net7),
    .Y(_00217_));
 sky130_fd_sc_hd__a32o_1 _23451_ (.A1(_03952_),
    .A2(net233),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net7),
    .X(_00218_));
 sky130_fd_sc_hd__a21o_1 _23452_ (.A1(_13294_),
    .A2(_13296_),
    .B1(_13291_),
    .X(_00219_));
 sky130_fd_sc_hd__a32oi_4 _23453_ (.A1(net229),
    .A2(net227),
    .A3(net239),
    .B1(_07308_),
    .B2(net8),
    .Y(_00221_));
 sky130_fd_sc_hd__o31a_1 _23454_ (.A1(net259),
    .A2(_03956_),
    .A3(_04407_),
    .B1(net269),
    .X(_00222_));
 sky130_fd_sc_hd__a22oi_4 _23455_ (.A1(net9),
    .A2(_07225_),
    .B1(_00222_),
    .B2(net225),
    .Y(_00223_));
 sky130_fd_sc_hd__o211ai_2 _23456_ (.A1(net233),
    .A2(_04557_),
    .B1(net240),
    .C1(net217),
    .Y(_00224_));
 sky130_fd_sc_hd__or3_1 _23457_ (.A(net51),
    .B(_04190_),
    .C(_04080_),
    .X(_00225_));
 sky130_fd_sc_hd__o32a_1 _23458_ (.A1(_06864_),
    .A2(net216),
    .A3(_04554_),
    .B1(_04080_),
    .B2(_06866_),
    .X(_00226_));
 sky130_fd_sc_hd__a21oi_1 _23459_ (.A1(_00224_),
    .A2(_00225_),
    .B1(_00223_),
    .Y(_00227_));
 sky130_fd_sc_hd__a21o_1 _23460_ (.A1(_00224_),
    .A2(_00225_),
    .B1(_00223_),
    .X(_00228_));
 sky130_fd_sc_hd__o311a_2 _23461_ (.A1(_04080_),
    .A2(_04190_),
    .A3(net51),
    .B1(_00224_),
    .C1(_00223_),
    .X(_00229_));
 sky130_fd_sc_hd__nand2_1 _23462_ (.A(_00223_),
    .B(_00226_),
    .Y(_00230_));
 sky130_fd_sc_hd__o21ai_1 _23463_ (.A1(_00227_),
    .A2(_00229_),
    .B1(_00221_),
    .Y(_00232_));
 sky130_fd_sc_hd__o21bai_2 _23464_ (.A1(_00223_),
    .A2(_00226_),
    .B1_N(_00221_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand3_1 _23465_ (.A(_00230_),
    .B(_00221_),
    .C(_00228_),
    .Y(_00234_));
 sky130_fd_sc_hd__o21bai_1 _23466_ (.A1(_00227_),
    .A2(_00229_),
    .B1_N(_00221_),
    .Y(_00235_));
 sky130_fd_sc_hd__o211ai_4 _23467_ (.A1(_00233_),
    .A2(_00229_),
    .B1(_00219_),
    .C1(_00232_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand4_4 _23468_ (.A(_13292_),
    .B(_13298_),
    .C(_00234_),
    .D(_00235_),
    .Y(_00237_));
 sky130_fd_sc_hd__a21o_1 _23469_ (.A1(_00236_),
    .A2(_00237_),
    .B1(_00218_),
    .X(_00238_));
 sky130_fd_sc_hd__nand3_1 _23470_ (.A(_00218_),
    .B(_00236_),
    .C(_00237_),
    .Y(_00239_));
 sky130_fd_sc_hd__a21o_1 _23471_ (.A1(_00236_),
    .A2(_00237_),
    .B1(_00217_),
    .X(_00240_));
 sky130_fd_sc_hd__nand3_2 _23472_ (.A(_00237_),
    .B(_00217_),
    .C(_00236_),
    .Y(_00241_));
 sky130_fd_sc_hd__a22oi_4 _23473_ (.A1(_13302_),
    .A2(_13305_),
    .B1(_00240_),
    .B2(_00241_),
    .Y(_00243_));
 sky130_fd_sc_hd__a22o_1 _23474_ (.A1(_13302_),
    .A2(_13305_),
    .B1(_00240_),
    .B2(_00241_),
    .X(_00244_));
 sky130_fd_sc_hd__a21oi_2 _23475_ (.A1(_00238_),
    .A2(_00239_),
    .B1(_00216_),
    .Y(_00245_));
 sky130_fd_sc_hd__a21o_1 _23476_ (.A1(_00238_),
    .A2(_00239_),
    .B1(_00216_),
    .X(_00246_));
 sky130_fd_sc_hd__o21a_1 _23477_ (.A1(_00243_),
    .A2(_00245_),
    .B1(_00214_),
    .X(_00247_));
 sky130_fd_sc_hd__and3_1 _23478_ (.A(_00215_),
    .B(_00244_),
    .C(_00246_),
    .X(_00248_));
 sky130_fd_sc_hd__o22a_1 _23479_ (.A1(_00212_),
    .A2(_00213_),
    .B1(_00243_),
    .B2(_00245_),
    .X(_00249_));
 sky130_fd_sc_hd__o21ai_1 _23480_ (.A1(_00243_),
    .A2(_00245_),
    .B1(_00215_),
    .Y(_00250_));
 sky130_fd_sc_hd__and3_1 _23481_ (.A(_00246_),
    .B(_00214_),
    .C(_00244_),
    .X(_00251_));
 sky130_fd_sc_hd__nand3_1 _23482_ (.A(_00246_),
    .B(_00214_),
    .C(_00244_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _23483_ (.A(_00250_),
    .B(_00252_),
    .Y(_00254_));
 sky130_fd_sc_hd__a21oi_1 _23484_ (.A1(_00210_),
    .A2(_00211_),
    .B1(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__o2bb2ai_1 _23485_ (.A1_N(_00210_),
    .A2_N(_00211_),
    .B1(_00247_),
    .B2(_00248_),
    .Y(_00256_));
 sky130_fd_sc_hd__o211a_1 _23486_ (.A1(_00249_),
    .A2(_00251_),
    .B1(_00210_),
    .C1(_00211_),
    .X(_00257_));
 sky130_fd_sc_hd__o211ai_4 _23487_ (.A1(_00249_),
    .A2(_00251_),
    .B1(_00210_),
    .C1(_00211_),
    .Y(_00258_));
 sky130_fd_sc_hd__a32oi_4 _23488_ (.A1(_13144_),
    .A2(_13228_),
    .A3(_13231_),
    .B1(_13233_),
    .B2(_13236_),
    .Y(_00259_));
 sky130_fd_sc_hd__o2bb2ai_2 _23489_ (.A1_N(_13236_),
    .A2_N(_13233_),
    .B1(_13234_),
    .B2(_13232_),
    .Y(_00260_));
 sky130_fd_sc_hd__a21oi_2 _23490_ (.A1(_00256_),
    .A2(_00258_),
    .B1(_00260_),
    .Y(_00261_));
 sky130_fd_sc_hd__o21ai_1 _23491_ (.A1(_00255_),
    .A2(_00257_),
    .B1(_00259_),
    .Y(_00262_));
 sky130_fd_sc_hd__nor3_2 _23492_ (.A(_00255_),
    .B(_00257_),
    .C(_00259_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand3_1 _23493_ (.A(_00256_),
    .B(_00258_),
    .C(_00260_),
    .Y(_00265_));
 sky130_fd_sc_hd__o21ai_2 _23494_ (.A1(_13312_),
    .A2(_13313_),
    .B1(_13286_),
    .Y(_00266_));
 sky130_fd_sc_hd__a21oi_1 _23495_ (.A1(_00262_),
    .A2(_00265_),
    .B1(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__o21bai_2 _23496_ (.A1(_00261_),
    .A2(_00263_),
    .B1_N(_00266_),
    .Y(_00268_));
 sky130_fd_sc_hd__a21oi_2 _23497_ (.A1(_13286_),
    .A2(_13315_),
    .B1(_00261_),
    .Y(_00269_));
 sky130_fd_sc_hd__and3_1 _23498_ (.A(_00262_),
    .B(_00265_),
    .C(_00266_),
    .X(_00270_));
 sky130_fd_sc_hd__nand3_1 _23499_ (.A(_00262_),
    .B(_00265_),
    .C(_00266_),
    .Y(_00271_));
 sky130_fd_sc_hd__o2bb2ai_2 _23500_ (.A1_N(_00159_),
    .A2_N(_00160_),
    .B1(_00267_),
    .B2(_00270_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand3_2 _23501_ (.A(_00160_),
    .B(_00268_),
    .C(_00271_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand4_1 _23502_ (.A(_00159_),
    .B(_00160_),
    .C(_00268_),
    .D(_00271_),
    .Y(_00274_));
 sky130_fd_sc_hd__o21ai_1 _23503_ (.A1(_00158_),
    .A2(_00273_),
    .B1(_00272_),
    .Y(_00276_));
 sky130_fd_sc_hd__a21oi_2 _23504_ (.A1(_00272_),
    .A2(_00274_),
    .B1(_13372_),
    .Y(_00277_));
 sky130_fd_sc_hd__a21o_1 _23505_ (.A1(_00272_),
    .A2(_00274_),
    .B1(_13372_),
    .X(_00278_));
 sky130_fd_sc_hd__o211a_2 _23506_ (.A1(_00158_),
    .A2(_00273_),
    .B1(_00272_),
    .C1(_13372_),
    .X(_00279_));
 sky130_fd_sc_hd__o211ai_1 _23507_ (.A1(_00158_),
    .A2(_00273_),
    .B1(_00272_),
    .C1(_13372_),
    .Y(_00280_));
 sky130_fd_sc_hd__o21ai_2 _23508_ (.A1(_00277_),
    .A2(_00279_),
    .B1(_13369_),
    .Y(_00281_));
 sky130_fd_sc_hd__a2bb2oi_1 _23509_ (.A1_N(_13322_),
    .A2_N(_13327_),
    .B1(_13370_),
    .B2(_00276_),
    .Y(_00282_));
 sky130_fd_sc_hd__o2bb2ai_2 _23510_ (.A1_N(_13370_),
    .A2_N(_00276_),
    .B1(_13322_),
    .B2(_13327_),
    .Y(_00283_));
 sky130_fd_sc_hd__o22ai_2 _23511_ (.A1(_13322_),
    .A2(_13327_),
    .B1(_00277_),
    .B2(_00279_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand3_1 _23512_ (.A(_00278_),
    .B(_00280_),
    .C(_13369_),
    .Y(_00285_));
 sky130_fd_sc_hd__o21ai_1 _23513_ (.A1(_12821_),
    .A2(_13341_),
    .B1(_13338_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _23514_ (.A(_13340_),
    .B(_00287_),
    .Y(_00288_));
 sky130_fd_sc_hd__o221a_2 _23515_ (.A1(_00279_),
    .A2(_00283_),
    .B1(_13337_),
    .B2(_13347_),
    .C1(_00281_),
    .X(_00289_));
 sky130_fd_sc_hd__o221ai_4 _23516_ (.A1(_00279_),
    .A2(_00283_),
    .B1(_13337_),
    .B2(_13347_),
    .C1(_00281_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand3_1 _23517_ (.A(_00284_),
    .B(_00285_),
    .C(_00288_),
    .Y(_00291_));
 sky130_fd_sc_hd__a21o_1 _23518_ (.A1(_00290_),
    .A2(_00291_),
    .B1(_13367_),
    .X(_00292_));
 sky130_fd_sc_hd__a31oi_2 _23519_ (.A1(_00284_),
    .A2(_00285_),
    .A3(_00288_),
    .B1(_13368_),
    .Y(_00293_));
 sky130_fd_sc_hd__a31o_1 _23520_ (.A1(_00284_),
    .A2(_00285_),
    .A3(_00288_),
    .B1(_13368_),
    .X(_00294_));
 sky130_fd_sc_hd__nand3_1 _23521_ (.A(_00290_),
    .B(_00291_),
    .C(_13368_),
    .Y(_00295_));
 sky130_fd_sc_hd__a21o_1 _23522_ (.A1(_00290_),
    .A2(_00291_),
    .B1(_13368_),
    .X(_00296_));
 sky130_fd_sc_hd__nand4_1 _23523_ (.A(_13352_),
    .B(_13356_),
    .C(_00295_),
    .D(_00296_),
    .Y(_00298_));
 sky130_fd_sc_hd__o221a_1 _23524_ (.A1(_13351_),
    .A2(_13355_),
    .B1(_00289_),
    .B2(_00294_),
    .C1(_00292_),
    .X(_00299_));
 sky130_fd_sc_hd__o221ai_4 _23525_ (.A1(_00289_),
    .A2(_00294_),
    .B1(_13351_),
    .B2(_13355_),
    .C1(_00292_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _23526_ (.A(_00298_),
    .B(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand4_4 _23527_ (.A(_13051_),
    .B(_13052_),
    .C(_13363_),
    .D(_13364_),
    .Y(_00302_));
 sky130_fd_sc_hd__and4_1 _23528_ (.A(_12388_),
    .B(_12389_),
    .C(_12721_),
    .D(_12723_),
    .X(_00303_));
 sky130_fd_sc_hd__or3_1 _23529_ (.A(_12390_),
    .B(_12724_),
    .C(_00302_),
    .X(_00304_));
 sky130_fd_sc_hd__a31oi_2 _23530_ (.A1(_12721_),
    .A2(_12384_),
    .A3(_12387_),
    .B1(_12722_),
    .Y(_00305_));
 sky130_fd_sc_hd__a32oi_4 _23531_ (.A1(_12728_),
    .A2(_13048_),
    .A3(_13050_),
    .B1(_13360_),
    .B2(_13057_),
    .Y(_00306_));
 sky130_fd_sc_hd__o22ai_4 _23532_ (.A1(_13362_),
    .A2(_00306_),
    .B1(_00305_),
    .B2(_00302_),
    .Y(_00307_));
 sky130_fd_sc_hd__o21bai_4 _23533_ (.A1(_00304_),
    .A2(_12402_),
    .B1_N(_00307_),
    .Y(_00309_));
 sky130_fd_sc_hd__xnor2_1 _23534_ (.A(_00301_),
    .B(_00309_),
    .Y(net103));
 sky130_fd_sc_hd__a21oi_1 _23535_ (.A1(_13367_),
    .A2(_00291_),
    .B1(_00289_),
    .Y(_00310_));
 sky130_fd_sc_hd__nor2_1 _23536_ (.A(_00215_),
    .B(_00243_),
    .Y(_00311_));
 sky130_fd_sc_hd__o21a_1 _23537_ (.A1(_00212_),
    .A2(_00213_),
    .B1(_00246_),
    .X(_00312_));
 sky130_fd_sc_hd__a41o_1 _23538_ (.A1(_13302_),
    .A2(_13305_),
    .A3(_00240_),
    .A4(_00241_),
    .B1(_00311_),
    .X(_00313_));
 sky130_fd_sc_hd__o21ai_2 _23539_ (.A1(_13375_),
    .A2(_00157_),
    .B1(_00273_),
    .Y(_00314_));
 sky130_fd_sc_hd__a31oi_1 _23540_ (.A1(_00160_),
    .A2(_00268_),
    .A3(_00271_),
    .B1(_00158_),
    .Y(_00315_));
 sky130_fd_sc_hd__o211ai_2 _23541_ (.A1(_00060_),
    .A2(_00058_),
    .B1(_00150_),
    .C1(_00149_),
    .Y(_00316_));
 sky130_fd_sc_hd__a2bb2o_1 _23542_ (.A1_N(_00016_),
    .A2_N(_00019_),
    .B1(_00018_),
    .B2(_12099_),
    .X(_00317_));
 sky130_fd_sc_hd__nand2_1 _23543_ (.A(net248),
    .B(_08657_),
    .Y(_00319_));
 sky130_fd_sc_hd__o22ai_4 _23544_ (.A1(_04026_),
    .A2(_08660_),
    .B1(_02410_),
    .B2(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__o2111a_2 _23545_ (.A1(net169),
    .A2(net268),
    .B1(net33),
    .C1(_00320_),
    .D1(net319),
    .X(_00321_));
 sky130_fd_sc_hd__a31oi_4 _23546_ (.A1(net161),
    .A2(net33),
    .A3(net319),
    .B1(_00320_),
    .Y(_00322_));
 sky130_fd_sc_hd__o21ai_4 _23547_ (.A1(_00321_),
    .A2(_00322_),
    .B1(net146),
    .Y(_00323_));
 sky130_fd_sc_hd__o22a_1 _23548_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_00320_),
    .B2(net156),
    .X(_00324_));
 sky130_fd_sc_hd__o21ai_2 _23549_ (.A1(_00320_),
    .A2(net156),
    .B1(_09300_),
    .Y(_00325_));
 sky130_fd_sc_hd__o21ai_4 _23550_ (.A1(net146),
    .A2(_13380_),
    .B1(_13379_),
    .Y(_00326_));
 sky130_fd_sc_hd__a21oi_4 _23551_ (.A1(_00323_),
    .A2(_00325_),
    .B1(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__a21o_1 _23552_ (.A1(_00323_),
    .A2(_00325_),
    .B1(_00326_),
    .X(_00328_));
 sky130_fd_sc_hd__o211a_1 _23553_ (.A1(net146),
    .A2(_00322_),
    .B1(_00326_),
    .C1(_00323_),
    .X(_00330_));
 sky130_fd_sc_hd__o211ai_4 _23554_ (.A1(net146),
    .A2(_00322_),
    .B1(_00326_),
    .C1(_00323_),
    .Y(_00331_));
 sky130_fd_sc_hd__o22ai_2 _23555_ (.A1(_10540_),
    .A2(net135),
    .B1(_00327_),
    .B2(_00330_),
    .Y(_00332_));
 sky130_fd_sc_hd__and3_1 _23556_ (.A(_00328_),
    .B(_00331_),
    .C(net133),
    .X(_00333_));
 sky130_fd_sc_hd__nand3_1 _23557_ (.A(_00328_),
    .B(_00331_),
    .C(net133),
    .Y(_00334_));
 sky130_fd_sc_hd__o211ai_2 _23558_ (.A1(_10540_),
    .A2(net135),
    .B1(_00328_),
    .C1(_00331_),
    .Y(_00335_));
 sky130_fd_sc_hd__o21ai_1 _23559_ (.A1(_00327_),
    .A2(_00330_),
    .B1(net133),
    .Y(_00336_));
 sky130_fd_sc_hd__o22ai_2 _23560_ (.A1(_00001_),
    .A2(_00010_),
    .B1(_10546_),
    .B2(_00008_),
    .Y(_00337_));
 sky130_fd_sc_hd__o22a_1 _23561_ (.A1(_00001_),
    .A2(_00010_),
    .B1(_10546_),
    .B2(_00008_),
    .X(_00338_));
 sky130_fd_sc_hd__a21oi_1 _23562_ (.A1(_00332_),
    .A2(_00334_),
    .B1(_00337_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand3_4 _23563_ (.A(_00335_),
    .B(_00336_),
    .C(_00338_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_2 _23564_ (.A(_00332_),
    .B(_00337_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand3_2 _23565_ (.A(_00332_),
    .B(_00334_),
    .C(_00337_),
    .Y(_00343_));
 sky130_fd_sc_hd__o311a_1 _23566_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_00341_),
    .C1(_00343_),
    .X(_00344_));
 sky130_fd_sc_hd__o221ai_4 _23567_ (.A1(_11042_),
    .A2(_11742_),
    .B1(_00333_),
    .B2(_00342_),
    .C1(_00341_),
    .Y(_00345_));
 sky130_fd_sc_hd__a21oi_2 _23568_ (.A1(_00341_),
    .A2(_00343_),
    .B1(_12099_),
    .Y(_00346_));
 sky130_fd_sc_hd__a21o_1 _23569_ (.A1(_00341_),
    .A2(_00343_),
    .B1(_12099_),
    .X(_00347_));
 sky130_fd_sc_hd__nand3_4 _23570_ (.A(_00317_),
    .B(_00345_),
    .C(_00347_),
    .Y(_00348_));
 sky130_fd_sc_hd__o221a_1 _23571_ (.A1(_00019_),
    .A2(_00016_),
    .B1(_00346_),
    .B2(_00344_),
    .C1(_00025_),
    .X(_00349_));
 sky130_fd_sc_hd__o221ai_4 _23572_ (.A1(_00019_),
    .A2(_00016_),
    .B1(_00346_),
    .B2(_00344_),
    .C1(_00025_),
    .Y(_00350_));
 sky130_fd_sc_hd__a21oi_4 _23573_ (.A1(_01293_),
    .A2(net159),
    .B1(_00031_),
    .Y(_00352_));
 sky130_fd_sc_hd__a31o_1 _23574_ (.A1(net319),
    .A2(net161),
    .A3(_01293_),
    .B1(_00031_),
    .X(_00353_));
 sky130_fd_sc_hd__nand2_2 _23575_ (.A(_00037_),
    .B(_00352_),
    .Y(_00354_));
 sky130_fd_sc_hd__a21oi_2 _23576_ (.A1(_13073_),
    .A2(_00036_),
    .B1(_00352_),
    .Y(_00355_));
 sky130_fd_sc_hd__a21o_4 _23577_ (.A1(_13073_),
    .A2(_00036_),
    .B1(_00352_),
    .X(_00356_));
 sky130_fd_sc_hd__and2_4 _23578_ (.A(_00354_),
    .B(_00356_),
    .X(_00357_));
 sky130_fd_sc_hd__nand2_4 _23579_ (.A(_00354_),
    .B(_00356_),
    .Y(_00358_));
 sky130_fd_sc_hd__o211ai_4 _23580_ (.A1(_12451_),
    .A2(_12454_),
    .B1(_00354_),
    .C1(_00356_),
    .Y(_00359_));
 sky130_fd_sc_hd__and3_4 _23581_ (.A(_00358_),
    .B(_12453_),
    .C(_12449_),
    .X(_00360_));
 sky130_fd_sc_hd__inv_2 _23582_ (.A(_00360_),
    .Y(_00361_));
 sky130_fd_sc_hd__a21oi_4 _23583_ (.A1(_00358_),
    .A2(_13065_),
    .B1(_11741_),
    .Y(_00363_));
 sky130_fd_sc_hd__a31o_4 _23584_ (.A1(_00358_),
    .A2(_12453_),
    .A3(_12449_),
    .B1(_11741_),
    .X(_00364_));
 sky130_fd_sc_hd__or3_4 _23585_ (.A(_12451_),
    .B(_12454_),
    .C(_11740_),
    .X(_00365_));
 sky130_fd_sc_hd__and3_4 _23586_ (.A(_11741_),
    .B(_00358_),
    .C(_13065_),
    .X(_00366_));
 sky130_fd_sc_hd__a221o_4 _23587_ (.A1(_11736_),
    .A2(net137),
    .B1(_00356_),
    .B2(_00354_),
    .C1(_13066_),
    .X(_00367_));
 sky130_fd_sc_hd__o21ai_2 _23588_ (.A1(_11740_),
    .A2(_00359_),
    .B1(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__inv_2 _23589_ (.A(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__a21oi_2 _23590_ (.A1(_00359_),
    .A2(net130),
    .B1(_00368_),
    .Y(_00370_));
 sky130_fd_sc_hd__nor2_1 _23591_ (.A(_00041_),
    .B(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__and2_1 _23592_ (.A(_00370_),
    .B(_00041_),
    .X(_00372_));
 sky130_fd_sc_hd__a31oi_4 _23593_ (.A1(_13066_),
    .A2(_00039_),
    .A3(_00040_),
    .B1(_00370_),
    .Y(_00374_));
 sky130_fd_sc_hd__and4_1 _23594_ (.A(_00370_),
    .B(_00040_),
    .C(_00039_),
    .D(_13066_),
    .X(_00375_));
 sky130_fd_sc_hd__o211ai_2 _23595_ (.A1(_00371_),
    .A2(_00372_),
    .B1(_00348_),
    .C1(_00350_),
    .Y(_00376_));
 sky130_fd_sc_hd__o2bb2ai_1 _23596_ (.A1_N(_00348_),
    .A2_N(_00350_),
    .B1(_00374_),
    .B2(_00375_),
    .Y(_00377_));
 sky130_fd_sc_hd__o211ai_2 _23597_ (.A1(_00374_),
    .A2(_00375_),
    .B1(_00348_),
    .C1(_00350_),
    .Y(_00378_));
 sky130_fd_sc_hd__o2bb2ai_1 _23598_ (.A1_N(_00348_),
    .A2_N(_00350_),
    .B1(_00371_),
    .B2(_00372_),
    .Y(_00379_));
 sky130_fd_sc_hd__a21oi_1 _23599_ (.A1(_00051_),
    .A2(_00027_),
    .B1(_00028_),
    .Y(_00380_));
 sky130_fd_sc_hd__nand3_4 _23600_ (.A(_00378_),
    .B(_00379_),
    .C(_00380_),
    .Y(_00381_));
 sky130_fd_sc_hd__o211ai_4 _23601_ (.A1(_00028_),
    .A2(_00056_),
    .B1(_00376_),
    .C1(_00377_),
    .Y(_00382_));
 sky130_fd_sc_hd__a21boi_2 _23602_ (.A1(_00043_),
    .A2(_13085_),
    .B1_N(_00045_),
    .Y(_00383_));
 sky130_fd_sc_hd__inv_2 _23603_ (.A(_00383_),
    .Y(_00384_));
 sky130_fd_sc_hd__o21a_1 _23604_ (.A1(_13158_),
    .A2(_00084_),
    .B1(_00082_),
    .X(_00385_));
 sky130_fd_sc_hd__o21ai_1 _23605_ (.A1(_13158_),
    .A2(_00084_),
    .B1(_00082_),
    .Y(_00386_));
 sky130_fd_sc_hd__nor2_1 _23606_ (.A(_00085_),
    .B(_00080_),
    .Y(_00387_));
 sky130_fd_sc_hd__o31a_1 _23607_ (.A1(_13158_),
    .A2(_00080_),
    .A3(_00084_),
    .B1(_00082_),
    .X(_00388_));
 sky130_fd_sc_hd__a21oi_2 _23608_ (.A1(_00064_),
    .A2(_00071_),
    .B1(_00072_),
    .Y(_00389_));
 sky130_fd_sc_hd__inv_2 _23609_ (.A(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__nor2_1 _23610_ (.A(_04245_),
    .B(_04218_),
    .Y(_00391_));
 sky130_fd_sc_hd__o311a_1 _23611_ (.A1(_03958_),
    .A2(_05927_),
    .A3(_07767_),
    .B1(_07771_),
    .C1(net281),
    .X(_00392_));
 sky130_fd_sc_hd__a31o_2 _23612_ (.A1(_07771_),
    .A2(net281),
    .A3(net165),
    .B1(_00391_),
    .X(_00393_));
 sky130_fd_sc_hd__nor2_2 _23613_ (.A(_04256_),
    .B(_03737_),
    .Y(_00395_));
 sky130_fd_sc_hd__o311a_1 _23614_ (.A1(net176),
    .A2(_07074_),
    .A3(net268),
    .B1(_03704_),
    .C1(net164),
    .X(_00396_));
 sky130_fd_sc_hd__a31oi_2 _23615_ (.A1(net164),
    .A2(net161),
    .A3(_03704_),
    .B1(_00395_),
    .Y(_00397_));
 sky130_fd_sc_hd__and3_2 _23616_ (.A(_04037_),
    .B(net25),
    .C(net37),
    .X(_00398_));
 sky130_fd_sc_hd__a21oi_2 _23617_ (.A1(net150),
    .A2(_08668_),
    .B1(_02869_),
    .Y(_00399_));
 sky130_fd_sc_hd__o21ai_1 _23618_ (.A1(net159),
    .A2(_08666_),
    .B1(_02858_),
    .Y(_00400_));
 sky130_fd_sc_hd__o22a_1 _23619_ (.A1(_00395_),
    .A2(_00396_),
    .B1(_00398_),
    .B2(_00399_),
    .X(_00401_));
 sky130_fd_sc_hd__o22ai_4 _23620_ (.A1(_00395_),
    .A2(_00396_),
    .B1(_00398_),
    .B2(_00399_),
    .Y(_00402_));
 sky130_fd_sc_hd__o211ai_4 _23621_ (.A1(net319),
    .A2(_02891_),
    .B1(_00397_),
    .C1(_00400_),
    .Y(_00403_));
 sky130_fd_sc_hd__o41a_1 _23622_ (.A1(_00395_),
    .A2(_00396_),
    .A3(_00398_),
    .A4(_00399_),
    .B1(_00393_),
    .X(_00404_));
 sky130_fd_sc_hd__a21oi_4 _23623_ (.A1(_00393_),
    .A2(_00403_),
    .B1(_00401_),
    .Y(_00406_));
 sky130_fd_sc_hd__a21oi_2 _23624_ (.A1(_00402_),
    .A2(_00403_),
    .B1(_00393_),
    .Y(_00407_));
 sky130_fd_sc_hd__a21o_1 _23625_ (.A1(_00402_),
    .A2(_00403_),
    .B1(_00393_),
    .X(_00408_));
 sky130_fd_sc_hd__o211a_1 _23626_ (.A1(_00391_),
    .A2(_00392_),
    .B1(_00402_),
    .C1(_00403_),
    .X(_00409_));
 sky130_fd_sc_hd__o211ai_4 _23627_ (.A1(_00391_),
    .A2(_00392_),
    .B1(_00402_),
    .C1(_00403_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _23628_ (.A(_00408_),
    .B(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__a22oi_1 _23629_ (.A1(_00035_),
    .A2(_00038_),
    .B1(_00408_),
    .B2(_00410_),
    .Y(_00412_));
 sky130_fd_sc_hd__o22ai_4 _23630_ (.A1(_00034_),
    .A2(_00037_),
    .B1(_00407_),
    .B2(_00409_),
    .Y(_00413_));
 sky130_fd_sc_hd__nor2_1 _23631_ (.A(_00039_),
    .B(_00407_),
    .Y(_00414_));
 sky130_fd_sc_hd__nor3_2 _23632_ (.A(_00039_),
    .B(_00407_),
    .C(_00409_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand3b_2 _23633_ (.A_N(_00039_),
    .B(_00408_),
    .C(_00410_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _23634_ (.A(_00413_),
    .B(_00417_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand4_2 _23635_ (.A(_00073_),
    .B(_00074_),
    .C(_00413_),
    .D(_00417_),
    .Y(_00419_));
 sky130_fd_sc_hd__o22ai_2 _23636_ (.A1(_00072_),
    .A2(_00075_),
    .B1(_00412_),
    .B2(_00415_),
    .Y(_00420_));
 sky130_fd_sc_hd__a21oi_2 _23637_ (.A1(_00413_),
    .A2(_00417_),
    .B1(_00390_),
    .Y(_00421_));
 sky130_fd_sc_hd__a221o_1 _23638_ (.A1(_00064_),
    .A2(_00071_),
    .B1(_00413_),
    .B2(_00417_),
    .C1(_00072_),
    .X(_00422_));
 sky130_fd_sc_hd__a21oi_2 _23639_ (.A1(_00411_),
    .A2(_00039_),
    .B1(_00389_),
    .Y(_00423_));
 sky130_fd_sc_hd__and3_1 _23640_ (.A(_00388_),
    .B(_00419_),
    .C(_00420_),
    .X(_00424_));
 sky130_fd_sc_hd__o211ai_4 _23641_ (.A1(_00080_),
    .A2(_00385_),
    .B1(_00419_),
    .C1(_00420_),
    .Y(_00425_));
 sky130_fd_sc_hd__and3_1 _23642_ (.A(_00081_),
    .B(_00386_),
    .C(_00422_),
    .X(_00426_));
 sky130_fd_sc_hd__o2bb2ai_2 _23643_ (.A1_N(_00389_),
    .A2_N(_00418_),
    .B1(_00083_),
    .B2(_00387_),
    .Y(_00428_));
 sky130_fd_sc_hd__a32o_1 _23644_ (.A1(_05933_),
    .A2(_05462_),
    .A3(net174),
    .B1(_05464_),
    .B2(net16),
    .X(_00429_));
 sky130_fd_sc_hd__a32oi_4 _23645_ (.A1(net202),
    .A2(net173),
    .A3(_05225_),
    .B1(_05228_),
    .B2(net17),
    .Y(_00430_));
 sky130_fd_sc_hd__o2111ai_2 _23646_ (.A1(net174),
    .A2(_06451_),
    .B1(net45),
    .C1(net197),
    .D1(_04102_),
    .Y(_00431_));
 sky130_fd_sc_hd__or3_1 _23647_ (.A(net45),
    .B(_04179_),
    .C(_04102_),
    .X(_00432_));
 sky130_fd_sc_hd__o221ai_4 _23648_ (.A1(_04179_),
    .A2(_04989_),
    .B1(_06454_),
    .B2(_04986_),
    .C1(_00430_),
    .Y(_00433_));
 sky130_fd_sc_hd__a21oi_2 _23649_ (.A1(_00431_),
    .A2(_00432_),
    .B1(_00430_),
    .Y(_00434_));
 sky130_fd_sc_hd__a21o_1 _23650_ (.A1(_00431_),
    .A2(_00432_),
    .B1(_00430_),
    .X(_00435_));
 sky130_fd_sc_hd__a21o_1 _23651_ (.A1(_00433_),
    .A2(_00435_),
    .B1(_00429_),
    .X(_00436_));
 sky130_fd_sc_hd__nand3_1 _23652_ (.A(_00429_),
    .B(_00433_),
    .C(_00435_),
    .Y(_00437_));
 sky130_fd_sc_hd__and2_1 _23653_ (.A(_00436_),
    .B(_00437_),
    .X(_00439_));
 sky130_fd_sc_hd__nand2_2 _23654_ (.A(_00436_),
    .B(_00437_),
    .Y(_00440_));
 sky130_fd_sc_hd__a21o_1 _23655_ (.A1(_00111_),
    .A2(_00118_),
    .B1(_00119_),
    .X(_00441_));
 sky130_fd_sc_hd__a32o_1 _23656_ (.A1(net194),
    .A2(net171),
    .A3(_04895_),
    .B1(_04897_),
    .B2(net19),
    .X(_00442_));
 sky130_fd_sc_hd__o211ai_4 _23657_ (.A1(net174),
    .A2(_07074_),
    .B1(_04480_),
    .C1(_07072_),
    .Y(_00443_));
 sky130_fd_sc_hd__or3b_2 _23658_ (.A(net42),
    .B(_04212_),
    .C_N(net41),
    .X(_00444_));
 sky130_fd_sc_hd__o211ai_4 _23659_ (.A1(net174),
    .A2(_07501_),
    .B1(_04267_),
    .C1(_07499_),
    .Y(_00445_));
 sky130_fd_sc_hd__or3b_1 _23660_ (.A(net41),
    .B(_04223_),
    .C_N(net40),
    .X(_00446_));
 sky130_fd_sc_hd__a22oi_2 _23661_ (.A1(_00443_),
    .A2(_00444_),
    .B1(_00445_),
    .B2(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__a22o_1 _23662_ (.A1(_00443_),
    .A2(_00444_),
    .B1(_00445_),
    .B2(_00446_),
    .X(_00448_));
 sky130_fd_sc_hd__o2111a_1 _23663_ (.A1(_04223_),
    .A2(_04270_),
    .B1(_00443_),
    .C1(_00444_),
    .D1(_00445_),
    .X(_00450_));
 sky130_fd_sc_hd__o2111ai_4 _23664_ (.A1(_04223_),
    .A2(_04270_),
    .B1(_00443_),
    .C1(_00444_),
    .D1(_00445_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand3_4 _23665_ (.A(_00442_),
    .B(_00448_),
    .C(_00451_),
    .Y(_00452_));
 sky130_fd_sc_hd__a21oi_1 _23666_ (.A1(_00448_),
    .A2(_00451_),
    .B1(_00442_),
    .Y(_00453_));
 sky130_fd_sc_hd__o21bai_2 _23667_ (.A1(_00447_),
    .A2(_00450_),
    .B1_N(_00442_),
    .Y(_00454_));
 sky130_fd_sc_hd__a21oi_2 _23668_ (.A1(_00120_),
    .A2(_00124_),
    .B1(_00453_),
    .Y(_00455_));
 sky130_fd_sc_hd__and3_1 _23669_ (.A(_00441_),
    .B(_00452_),
    .C(_00454_),
    .X(_00456_));
 sky130_fd_sc_hd__nand2_1 _23670_ (.A(_00455_),
    .B(_00452_),
    .Y(_00457_));
 sky130_fd_sc_hd__a21oi_2 _23671_ (.A1(_00452_),
    .A2(_00454_),
    .B1(_00441_),
    .Y(_00458_));
 sky130_fd_sc_hd__a21o_1 _23672_ (.A1(_00452_),
    .A2(_00454_),
    .B1(_00441_),
    .X(_00459_));
 sky130_fd_sc_hd__and3_1 _23673_ (.A(_00440_),
    .B(_00457_),
    .C(_00459_),
    .X(_00461_));
 sky130_fd_sc_hd__o211a_1 _23674_ (.A1(_00456_),
    .A2(_00458_),
    .B1(_00436_),
    .C1(_00437_),
    .X(_00462_));
 sky130_fd_sc_hd__nand2_1 _23675_ (.A(_00439_),
    .B(_00459_),
    .Y(_00463_));
 sky130_fd_sc_hd__a211oi_4 _23676_ (.A1(_00455_),
    .A2(_00452_),
    .B1(_00440_),
    .C1(_00458_),
    .Y(_00464_));
 sky130_fd_sc_hd__a21oi_2 _23677_ (.A1(_00457_),
    .A2(_00459_),
    .B1(_00439_),
    .Y(_00465_));
 sky130_fd_sc_hd__a22o_1 _23678_ (.A1(_00436_),
    .A2(_00437_),
    .B1(_00457_),
    .B2(_00459_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_1 _23679_ (.A(_00464_),
    .B(_00465_),
    .Y(_00467_));
 sky130_fd_sc_hd__o221ai_4 _23680_ (.A1(_00464_),
    .A2(_00465_),
    .B1(_00421_),
    .B2(_00388_),
    .C1(_00425_),
    .Y(_00468_));
 sky130_fd_sc_hd__o2bb2ai_1 _23681_ (.A1_N(_00425_),
    .A2_N(_00428_),
    .B1(_00461_),
    .B2(_00462_),
    .Y(_00469_));
 sky130_fd_sc_hd__o2bb2ai_2 _23682_ (.A1_N(_00425_),
    .A2_N(_00428_),
    .B1(_00464_),
    .B2(_00465_),
    .Y(_00470_));
 sky130_fd_sc_hd__o211a_1 _23683_ (.A1(_00456_),
    .A2(_00463_),
    .B1(_00466_),
    .C1(_00425_),
    .X(_00472_));
 sky130_fd_sc_hd__o2111ai_4 _23684_ (.A1(_00456_),
    .A2(_00463_),
    .B1(_00466_),
    .C1(_00428_),
    .D1(_00425_),
    .Y(_00473_));
 sky130_fd_sc_hd__a21oi_1 _23685_ (.A1(_00470_),
    .A2(_00473_),
    .B1(_00384_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand3_4 _23686_ (.A(_00383_),
    .B(_00468_),
    .C(_00469_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand3_4 _23687_ (.A(_00470_),
    .B(_00473_),
    .C(_00384_),
    .Y(_00476_));
 sky130_fd_sc_hd__o211a_1 _23688_ (.A1(_00127_),
    .A2(_00130_),
    .B1(_00133_),
    .C1(_00092_),
    .X(_00477_));
 sky130_fd_sc_hd__o21a_1 _23689_ (.A1(_00091_),
    .A2(_00135_),
    .B1(_00094_),
    .X(_00478_));
 sky130_fd_sc_hd__o211a_1 _23690_ (.A1(_00093_),
    .A2(_00477_),
    .B1(_00476_),
    .C1(_00475_),
    .X(_00479_));
 sky130_fd_sc_hd__o211ai_1 _23691_ (.A1(_00093_),
    .A2(_00477_),
    .B1(_00476_),
    .C1(_00475_),
    .Y(_00480_));
 sky130_fd_sc_hd__a211oi_1 _23692_ (.A1(_00475_),
    .A2(_00476_),
    .B1(_00477_),
    .C1(_00093_),
    .Y(_00481_));
 sky130_fd_sc_hd__a21bo_1 _23693_ (.A1(_00475_),
    .A2(_00476_),
    .B1_N(_00478_),
    .X(_00483_));
 sky130_fd_sc_hd__a21oi_1 _23694_ (.A1(_00475_),
    .A2(_00476_),
    .B1(_00478_),
    .Y(_00484_));
 sky130_fd_sc_hd__a21o_1 _23695_ (.A1(_00475_),
    .A2(_00476_),
    .B1(_00478_),
    .X(_00485_));
 sky130_fd_sc_hd__and3_1 _23696_ (.A(_00475_),
    .B(_00476_),
    .C(_00478_),
    .X(_00486_));
 sky130_fd_sc_hd__o2111ai_4 _23697_ (.A1(_00091_),
    .A2(_00135_),
    .B1(_00475_),
    .C1(_00476_),
    .D1(_00094_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand4_2 _23698_ (.A(_00381_),
    .B(_00382_),
    .C(_00485_),
    .D(_00487_),
    .Y(_00488_));
 sky130_fd_sc_hd__o2bb2ai_2 _23699_ (.A1_N(_00381_),
    .A2_N(_00382_),
    .B1(_00484_),
    .B2(_00486_),
    .Y(_00489_));
 sky130_fd_sc_hd__o2bb2ai_1 _23700_ (.A1_N(_00381_),
    .A2_N(_00382_),
    .B1(_00479_),
    .B2(_00481_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand4_2 _23701_ (.A(_00381_),
    .B(_00382_),
    .C(_00480_),
    .D(_00483_),
    .Y(_00491_));
 sky130_fd_sc_hd__o2111a_1 _23702_ (.A1(_00060_),
    .A2(_00058_),
    .B1(_00488_),
    .C1(_00152_),
    .D1(_00489_),
    .X(_00492_));
 sky130_fd_sc_hd__o2111ai_4 _23703_ (.A1(_00060_),
    .A2(_00058_),
    .B1(_00488_),
    .C1(_00152_),
    .D1(_00489_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand4_4 _23704_ (.A(_00062_),
    .B(_00316_),
    .C(_00490_),
    .D(_00491_),
    .Y(_00495_));
 sky130_fd_sc_hd__a21boi_4 _23705_ (.A1(_00210_),
    .A2(_00254_),
    .B1_N(_00211_),
    .Y(_00496_));
 sky130_fd_sc_hd__a31oi_2 _23706_ (.A1(_00136_),
    .A2(_00137_),
    .A3(_00139_),
    .B1(_00146_),
    .Y(_00497_));
 sky130_fd_sc_hd__a31o_2 _23707_ (.A1(_00136_),
    .A2(_00137_),
    .A3(_00139_),
    .B1(_00146_),
    .X(_00498_));
 sky130_fd_sc_hd__a21oi_1 _23708_ (.A1(_00141_),
    .A2(_00146_),
    .B1(_00142_),
    .Y(_00499_));
 sky130_fd_sc_hd__nor2_1 _23709_ (.A(_00163_),
    .B(_00201_),
    .Y(_00500_));
 sky130_fd_sc_hd__a21o_1 _23710_ (.A1(_00163_),
    .A2(_00204_),
    .B1(_00201_),
    .X(_00501_));
 sky130_fd_sc_hd__a2bb2o_1 _23711_ (.A1_N(_00191_),
    .A2_N(_00186_),
    .B1(_00167_),
    .B2(_00194_),
    .X(_00502_));
 sky130_fd_sc_hd__o2bb2ai_1 _23712_ (.A1_N(_00106_),
    .A2_N(_00129_),
    .B1(_00126_),
    .B2(_00123_),
    .Y(_00503_));
 sky130_fd_sc_hd__a21oi_1 _23713_ (.A1(_00106_),
    .A2(_00129_),
    .B1(_00127_),
    .Y(_00505_));
 sky130_fd_sc_hd__a21o_1 _23714_ (.A1(_00173_),
    .A2(_00182_),
    .B1(_00183_),
    .X(_00506_));
 sky130_fd_sc_hd__a32o_1 _23715_ (.A1(net209),
    .A2(_05074_),
    .A3(net273),
    .B1(_06326_),
    .B2(net13),
    .X(_00507_));
 sky130_fd_sc_hd__nor2_1 _23716_ (.A(_04146_),
    .B(_05766_),
    .Y(_00508_));
 sky130_fd_sc_hd__a211oi_2 _23717_ (.A1(_04788_),
    .A2(_05550_),
    .B1(_05763_),
    .C1(_05548_),
    .Y(_00509_));
 sky130_fd_sc_hd__o211ai_1 _23718_ (.A1(net184),
    .A2(_05551_),
    .B1(_05762_),
    .C1(net178),
    .Y(_00510_));
 sky130_fd_sc_hd__nand3_1 _23719_ (.A(_05290_),
    .B(_05292_),
    .C(net274),
    .Y(_00511_));
 sky130_fd_sc_hd__or3b_1 _23720_ (.A(_04135_),
    .B(net49),
    .C_N(net48),
    .X(_00512_));
 sky130_fd_sc_hd__o21ai_1 _23721_ (.A1(_04135_),
    .A2(_06030_),
    .B1(_00511_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand3_1 _23722_ (.A(_00510_),
    .B(_00511_),
    .C(_00512_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand4b_1 _23723_ (.A_N(_00508_),
    .B(_00510_),
    .C(_00511_),
    .D(_00512_),
    .Y(_00516_));
 sky130_fd_sc_hd__o21ai_2 _23724_ (.A1(_00508_),
    .A2(_00509_),
    .B1(_00513_),
    .Y(_00517_));
 sky130_fd_sc_hd__inv_2 _23725_ (.A(_00517_),
    .Y(_00518_));
 sky130_fd_sc_hd__o211a_2 _23726_ (.A1(_00514_),
    .A2(_00508_),
    .B1(_00507_),
    .C1(_00517_),
    .X(_00519_));
 sky130_fd_sc_hd__o211ai_2 _23727_ (.A1(_00514_),
    .A2(_00508_),
    .B1(_00507_),
    .C1(_00517_),
    .Y(_00520_));
 sky130_fd_sc_hd__a21oi_1 _23728_ (.A1(_00516_),
    .A2(_00517_),
    .B1(_00507_),
    .Y(_00521_));
 sky130_fd_sc_hd__a21o_1 _23729_ (.A1(_00516_),
    .A2(_00517_),
    .B1(_00507_),
    .X(_00522_));
 sky130_fd_sc_hd__and3_1 _23730_ (.A(_00522_),
    .B(_00104_),
    .C(_00520_),
    .X(_00523_));
 sky130_fd_sc_hd__nand3_1 _23731_ (.A(_00522_),
    .B(_00104_),
    .C(_00520_),
    .Y(_00524_));
 sky130_fd_sc_hd__o22ai_4 _23732_ (.A1(_00100_),
    .A2(_00103_),
    .B1(_00519_),
    .B2(_00521_),
    .Y(_00525_));
 sky130_fd_sc_hd__a22o_1 _23733_ (.A1(_00184_),
    .A2(_00188_),
    .B1(_00524_),
    .B2(_00525_),
    .X(_00527_));
 sky130_fd_sc_hd__o2111ai_1 _23734_ (.A1(_00185_),
    .A2(_00172_),
    .B1(_00184_),
    .C1(_00524_),
    .D1(_00525_),
    .Y(_00528_));
 sky130_fd_sc_hd__o21a_2 _23735_ (.A1(_00183_),
    .A2(_00186_),
    .B1(_00525_),
    .X(_00529_));
 sky130_fd_sc_hd__o211ai_1 _23736_ (.A1(_00183_),
    .A2(_00186_),
    .B1(_00524_),
    .C1(_00525_),
    .Y(_00530_));
 sky130_fd_sc_hd__a21o_1 _23737_ (.A1(_00524_),
    .A2(_00525_),
    .B1(_00506_),
    .X(_00531_));
 sky130_fd_sc_hd__and3_2 _23738_ (.A(_00531_),
    .B(_00503_),
    .C(_00530_),
    .X(_00532_));
 sky130_fd_sc_hd__nand3_2 _23739_ (.A(_00531_),
    .B(_00503_),
    .C(_00530_),
    .Y(_00533_));
 sky130_fd_sc_hd__nand3_2 _23740_ (.A(_00505_),
    .B(_00527_),
    .C(_00528_),
    .Y(_00534_));
 sky130_fd_sc_hd__o211a_2 _23741_ (.A1(_00192_),
    .A2(_00196_),
    .B1(_00533_),
    .C1(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__o211ai_2 _23742_ (.A1(_00192_),
    .A2(_00196_),
    .B1(_00533_),
    .C1(_00534_),
    .Y(_00536_));
 sky130_fd_sc_hd__a21oi_1 _23743_ (.A1(_00533_),
    .A2(_00534_),
    .B1(_00502_),
    .Y(_00538_));
 sky130_fd_sc_hd__a21o_1 _23744_ (.A1(_00533_),
    .A2(_00534_),
    .B1(_00502_),
    .X(_00539_));
 sky130_fd_sc_hd__nand3_4 _23745_ (.A(_00539_),
    .B(_00501_),
    .C(_00536_),
    .Y(_00540_));
 sky130_fd_sc_hd__o22ai_4 _23746_ (.A1(_00203_),
    .A2(_00500_),
    .B1(_00535_),
    .B2(_00538_),
    .Y(_00541_));
 sky130_fd_sc_hd__or4_2 _23747_ (.A(net54),
    .B(_04266_),
    .C(_03951_),
    .D(_03957_),
    .X(_00542_));
 sky130_fd_sc_hd__o2bb2a_2 _23748_ (.A1_N(_03959_),
    .A2_N(net238),
    .B1(_08007_),
    .B2(_04048_),
    .X(_00543_));
 sky130_fd_sc_hd__a21boi_2 _23749_ (.A1(_00218_),
    .A2(_00237_),
    .B1_N(_00236_),
    .Y(_00544_));
 sky130_fd_sc_hd__a32oi_2 _23750_ (.A1(net229),
    .A2(net227),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net8),
    .Y(_00545_));
 sky130_fd_sc_hd__a32o_1 _23751_ (.A1(net229),
    .A2(net227),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net8),
    .X(_00546_));
 sky130_fd_sc_hd__or3b_1 _23752_ (.A(_04080_),
    .B(net52),
    .C_N(net51),
    .X(_00547_));
 sky130_fd_sc_hd__o211ai_2 _23753_ (.A1(net233),
    .A2(_04557_),
    .B1(net269),
    .C1(net217),
    .Y(_00549_));
 sky130_fd_sc_hd__nor2_1 _23754_ (.A(_04091_),
    .B(_06866_),
    .Y(_00550_));
 sky130_fd_sc_hd__o311a_1 _23755_ (.A1(net7),
    .A2(net248),
    .A3(_04787_),
    .B1(net240),
    .C1(net213),
    .X(_00551_));
 sky130_fd_sc_hd__a31oi_1 _23756_ (.A1(net184),
    .A2(net213),
    .A3(net240),
    .B1(_00550_),
    .Y(_00552_));
 sky130_fd_sc_hd__o211ai_2 _23757_ (.A1(_04080_),
    .A2(_07226_),
    .B1(_00549_),
    .C1(_00552_),
    .Y(_00553_));
 sky130_fd_sc_hd__o2bb2ai_1 _23758_ (.A1_N(_00547_),
    .A2_N(_00549_),
    .B1(_00550_),
    .B2(_00551_),
    .Y(_00554_));
 sky130_fd_sc_hd__a32o_1 _23759_ (.A1(_04409_),
    .A2(net225),
    .A3(net239),
    .B1(_07308_),
    .B2(net9),
    .X(_00555_));
 sky130_fd_sc_hd__a21o_1 _23760_ (.A1(_00553_),
    .A2(_00554_),
    .B1(_00555_),
    .X(_00556_));
 sky130_fd_sc_hd__nand3_2 _23761_ (.A(_00553_),
    .B(_00554_),
    .C(_00555_),
    .Y(_00557_));
 sky130_fd_sc_hd__o21ai_2 _23762_ (.A1(_00221_),
    .A2(_00229_),
    .B1(_00228_),
    .Y(_00558_));
 sky130_fd_sc_hd__a21oi_1 _23763_ (.A1(_00556_),
    .A2(_00557_),
    .B1(_00558_),
    .Y(_00560_));
 sky130_fd_sc_hd__a21o_1 _23764_ (.A1(_00556_),
    .A2(_00557_),
    .B1(_00558_),
    .X(_00561_));
 sky130_fd_sc_hd__and3_1 _23765_ (.A(_00556_),
    .B(_00558_),
    .C(_00557_),
    .X(_00562_));
 sky130_fd_sc_hd__nand3_1 _23766_ (.A(_00556_),
    .B(_00557_),
    .C(_00558_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand3_1 _23767_ (.A(_00546_),
    .B(_00561_),
    .C(_00563_),
    .Y(_00564_));
 sky130_fd_sc_hd__o21ai_1 _23768_ (.A1(_00560_),
    .A2(_00562_),
    .B1(_00545_),
    .Y(_00565_));
 sky130_fd_sc_hd__o21ai_1 _23769_ (.A1(_00560_),
    .A2(_00562_),
    .B1(_00546_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand3_1 _23770_ (.A(_00561_),
    .B(_00563_),
    .C(_00545_),
    .Y(_00567_));
 sky130_fd_sc_hd__a21oi_2 _23771_ (.A1(_00566_),
    .A2(_00567_),
    .B1(_00544_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand3b_2 _23772_ (.A_N(_00544_),
    .B(_00564_),
    .C(_00565_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand3_2 _23773_ (.A(_00544_),
    .B(_00566_),
    .C(_00567_),
    .Y(_00571_));
 sky130_fd_sc_hd__inv_2 _23774_ (.A(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _23775_ (.A(_00569_),
    .B(_00571_),
    .Y(_00573_));
 sky130_fd_sc_hd__a21oi_2 _23776_ (.A1(_00569_),
    .A2(_00571_),
    .B1(_00543_),
    .Y(_00574_));
 sky130_fd_sc_hd__and3_1 _23777_ (.A(_00569_),
    .B(_00571_),
    .C(_00543_),
    .X(_00575_));
 sky130_fd_sc_hd__o211a_1 _23778_ (.A1(_04048_),
    .A2(_08007_),
    .B1(_00542_),
    .C1(_00573_),
    .X(_00576_));
 sky130_fd_sc_hd__nor2_2 _23779_ (.A(_00543_),
    .B(_00573_),
    .Y(_00577_));
 sky130_fd_sc_hd__nor2_1 _23780_ (.A(_00574_),
    .B(_00575_),
    .Y(_00578_));
 sky130_fd_sc_hd__o21a_1 _23781_ (.A1(_00574_),
    .A2(_00575_),
    .B1(_00541_),
    .X(_00579_));
 sky130_fd_sc_hd__o211a_1 _23782_ (.A1(_00574_),
    .A2(_00575_),
    .B1(_00540_),
    .C1(_00541_),
    .X(_00580_));
 sky130_fd_sc_hd__o211ai_4 _23783_ (.A1(_00574_),
    .A2(_00575_),
    .B1(_00540_),
    .C1(_00541_),
    .Y(_00582_));
 sky130_fd_sc_hd__a21boi_1 _23784_ (.A1(_00540_),
    .A2(_00541_),
    .B1_N(_00578_),
    .Y(_00583_));
 sky130_fd_sc_hd__o2bb2ai_4 _23785_ (.A1_N(_00540_),
    .A2_N(_00541_),
    .B1(_00576_),
    .B2(_00577_),
    .Y(_00584_));
 sky130_fd_sc_hd__a31o_2 _23786_ (.A1(_00501_),
    .A2(_00536_),
    .A3(_00539_),
    .B1(_00579_),
    .X(_00585_));
 sky130_fd_sc_hd__nand3_2 _23787_ (.A(_00141_),
    .B(_00498_),
    .C(_00584_),
    .Y(_00586_));
 sky130_fd_sc_hd__and4_1 _23788_ (.A(_00141_),
    .B(_00498_),
    .C(_00582_),
    .D(_00584_),
    .X(_00587_));
 sky130_fd_sc_hd__nand4_4 _23789_ (.A(_00141_),
    .B(_00498_),
    .C(_00582_),
    .D(_00584_),
    .Y(_00588_));
 sky130_fd_sc_hd__a2bb2oi_4 _23790_ (.A1_N(_00140_),
    .A2_N(_00497_),
    .B1(_00582_),
    .B2(_00584_),
    .Y(_00589_));
 sky130_fd_sc_hd__a22o_1 _23791_ (.A1(_00141_),
    .A2(_00498_),
    .B1(_00582_),
    .B2(_00584_),
    .X(_00590_));
 sky130_fd_sc_hd__a21oi_1 _23792_ (.A1(_00211_),
    .A2(_00258_),
    .B1(_00589_),
    .Y(_00591_));
 sky130_fd_sc_hd__nor3b_1 _23793_ (.A(_00589_),
    .B(_00496_),
    .C_N(_00588_),
    .Y(_00593_));
 sky130_fd_sc_hd__a21boi_1 _23794_ (.A1(_00588_),
    .A2(_00590_),
    .B1_N(_00496_),
    .Y(_00594_));
 sky130_fd_sc_hd__a21oi_1 _23795_ (.A1(_00211_),
    .A2(_00258_),
    .B1(_00588_),
    .Y(_00595_));
 sky130_fd_sc_hd__a211o_1 _23796_ (.A1(_00579_),
    .A2(_00540_),
    .B1(_00496_),
    .C1(_00586_),
    .X(_00596_));
 sky130_fd_sc_hd__o211ai_2 _23797_ (.A1(_00580_),
    .A2(_00583_),
    .B1(_00496_),
    .C1(_00499_),
    .Y(_00597_));
 sky130_fd_sc_hd__and3_1 _23798_ (.A(_00211_),
    .B(_00258_),
    .C(_00588_),
    .X(_00598_));
 sky130_fd_sc_hd__a31o_1 _23799_ (.A1(_00211_),
    .A2(_00258_),
    .A3(_00588_),
    .B1(_00589_),
    .X(_00599_));
 sky130_fd_sc_hd__inv_2 _23800_ (.A(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__o221a_1 _23801_ (.A1(_00580_),
    .A2(_00586_),
    .B1(_00496_),
    .B2(_00589_),
    .C1(_00597_),
    .X(_00601_));
 sky130_fd_sc_hd__o221ai_4 _23802_ (.A1(_00580_),
    .A2(_00586_),
    .B1(_00496_),
    .B2(_00589_),
    .C1(_00597_),
    .Y(_00602_));
 sky130_fd_sc_hd__o21ai_1 _23803_ (.A1(_00496_),
    .A2(_00588_),
    .B1(_00602_),
    .Y(_00604_));
 sky130_fd_sc_hd__o2111ai_2 _23804_ (.A1(_00496_),
    .A2(_00588_),
    .B1(_00602_),
    .C1(_00495_),
    .D1(_00494_),
    .Y(_00605_));
 sky130_fd_sc_hd__o2bb2ai_1 _23805_ (.A1_N(_00494_),
    .A2_N(_00495_),
    .B1(_00595_),
    .B2(_00601_),
    .Y(_00606_));
 sky130_fd_sc_hd__o2bb2ai_1 _23806_ (.A1_N(_00494_),
    .A2_N(_00495_),
    .B1(_00593_),
    .B2(_00594_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand3_1 _23807_ (.A(_00604_),
    .B(_00495_),
    .C(_00494_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand3_2 _23808_ (.A(_00315_),
    .B(_00605_),
    .C(_00606_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand3_4 _23809_ (.A(_00314_),
    .B(_00607_),
    .C(_00608_),
    .Y(_00610_));
 sky130_fd_sc_hd__and3_1 _23810_ (.A(_13286_),
    .B(_13315_),
    .C(_00265_),
    .X(_00611_));
 sky130_fd_sc_hd__o2bb2ai_2 _23811_ (.A1_N(_00609_),
    .A2_N(_00610_),
    .B1(_00611_),
    .B2(_00261_),
    .Y(_00612_));
 sky130_fd_sc_hd__o211ai_4 _23812_ (.A1(_00263_),
    .A2(_00269_),
    .B1(_00609_),
    .C1(_00610_),
    .Y(_00613_));
 sky130_fd_sc_hd__o21ai_1 _23813_ (.A1(_13369_),
    .A2(_00277_),
    .B1(_00280_),
    .Y(_00615_));
 sky130_fd_sc_hd__a21oi_2 _23814_ (.A1(_00612_),
    .A2(_00613_),
    .B1(_00615_),
    .Y(_00616_));
 sky130_fd_sc_hd__a21o_1 _23815_ (.A1(_00612_),
    .A2(_00613_),
    .B1(_00615_),
    .X(_00617_));
 sky130_fd_sc_hd__o211a_2 _23816_ (.A1(_00279_),
    .A2(_00282_),
    .B1(_00612_),
    .C1(_00613_),
    .X(_00618_));
 sky130_fd_sc_hd__o211ai_1 _23817_ (.A1(_00279_),
    .A2(_00282_),
    .B1(_00612_),
    .C1(_00613_),
    .Y(_00619_));
 sky130_fd_sc_hd__o22ai_1 _23818_ (.A1(_00243_),
    .A2(_00312_),
    .B1(_00616_),
    .B2(_00618_),
    .Y(_00620_));
 sky130_fd_sc_hd__o211ai_1 _23819_ (.A1(_00245_),
    .A2(_00311_),
    .B1(_00617_),
    .C1(_00619_),
    .Y(_00621_));
 sky130_fd_sc_hd__o211a_1 _23820_ (.A1(_00214_),
    .A2(_00245_),
    .B1(_00619_),
    .C1(_00244_),
    .X(_00622_));
 sky130_fd_sc_hd__nor2_1 _23821_ (.A(_00313_),
    .B(_00616_),
    .Y(_00623_));
 sky130_fd_sc_hd__o21ai_1 _23822_ (.A1(_00243_),
    .A2(_00312_),
    .B1(_00617_),
    .Y(_00624_));
 sky130_fd_sc_hd__o21ai_1 _23823_ (.A1(_00616_),
    .A2(_00618_),
    .B1(_00313_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand3_1 _23824_ (.A(_00310_),
    .B(_00620_),
    .C(_00621_),
    .Y(_00627_));
 sky130_fd_sc_hd__o221ai_4 _23825_ (.A1(_00289_),
    .A2(_00293_),
    .B1(_00618_),
    .B2(_00624_),
    .C1(_00626_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _23826_ (.A(_00627_),
    .B(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__o21a_1 _23827_ (.A1(_00299_),
    .A2(_00309_),
    .B1(_00298_),
    .X(_00630_));
 sky130_fd_sc_hd__xnor2_1 _23828_ (.A(_00629_),
    .B(_00630_),
    .Y(net104));
 sky130_fd_sc_hd__o211a_1 _23829_ (.A1(_04048_),
    .A2(_08007_),
    .B1(_00542_),
    .C1(_00569_),
    .X(_00631_));
 sky130_fd_sc_hd__o21a_1 _23830_ (.A1(_00543_),
    .A2(_00573_),
    .B1(_00569_),
    .X(_00632_));
 sky130_fd_sc_hd__o211ai_4 _23831_ (.A1(_00496_),
    .A2(_00588_),
    .B1(_00602_),
    .C1(_00495_),
    .Y(_00633_));
 sky130_fd_sc_hd__a31o_1 _23832_ (.A1(_00495_),
    .A2(_00596_),
    .A3(_00602_),
    .B1(_00492_),
    .X(_00634_));
 sky130_fd_sc_hd__a31oi_1 _23833_ (.A1(_00495_),
    .A2(_00596_),
    .A3(_00602_),
    .B1(_00492_),
    .Y(_00636_));
 sky130_fd_sc_hd__a21oi_1 _23834_ (.A1(_00502_),
    .A2(_00534_),
    .B1(_00532_),
    .Y(_00637_));
 sky130_fd_sc_hd__a21o_1 _23835_ (.A1(_00502_),
    .A2(_00534_),
    .B1(_00532_),
    .X(_00638_));
 sky130_fd_sc_hd__a21o_1 _23836_ (.A1(_00507_),
    .A2(_00516_),
    .B1(_00518_),
    .X(_00639_));
 sky130_fd_sc_hd__a221oi_4 _23837_ (.A1(_03957_),
    .A2(_05926_),
    .B1(_05553_),
    .B2(net16),
    .C1(_05763_),
    .Y(_00640_));
 sky130_fd_sc_hd__a221o_1 _23838_ (.A1(_03957_),
    .A2(_05926_),
    .B1(_05553_),
    .B2(net16),
    .C1(_05763_),
    .X(_00641_));
 sky130_fd_sc_hd__nor2_1 _23839_ (.A(_04157_),
    .B(_05766_),
    .Y(_00642_));
 sky130_fd_sc_hd__or3b_1 _23840_ (.A(net48),
    .B(_04157_),
    .C_N(net47),
    .X(_00643_));
 sky130_fd_sc_hd__o211ai_1 _23841_ (.A1(net184),
    .A2(_05551_),
    .B1(net274),
    .C1(net178),
    .Y(_00644_));
 sky130_fd_sc_hd__nor2_1 _23842_ (.A(_04146_),
    .B(_06030_),
    .Y(_00645_));
 sky130_fd_sc_hd__or3b_1 _23843_ (.A(_04146_),
    .B(net49),
    .C_N(net48),
    .X(_00647_));
 sky130_fd_sc_hd__a31o_1 _23844_ (.A1(net178),
    .A2(_05553_),
    .A3(net274),
    .B1(_00645_),
    .X(_00648_));
 sky130_fd_sc_hd__o21a_1 _23845_ (.A1(_00640_),
    .A2(_00642_),
    .B1(_00648_),
    .X(_00649_));
 sky130_fd_sc_hd__o21ai_2 _23846_ (.A1(_00640_),
    .A2(_00642_),
    .B1(_00648_),
    .Y(_00650_));
 sky130_fd_sc_hd__a31o_1 _23847_ (.A1(net178),
    .A2(_05553_),
    .A3(net274),
    .B1(_00642_),
    .X(_00651_));
 sky130_fd_sc_hd__nand4_2 _23848_ (.A(_00641_),
    .B(_00643_),
    .C(_00644_),
    .D(_00647_),
    .Y(_00652_));
 sky130_fd_sc_hd__a32o_1 _23849_ (.A1(_05290_),
    .A2(_05292_),
    .A3(net273),
    .B1(_06326_),
    .B2(net14),
    .X(_00653_));
 sky130_fd_sc_hd__a21oi_2 _23850_ (.A1(_00650_),
    .A2(_00652_),
    .B1(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__a21o_1 _23851_ (.A1(_00650_),
    .A2(_00652_),
    .B1(_00653_),
    .X(_00655_));
 sky130_fd_sc_hd__o311a_2 _23852_ (.A1(_00640_),
    .A2(_00645_),
    .A3(_00651_),
    .B1(_00653_),
    .C1(_00650_),
    .X(_00656_));
 sky130_fd_sc_hd__nand3_1 _23853_ (.A(_00650_),
    .B(_00652_),
    .C(_00653_),
    .Y(_00658_));
 sky130_fd_sc_hd__a21o_1 _23854_ (.A1(_00429_),
    .A2(_00433_),
    .B1(_00434_),
    .X(_00659_));
 sky130_fd_sc_hd__a21oi_4 _23855_ (.A1(_00429_),
    .A2(_00433_),
    .B1(_00434_),
    .Y(_00660_));
 sky130_fd_sc_hd__o21ai_4 _23856_ (.A1(_00654_),
    .A2(_00656_),
    .B1(_00660_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand3_4 _23857_ (.A(_00655_),
    .B(_00659_),
    .C(_00658_),
    .Y(_00662_));
 sky130_fd_sc_hd__a21oi_1 _23858_ (.A1(_00661_),
    .A2(_00662_),
    .B1(_00639_),
    .Y(_00663_));
 sky130_fd_sc_hd__a21o_1 _23859_ (.A1(_00661_),
    .A2(_00662_),
    .B1(_00639_),
    .X(_00664_));
 sky130_fd_sc_hd__o21ai_2 _23860_ (.A1(_00518_),
    .A2(_00519_),
    .B1(_00661_),
    .Y(_00665_));
 sky130_fd_sc_hd__o211a_1 _23861_ (.A1(_00518_),
    .A2(_00519_),
    .B1(_00661_),
    .C1(_00662_),
    .X(_00666_));
 sky130_fd_sc_hd__o211ai_2 _23862_ (.A1(_00518_),
    .A2(_00519_),
    .B1(_00661_),
    .C1(_00662_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _23863_ (.A(_00664_),
    .B(_00667_),
    .Y(_00669_));
 sky130_fd_sc_hd__o2bb2ai_2 _23864_ (.A1_N(_00452_),
    .A2_N(_00455_),
    .B1(_00440_),
    .B2(_00458_),
    .Y(_00670_));
 sky130_fd_sc_hd__o2bb2a_1 _23865_ (.A1_N(_00452_),
    .A2_N(_00455_),
    .B1(_00440_),
    .B2(_00458_),
    .X(_00671_));
 sky130_fd_sc_hd__o21bai_4 _23866_ (.A1(_00663_),
    .A2(_00666_),
    .B1_N(_00670_),
    .Y(_00672_));
 sky130_fd_sc_hd__and3_1 _23867_ (.A(_00664_),
    .B(_00667_),
    .C(_00670_),
    .X(_00673_));
 sky130_fd_sc_hd__nand3_2 _23868_ (.A(_00664_),
    .B(_00667_),
    .C(_00670_),
    .Y(_00674_));
 sky130_fd_sc_hd__a31o_1 _23869_ (.A1(_00104_),
    .A2(_00520_),
    .A3(_00522_),
    .B1(_00529_),
    .X(_00675_));
 sky130_fd_sc_hd__a21oi_1 _23870_ (.A1(_00672_),
    .A2(_00674_),
    .B1(_00675_),
    .Y(_00676_));
 sky130_fd_sc_hd__a21o_1 _23871_ (.A1(_00672_),
    .A2(_00674_),
    .B1(_00675_),
    .X(_00677_));
 sky130_fd_sc_hd__a2bb2oi_2 _23872_ (.A1_N(_00523_),
    .A2_N(_00529_),
    .B1(_00669_),
    .B2(_00671_),
    .Y(_00678_));
 sky130_fd_sc_hd__o211a_1 _23873_ (.A1(_00523_),
    .A2(_00529_),
    .B1(_00672_),
    .C1(_00674_),
    .X(_00680_));
 sky130_fd_sc_hd__o211ai_4 _23874_ (.A1(_00523_),
    .A2(_00529_),
    .B1(_00672_),
    .C1(_00674_),
    .Y(_00681_));
 sky130_fd_sc_hd__a21oi_1 _23875_ (.A1(_00677_),
    .A2(_00681_),
    .B1(_00638_),
    .Y(_00682_));
 sky130_fd_sc_hd__o21ai_2 _23876_ (.A1(_00676_),
    .A2(_00680_),
    .B1(_00637_),
    .Y(_00683_));
 sky130_fd_sc_hd__o211a_1 _23877_ (.A1(_00532_),
    .A2(_00535_),
    .B1(_00677_),
    .C1(_00681_),
    .X(_00684_));
 sky130_fd_sc_hd__o211ai_4 _23878_ (.A1(_00532_),
    .A2(_00535_),
    .B1(_00677_),
    .C1(_00681_),
    .Y(_00685_));
 sky130_fd_sc_hd__a32o_1 _23879_ (.A1(_04409_),
    .A2(net225),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net9),
    .X(_00686_));
 sky130_fd_sc_hd__a21boi_2 _23880_ (.A1(_00553_),
    .A2(_00555_),
    .B1_N(_00554_),
    .Y(_00687_));
 sky130_fd_sc_hd__a32oi_4 _23881_ (.A1(net220),
    .A2(net186),
    .A3(net239),
    .B1(_07308_),
    .B2(net10),
    .Y(_00688_));
 sky130_fd_sc_hd__a32o_1 _23882_ (.A1(net220),
    .A2(net186),
    .A3(net239),
    .B1(_07308_),
    .B2(net10),
    .X(_00689_));
 sky130_fd_sc_hd__nor2_1 _23883_ (.A(_04113_),
    .B(_06866_),
    .Y(_00691_));
 sky130_fd_sc_hd__a31oi_4 _23884_ (.A1(net209),
    .A2(_05074_),
    .A3(net240),
    .B1(_00691_),
    .Y(_00692_));
 sky130_fd_sc_hd__or3b_1 _23885_ (.A(_04091_),
    .B(net52),
    .C_N(net51),
    .X(_00693_));
 sky130_fd_sc_hd__o221ai_4 _23886_ (.A1(net233),
    .A2(_04787_),
    .B1(_04091_),
    .B2(net216),
    .C1(net269),
    .Y(_00694_));
 sky130_fd_sc_hd__o211ai_4 _23887_ (.A1(_04091_),
    .A2(_07226_),
    .B1(_00694_),
    .C1(_00692_),
    .Y(_00695_));
 sky130_fd_sc_hd__a21oi_1 _23888_ (.A1(_00693_),
    .A2(_00694_),
    .B1(_00692_),
    .Y(_00696_));
 sky130_fd_sc_hd__a21o_1 _23889_ (.A1(_00693_),
    .A2(_00694_),
    .B1(_00692_),
    .X(_00697_));
 sky130_fd_sc_hd__nand3_1 _23890_ (.A(_00689_),
    .B(_00695_),
    .C(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__a21o_1 _23891_ (.A1(_00695_),
    .A2(_00697_),
    .B1(_00689_),
    .X(_00699_));
 sky130_fd_sc_hd__nand3_1 _23892_ (.A(_00697_),
    .B(_00688_),
    .C(_00695_),
    .Y(_00700_));
 sky130_fd_sc_hd__a21o_1 _23893_ (.A1(_00695_),
    .A2(_00697_),
    .B1(_00688_),
    .X(_00702_));
 sky130_fd_sc_hd__nand3b_4 _23894_ (.A_N(_00687_),
    .B(_00698_),
    .C(_00699_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand3_2 _23895_ (.A(_00702_),
    .B(_00687_),
    .C(_00700_),
    .Y(_00704_));
 sky130_fd_sc_hd__a21o_1 _23896_ (.A1(_00703_),
    .A2(_00704_),
    .B1(_00686_),
    .X(_00705_));
 sky130_fd_sc_hd__nand3_4 _23897_ (.A(_00686_),
    .B(_00703_),
    .C(_00704_),
    .Y(_00706_));
 sky130_fd_sc_hd__nor2_1 _23898_ (.A(_00545_),
    .B(_00560_),
    .Y(_00707_));
 sky130_fd_sc_hd__a32o_1 _23899_ (.A1(_00556_),
    .A2(_00557_),
    .A3(_00558_),
    .B1(_00561_),
    .B2(_00546_),
    .X(_00708_));
 sky130_fd_sc_hd__a21oi_2 _23900_ (.A1(_00705_),
    .A2(_00706_),
    .B1(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__o211a_2 _23901_ (.A1(_00562_),
    .A2(_00707_),
    .B1(_00706_),
    .C1(_00705_),
    .X(_00710_));
 sky130_fd_sc_hd__a32o_1 _23902_ (.A1(net229),
    .A2(net227),
    .A3(net238),
    .B1(_08006_),
    .B2(net8),
    .X(_00711_));
 sky130_fd_sc_hd__o21ba_1 _23903_ (.A1(_00709_),
    .A2(_00710_),
    .B1_N(_00711_),
    .X(_00713_));
 sky130_fd_sc_hd__nor3b_4 _23904_ (.A(_00709_),
    .B(_00710_),
    .C_N(_00711_),
    .Y(_00714_));
 sky130_fd_sc_hd__nor2_1 _23905_ (.A(_00713_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__a21oi_2 _23906_ (.A1(_00683_),
    .A2(_00685_),
    .B1(_00715_),
    .Y(_00716_));
 sky130_fd_sc_hd__o2bb2ai_1 _23907_ (.A1_N(_00683_),
    .A2_N(_00685_),
    .B1(_00713_),
    .B2(_00714_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand3_1 _23908_ (.A(_00715_),
    .B(_00685_),
    .C(_00683_),
    .Y(_00718_));
 sky130_fd_sc_hd__o21ai_1 _23909_ (.A1(_00682_),
    .A2(_00684_),
    .B1(_00715_),
    .Y(_00719_));
 sky130_fd_sc_hd__o211ai_2 _23910_ (.A1(_00713_),
    .A2(_00714_),
    .B1(_00683_),
    .C1(_00685_),
    .Y(_00720_));
 sky130_fd_sc_hd__a21o_1 _23911_ (.A1(_00476_),
    .A2(_00478_),
    .B1(_00474_),
    .X(_00721_));
 sky130_fd_sc_hd__a21oi_1 _23912_ (.A1(_00476_),
    .A2(_00478_),
    .B1(_00474_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand3_4 _23913_ (.A(_00719_),
    .B(_00720_),
    .C(_00721_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _23914_ (.A(_00718_),
    .B(_00722_),
    .Y(_00725_));
 sky130_fd_sc_hd__nand3_2 _23915_ (.A(_00717_),
    .B(_00718_),
    .C(_00722_),
    .Y(_00726_));
 sky130_fd_sc_hd__a21oi_4 _23916_ (.A1(_00724_),
    .A2(_00726_),
    .B1(_00585_),
    .Y(_00727_));
 sky130_fd_sc_hd__a21o_1 _23917_ (.A1(_00724_),
    .A2(_00726_),
    .B1(_00585_),
    .X(_00728_));
 sky130_fd_sc_hd__o211a_2 _23918_ (.A1(_00716_),
    .A2(_00725_),
    .B1(_00724_),
    .C1(_00585_),
    .X(_00729_));
 sky130_fd_sc_hd__o211ai_4 _23919_ (.A1(_00716_),
    .A2(_00725_),
    .B1(_00724_),
    .C1(_00585_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand3_2 _23920_ (.A(_00382_),
    .B(_00485_),
    .C(_00487_),
    .Y(_00731_));
 sky130_fd_sc_hd__o21ai_2 _23921_ (.A1(_00484_),
    .A2(_00486_),
    .B1(_00381_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand2_1 _23922_ (.A(_00381_),
    .B(_00731_),
    .Y(_00733_));
 sky130_fd_sc_hd__inv_2 _23923_ (.A(_00733_),
    .Y(_00735_));
 sky130_fd_sc_hd__o21a_4 _23924_ (.A1(_00357_),
    .A2(_00365_),
    .B1(_00364_),
    .X(_00736_));
 sky130_fd_sc_hd__o21ai_4 _23925_ (.A1(_00357_),
    .A2(_00365_),
    .B1(_00364_),
    .Y(_00737_));
 sky130_fd_sc_hd__o22a_4 _23926_ (.A1(_00342_),
    .A2(_00333_),
    .B1(net132),
    .B2(_00339_),
    .X(_00738_));
 sky130_fd_sc_hd__o22ai_1 _23927_ (.A1(_00342_),
    .A2(_00333_),
    .B1(net132),
    .B2(_00339_),
    .Y(_00739_));
 sky130_fd_sc_hd__o21ba_1 _23928_ (.A1(net146),
    .A2(_00322_),
    .B1_N(_00321_),
    .X(_00740_));
 sky130_fd_sc_hd__nor2_1 _23929_ (.A(_04048_),
    .B(_08660_),
    .Y(_00741_));
 sky130_fd_sc_hd__a31oi_4 _23930_ (.A1(_03952_),
    .A2(net233),
    .A3(_08657_),
    .B1(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__a31o_1 _23931_ (.A1(_03952_),
    .A2(net233),
    .A3(_08657_),
    .B1(_00741_),
    .X(_00743_));
 sky130_fd_sc_hd__nand3_4 _23932_ (.A(_00743_),
    .B(net159),
    .C(net33),
    .Y(_00744_));
 sky130_fd_sc_hd__o221a_1 _23933_ (.A1(_03961_),
    .A2(_08658_),
    .B1(_08660_),
    .B2(_04048_),
    .C1(_08878_),
    .X(_00746_));
 sky130_fd_sc_hd__nand2_2 _23934_ (.A(_08878_),
    .B(_00742_),
    .Y(_00747_));
 sky130_fd_sc_hd__o2bb2ai_2 _23935_ (.A1_N(_00742_),
    .A2_N(_08878_),
    .B1(_08881_),
    .B2(_09297_),
    .Y(_00748_));
 sky130_fd_sc_hd__a2bb2oi_2 _23936_ (.A1_N(_08881_),
    .A2_N(_09297_),
    .B1(_00744_),
    .B2(_00747_),
    .Y(_00749_));
 sky130_fd_sc_hd__a22o_1 _23937_ (.A1(_08882_),
    .A2(_09298_),
    .B1(_00744_),
    .B2(_00747_),
    .X(_00750_));
 sky130_fd_sc_hd__o2111a_1 _23938_ (.A1(_04495_),
    .A2(net150),
    .B1(_08882_),
    .C1(_00744_),
    .D1(_00747_),
    .X(_00751_));
 sky130_fd_sc_hd__o2111ai_4 _23939_ (.A1(_04495_),
    .A2(net150),
    .B1(_08882_),
    .C1(_00744_),
    .D1(_00747_),
    .Y(_00752_));
 sky130_fd_sc_hd__nand3_4 _23940_ (.A(_00740_),
    .B(_00750_),
    .C(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__o22a_1 _23941_ (.A1(_00321_),
    .A2(_00324_),
    .B1(_00749_),
    .B2(_00751_),
    .X(_00754_));
 sky130_fd_sc_hd__o22ai_4 _23942_ (.A1(_00321_),
    .A2(_00324_),
    .B1(_00749_),
    .B2(_00751_),
    .Y(_00755_));
 sky130_fd_sc_hd__a22o_1 _23943_ (.A1(net138),
    .A2(net134),
    .B1(_00753_),
    .B2(_00755_),
    .X(_00757_));
 sky130_fd_sc_hd__a31oi_2 _23944_ (.A1(_00740_),
    .A2(_00750_),
    .A3(_00752_),
    .B1(_10546_),
    .Y(_00758_));
 sky130_fd_sc_hd__nand4_2 _23945_ (.A(net138),
    .B(net134),
    .C(_00753_),
    .D(_00755_),
    .Y(_00759_));
 sky130_fd_sc_hd__o211ai_4 _23946_ (.A1(_10540_),
    .A2(net135),
    .B1(_00753_),
    .C1(_00755_),
    .Y(_00760_));
 sky130_fd_sc_hd__a21o_1 _23947_ (.A1(_00753_),
    .A2(_00755_),
    .B1(_10546_),
    .X(_00761_));
 sky130_fd_sc_hd__o21ai_2 _23948_ (.A1(_10546_),
    .A2(_00327_),
    .B1(_00331_),
    .Y(_00762_));
 sky130_fd_sc_hd__a21oi_1 _23949_ (.A1(_00328_),
    .A2(net133),
    .B1(_00330_),
    .Y(_00763_));
 sky130_fd_sc_hd__and3_1 _23950_ (.A(_00757_),
    .B(_00759_),
    .C(_00762_),
    .X(_00764_));
 sky130_fd_sc_hd__nand3_4 _23951_ (.A(_00757_),
    .B(_00759_),
    .C(_00762_),
    .Y(_00765_));
 sky130_fd_sc_hd__o2111ai_4 _23952_ (.A1(_10546_),
    .A2(_00327_),
    .B1(_00331_),
    .C1(_00760_),
    .D1(_00761_),
    .Y(_00766_));
 sky130_fd_sc_hd__a31oi_2 _23953_ (.A1(_00760_),
    .A2(_00761_),
    .A3(_00763_),
    .B1(net132),
    .Y(_00768_));
 sky130_fd_sc_hd__o311a_1 _23954_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_00765_),
    .C1(_00766_),
    .X(_00769_));
 sky130_fd_sc_hd__a21oi_2 _23955_ (.A1(_00765_),
    .A2(_00766_),
    .B1(_12099_),
    .Y(_00770_));
 sky130_fd_sc_hd__a22oi_1 _23956_ (.A1(_11743_),
    .A2(net142),
    .B1(_00766_),
    .B2(_00765_),
    .Y(_00771_));
 sky130_fd_sc_hd__o2bb2ai_2 _23957_ (.A1_N(_00765_),
    .A2_N(_00766_),
    .B1(_11042_),
    .B2(_11742_),
    .Y(_00772_));
 sky130_fd_sc_hd__o2111a_1 _23958_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net142),
    .C1(_00765_),
    .D1(_00766_),
    .X(_00773_));
 sky130_fd_sc_hd__o2111ai_4 _23959_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net142),
    .C1(_00765_),
    .D1(_00766_),
    .Y(_00774_));
 sky130_fd_sc_hd__a21oi_4 _23960_ (.A1(_00772_),
    .A2(_00774_),
    .B1(_00738_),
    .Y(_00775_));
 sky130_fd_sc_hd__nor3_2 _23961_ (.A(_00739_),
    .B(_00771_),
    .C(_00773_),
    .Y(_00776_));
 sky130_fd_sc_hd__o22ai_4 _23962_ (.A1(net130),
    .A2(_00366_),
    .B1(_00775_),
    .B2(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__a31oi_4 _23963_ (.A1(_00738_),
    .A2(_00772_),
    .A3(_00774_),
    .B1(_00737_),
    .Y(_00779_));
 sky130_fd_sc_hd__o31ai_4 _23964_ (.A1(_00738_),
    .A2(_00769_),
    .A3(_00770_),
    .B1(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__o21a_1 _23965_ (.A1(_00374_),
    .A2(_00375_),
    .B1(_00348_),
    .X(_00781_));
 sky130_fd_sc_hd__o21ai_2 _23966_ (.A1(_00374_),
    .A2(_00375_),
    .B1(_00348_),
    .Y(_00782_));
 sky130_fd_sc_hd__nand4_4 _23967_ (.A(_00350_),
    .B(_00777_),
    .C(_00780_),
    .D(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__a22oi_4 _23968_ (.A1(_00777_),
    .A2(_00780_),
    .B1(_00782_),
    .B2(_00350_),
    .Y(_00784_));
 sky130_fd_sc_hd__o2bb2ai_4 _23969_ (.A1_N(_00777_),
    .A2_N(_00780_),
    .B1(_00781_),
    .B2(_00349_),
    .Y(_00785_));
 sky130_fd_sc_hd__a32o_1 _23970_ (.A1(_13066_),
    .A2(_00039_),
    .A3(_00040_),
    .B1(net130),
    .B2(_00359_),
    .X(_00786_));
 sky130_fd_sc_hd__o211a_1 _23971_ (.A1(_11740_),
    .A2(_00359_),
    .B1(_00367_),
    .C1(_00786_),
    .X(_00787_));
 sky130_fd_sc_hd__o2bb2a_2 _23972_ (.A1_N(_00359_),
    .A2_N(net130),
    .B1(_00041_),
    .B2(_00368_),
    .X(_00788_));
 sky130_fd_sc_hd__nor2_2 _23973_ (.A(net319),
    .B(_03737_),
    .Y(_00790_));
 sky130_fd_sc_hd__or3_1 _23974_ (.A(net39),
    .B(net319),
    .C(_04037_),
    .X(_00791_));
 sky130_fd_sc_hd__a21oi_1 _23975_ (.A1(net150),
    .A2(_08668_),
    .B1(_03714_),
    .Y(_00792_));
 sky130_fd_sc_hd__o21ai_1 _23976_ (.A1(net159),
    .A2(_08666_),
    .B1(_03704_),
    .Y(_00793_));
 sky130_fd_sc_hd__nor2_1 _23977_ (.A(net25),
    .B(_02869_),
    .Y(_00794_));
 sky130_fd_sc_hd__a22oi_4 _23978_ (.A1(net25),
    .A2(_02880_),
    .B1(net163),
    .B2(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__a31o_4 _23979_ (.A1(net319),
    .A2(net161),
    .A3(_02858_),
    .B1(_00398_),
    .X(_00796_));
 sky130_fd_sc_hd__o21bai_2 _23980_ (.A1(_00790_),
    .A2(_00792_),
    .B1_N(_00795_),
    .Y(_00797_));
 sky130_fd_sc_hd__o211ai_4 _23981_ (.A1(net319),
    .A2(_03737_),
    .B1(_00795_),
    .C1(_00793_),
    .Y(_00798_));
 sky130_fd_sc_hd__a32o_2 _23982_ (.A1(net164),
    .A2(net161),
    .A3(net281),
    .B1(_04217_),
    .B2(net24),
    .X(_00799_));
 sky130_fd_sc_hd__a21oi_4 _23983_ (.A1(_00797_),
    .A2(_00798_),
    .B1(_00799_),
    .Y(_00801_));
 sky130_fd_sc_hd__a21o_1 _23984_ (.A1(_00797_),
    .A2(_00798_),
    .B1(_00799_),
    .X(_00802_));
 sky130_fd_sc_hd__o31a_2 _23985_ (.A1(_00790_),
    .A2(_00796_),
    .A3(_00792_),
    .B1(_00799_),
    .X(_00803_));
 sky130_fd_sc_hd__nand2_1 _23986_ (.A(_00798_),
    .B(_00799_),
    .Y(_00804_));
 sky130_fd_sc_hd__a22oi_2 _23987_ (.A1(_00038_),
    .A2(_00353_),
    .B1(_00802_),
    .B2(_00804_),
    .Y(_00805_));
 sky130_fd_sc_hd__o21ai_4 _23988_ (.A1(_00801_),
    .A2(_00803_),
    .B1(_00356_),
    .Y(_00806_));
 sky130_fd_sc_hd__a211oi_1 _23989_ (.A1(_00798_),
    .A2(_00799_),
    .B1(_00356_),
    .C1(_00801_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand4_1 _23990_ (.A(_00038_),
    .B(_00353_),
    .C(_00802_),
    .D(_00804_),
    .Y(_00808_));
 sky130_fd_sc_hd__nand2_1 _23991_ (.A(_00806_),
    .B(_00808_),
    .Y(_00809_));
 sky130_fd_sc_hd__o21a_2 _23992_ (.A1(_00805_),
    .A2(_00807_),
    .B1(_00406_),
    .X(_00810_));
 sky130_fd_sc_hd__o22ai_2 _23993_ (.A1(_00401_),
    .A2(_00404_),
    .B1(_00805_),
    .B2(_00807_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand3_1 _23994_ (.A(_00806_),
    .B(_00808_),
    .C(_00406_),
    .Y(_00813_));
 sky130_fd_sc_hd__a22oi_4 _23995_ (.A1(_00414_),
    .A2(_00410_),
    .B1(_00390_),
    .B2(_00413_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand3_4 _23996_ (.A(_00812_),
    .B(_00813_),
    .C(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__o2bb2a_2 _23997_ (.A1_N(_00406_),
    .A2_N(_00809_),
    .B1(_00423_),
    .B2(_00415_),
    .X(_00816_));
 sky130_fd_sc_hd__o2bb2ai_4 _23998_ (.A1_N(_00406_),
    .A2_N(_00809_),
    .B1(_00423_),
    .B2(_00415_),
    .Y(_00817_));
 sky130_fd_sc_hd__a21o_2 _23999_ (.A1(_00442_),
    .A2(_00451_),
    .B1(_00447_),
    .X(_00818_));
 sky130_fd_sc_hd__and3_1 _24000_ (.A(_04102_),
    .B(net20),
    .C(net42),
    .X(_00819_));
 sky130_fd_sc_hd__o311a_1 _24001_ (.A1(net244),
    .A2(net241),
    .A3(_07074_),
    .B1(_04895_),
    .C1(_07072_),
    .X(_00820_));
 sky130_fd_sc_hd__a31o_1 _24002_ (.A1(_07072_),
    .A2(net169),
    .A3(_04895_),
    .B1(_00819_),
    .X(_00821_));
 sky130_fd_sc_hd__o211ai_4 _24003_ (.A1(net169),
    .A2(_07765_),
    .B1(_04267_),
    .C1(_07771_),
    .Y(_00823_));
 sky130_fd_sc_hd__or3b_1 _24004_ (.A(net41),
    .B(_04245_),
    .C_N(net40),
    .X(_00824_));
 sky130_fd_sc_hd__a31oi_2 _24005_ (.A1(_03957_),
    .A2(_05926_),
    .A3(_07500_),
    .B1(_04481_),
    .Y(_00825_));
 sky130_fd_sc_hd__o21ai_2 _24006_ (.A1(_04223_),
    .A2(_07075_),
    .B1(_00825_),
    .Y(_00826_));
 sky130_fd_sc_hd__or3b_1 _24007_ (.A(net42),
    .B(_04223_),
    .C_N(net41),
    .X(_00827_));
 sky130_fd_sc_hd__a22oi_1 _24008_ (.A1(net21),
    .A2(_04482_),
    .B1(_00825_),
    .B2(_07499_),
    .Y(_00828_));
 sky130_fd_sc_hd__a21oi_1 _24009_ (.A1(_00823_),
    .A2(_00824_),
    .B1(_00828_),
    .Y(_00829_));
 sky130_fd_sc_hd__a22o_1 _24010_ (.A1(_00823_),
    .A2(_00824_),
    .B1(_00826_),
    .B2(_00827_),
    .X(_00830_));
 sky130_fd_sc_hd__o2111ai_4 _24011_ (.A1(_04245_),
    .A2(_04270_),
    .B1(_00823_),
    .C1(_00826_),
    .D1(_00827_),
    .Y(_00831_));
 sky130_fd_sc_hd__a21o_2 _24012_ (.A1(_00830_),
    .A2(_00831_),
    .B1(_00821_),
    .X(_00832_));
 sky130_fd_sc_hd__o211ai_4 _24013_ (.A1(_00819_),
    .A2(_00820_),
    .B1(_00830_),
    .C1(_00831_),
    .Y(_00834_));
 sky130_fd_sc_hd__a21oi_2 _24014_ (.A1(_00832_),
    .A2(_00834_),
    .B1(_00818_),
    .Y(_00835_));
 sky130_fd_sc_hd__a21o_2 _24015_ (.A1(_00832_),
    .A2(_00834_),
    .B1(_00818_),
    .X(_00836_));
 sky130_fd_sc_hd__nand3_4 _24016_ (.A(_00818_),
    .B(_00832_),
    .C(_00834_),
    .Y(_00837_));
 sky130_fd_sc_hd__o22a_1 _24017_ (.A1(_04168_),
    .A2(_05465_),
    .B1(_06222_),
    .B2(_05463_),
    .X(_00838_));
 sky130_fd_sc_hd__a32o_1 _24018_ (.A1(net202),
    .A2(net173),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net17),
    .X(_00839_));
 sky130_fd_sc_hd__a32oi_4 _24019_ (.A1(net197),
    .A2(_06452_),
    .A3(_05225_),
    .B1(_05228_),
    .B2(net18),
    .Y(_00840_));
 sky130_fd_sc_hd__a32o_1 _24020_ (.A1(net197),
    .A2(_06452_),
    .A3(_05225_),
    .B1(_05228_),
    .B2(net18),
    .X(_00841_));
 sky130_fd_sc_hd__a32oi_4 _24021_ (.A1(net191),
    .A2(_06762_),
    .A3(net242),
    .B1(_04988_),
    .B2(net19),
    .Y(_00842_));
 sky130_fd_sc_hd__a32o_1 _24022_ (.A1(net191),
    .A2(_06762_),
    .A3(net242),
    .B1(_04988_),
    .B2(net19),
    .X(_00843_));
 sky130_fd_sc_hd__nand2_2 _24023_ (.A(_00840_),
    .B(_00842_),
    .Y(_00845_));
 sky130_fd_sc_hd__nor2_1 _24024_ (.A(_00840_),
    .B(_00842_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _24025_ (.A(_00841_),
    .B(_00843_),
    .Y(_00847_));
 sky130_fd_sc_hd__a21o_2 _24026_ (.A1(_00845_),
    .A2(_00847_),
    .B1(_00839_),
    .X(_00848_));
 sky130_fd_sc_hd__nand3_4 _24027_ (.A(_00839_),
    .B(_00845_),
    .C(_00847_),
    .Y(_00849_));
 sky130_fd_sc_hd__nand2_2 _24028_ (.A(_00848_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__a22oi_4 _24029_ (.A1(_00836_),
    .A2(_00837_),
    .B1(_00848_),
    .B2(_00849_),
    .Y(_00851_));
 sky130_fd_sc_hd__and4_1 _24030_ (.A(_00836_),
    .B(_00837_),
    .C(_00848_),
    .D(_00849_),
    .X(_00852_));
 sky130_fd_sc_hd__and3_2 _24031_ (.A(_00836_),
    .B(_00837_),
    .C(_00850_),
    .X(_00853_));
 sky130_fd_sc_hd__a21oi_4 _24032_ (.A1(_00836_),
    .A2(_00837_),
    .B1(_00850_),
    .Y(_00854_));
 sky130_fd_sc_hd__o221ai_4 _24033_ (.A1(_00851_),
    .A2(_00852_),
    .B1(_00814_),
    .B2(_00810_),
    .C1(_00815_),
    .Y(_00856_));
 sky130_fd_sc_hd__o2bb2ai_2 _24034_ (.A1_N(_00815_),
    .A2_N(_00817_),
    .B1(_00853_),
    .B2(_00854_),
    .Y(_00857_));
 sky130_fd_sc_hd__o2bb2ai_2 _24035_ (.A1_N(_00815_),
    .A2_N(_00817_),
    .B1(_00851_),
    .B2(_00852_),
    .Y(_00858_));
 sky130_fd_sc_hd__o21a_1 _24036_ (.A1(_00853_),
    .A2(_00854_),
    .B1(_00815_),
    .X(_00859_));
 sky130_fd_sc_hd__o21ai_4 _24037_ (.A1(_00853_),
    .A2(_00854_),
    .B1(_00815_),
    .Y(_00860_));
 sky130_fd_sc_hd__o221ai_4 _24038_ (.A1(_00853_),
    .A2(_00854_),
    .B1(_00814_),
    .B2(_00810_),
    .C1(_00815_),
    .Y(_00861_));
 sky130_fd_sc_hd__a22oi_2 _24039_ (.A1(_00369_),
    .A2(_00786_),
    .B1(_00858_),
    .B2(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand3_4 _24040_ (.A(_00788_),
    .B(_00856_),
    .C(_00857_),
    .Y(_00863_));
 sky130_fd_sc_hd__o211a_4 _24041_ (.A1(_00816_),
    .A2(_00860_),
    .B1(_00787_),
    .C1(_00858_),
    .X(_00864_));
 sky130_fd_sc_hd__nand3_4 _24042_ (.A(_00858_),
    .B(_00861_),
    .C(_00787_),
    .Y(_00865_));
 sky130_fd_sc_hd__o32a_1 _24043_ (.A1(_00080_),
    .A2(_00385_),
    .A3(_00421_),
    .B1(_00464_),
    .B2(_00465_),
    .X(_00867_));
 sky130_fd_sc_hd__a32o_1 _24044_ (.A1(_00081_),
    .A2(_00386_),
    .A3(_00422_),
    .B1(_00425_),
    .B2(_00467_),
    .X(_00868_));
 sky130_fd_sc_hd__o2bb2a_1 _24045_ (.A1_N(_00425_),
    .A2_N(_00467_),
    .B1(_00388_),
    .B2(_00421_),
    .X(_00869_));
 sky130_fd_sc_hd__a21oi_1 _24046_ (.A1(_00863_),
    .A2(_00865_),
    .B1(_00868_),
    .Y(_00870_));
 sky130_fd_sc_hd__a21o_1 _24047_ (.A1(_00863_),
    .A2(_00865_),
    .B1(_00868_),
    .X(_00871_));
 sky130_fd_sc_hd__a31oi_2 _24048_ (.A1(_00788_),
    .A2(_00856_),
    .A3(_00857_),
    .B1(_00869_),
    .Y(_00872_));
 sky130_fd_sc_hd__a31o_1 _24049_ (.A1(_00788_),
    .A2(_00856_),
    .A3(_00857_),
    .B1(_00869_),
    .X(_00873_));
 sky130_fd_sc_hd__and3_1 _24050_ (.A(_00863_),
    .B(_00865_),
    .C(_00868_),
    .X(_00874_));
 sky130_fd_sc_hd__a21oi_1 _24051_ (.A1(_00863_),
    .A2(_00865_),
    .B1(_00869_),
    .Y(_00875_));
 sky130_fd_sc_hd__o22ai_4 _24052_ (.A1(_00426_),
    .A2(_00472_),
    .B1(_00862_),
    .B2(_00864_),
    .Y(_00876_));
 sky130_fd_sc_hd__and3_1 _24053_ (.A(_00863_),
    .B(_00865_),
    .C(_00869_),
    .X(_00878_));
 sky130_fd_sc_hd__o211ai_4 _24054_ (.A1(_00424_),
    .A2(_00867_),
    .B1(_00865_),
    .C1(_00863_),
    .Y(_00879_));
 sky130_fd_sc_hd__o21ai_1 _24055_ (.A1(_00864_),
    .A2(_00873_),
    .B1(_00871_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand4_4 _24056_ (.A(_00783_),
    .B(_00785_),
    .C(_00876_),
    .D(_00879_),
    .Y(_00881_));
 sky130_fd_sc_hd__o2bb2ai_2 _24057_ (.A1_N(_00783_),
    .A2_N(_00785_),
    .B1(_00875_),
    .B2(_00878_),
    .Y(_00882_));
 sky130_fd_sc_hd__o2bb2ai_4 _24058_ (.A1_N(_00783_),
    .A2_N(_00785_),
    .B1(_00870_),
    .B2(_00874_),
    .Y(_00883_));
 sky130_fd_sc_hd__o211ai_1 _24059_ (.A1(_00864_),
    .A2(_00873_),
    .B1(_00871_),
    .C1(_00783_),
    .Y(_00884_));
 sky130_fd_sc_hd__o2111ai_4 _24060_ (.A1(_00864_),
    .A2(_00873_),
    .B1(_00871_),
    .C1(_00783_),
    .D1(_00785_),
    .Y(_00885_));
 sky130_fd_sc_hd__o21ai_1 _24061_ (.A1(_00784_),
    .A2(_00884_),
    .B1(_00883_),
    .Y(_00886_));
 sky130_fd_sc_hd__o21a_1 _24062_ (.A1(_00784_),
    .A2(_00884_),
    .B1(_00883_),
    .X(_00887_));
 sky130_fd_sc_hd__a22oi_4 _24063_ (.A1(_00381_),
    .A2(_00731_),
    .B1(_00883_),
    .B2(_00885_),
    .Y(_00889_));
 sky130_fd_sc_hd__nand4_4 _24064_ (.A(_00382_),
    .B(_00732_),
    .C(_00881_),
    .D(_00882_),
    .Y(_00890_));
 sky130_fd_sc_hd__a22oi_4 _24065_ (.A1(_00382_),
    .A2(_00732_),
    .B1(_00881_),
    .B2(_00882_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand4_4 _24066_ (.A(_00381_),
    .B(_00731_),
    .C(_00883_),
    .D(_00885_),
    .Y(_00892_));
 sky130_fd_sc_hd__o211ai_2 _24067_ (.A1(_00727_),
    .A2(_00729_),
    .B1(_00890_),
    .C1(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__o211ai_2 _24068_ (.A1(_00889_),
    .A2(_00891_),
    .B1(_00728_),
    .C1(_00730_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand4_4 _24069_ (.A(_00728_),
    .B(_00730_),
    .C(_00890_),
    .D(_00892_),
    .Y(_00895_));
 sky130_fd_sc_hd__o22ai_4 _24070_ (.A1(_00727_),
    .A2(_00729_),
    .B1(_00889_),
    .B2(_00891_),
    .Y(_00896_));
 sky130_fd_sc_hd__nand4_4 _24071_ (.A(_00494_),
    .B(_00633_),
    .C(_00895_),
    .D(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__a22oi_4 _24072_ (.A1(_00494_),
    .A2(_00633_),
    .B1(_00895_),
    .B2(_00896_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand3_1 _24073_ (.A(_00894_),
    .B(_00634_),
    .C(_00893_),
    .Y(_00900_));
 sky130_fd_sc_hd__a2bb2oi_1 _24074_ (.A1_N(_00589_),
    .A2_N(_00598_),
    .B1(_00897_),
    .B2(_00900_),
    .Y(_00901_));
 sky130_fd_sc_hd__a21o_1 _24075_ (.A1(_00897_),
    .A2(_00900_),
    .B1(_00600_),
    .X(_00902_));
 sky130_fd_sc_hd__a31oi_2 _24076_ (.A1(_00894_),
    .A2(_00634_),
    .A3(_00893_),
    .B1(_00599_),
    .Y(_00903_));
 sky130_fd_sc_hd__o211a_1 _24077_ (.A1(_00587_),
    .A2(_00591_),
    .B1(_00897_),
    .C1(_00900_),
    .X(_00904_));
 sky130_fd_sc_hd__nand2_1 _24078_ (.A(_00903_),
    .B(_00897_),
    .Y(_00905_));
 sky130_fd_sc_hd__a31oi_2 _24079_ (.A1(_00636_),
    .A2(_00895_),
    .A3(_00896_),
    .B1(_00600_),
    .Y(_00906_));
 sky130_fd_sc_hd__o21ai_2 _24080_ (.A1(_00599_),
    .A2(_00898_),
    .B1(_00897_),
    .Y(_00907_));
 sky130_fd_sc_hd__o21ai_1 _24081_ (.A1(_00263_),
    .A2(_00269_),
    .B1(_00609_),
    .Y(_00908_));
 sky130_fd_sc_hd__nand2_1 _24082_ (.A(_00610_),
    .B(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__a221oi_2 _24083_ (.A1(_00610_),
    .A2(_00908_),
    .B1(_00903_),
    .B2(_00897_),
    .C1(_00901_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand3_2 _24084_ (.A(_00902_),
    .B(_00905_),
    .C(_00909_),
    .Y(_00912_));
 sky130_fd_sc_hd__a21oi_2 _24085_ (.A1(_00902_),
    .A2(_00905_),
    .B1(_00909_),
    .Y(_00913_));
 sky130_fd_sc_hd__o21bai_2 _24086_ (.A1(_00901_),
    .A2(_00904_),
    .B1_N(_00909_),
    .Y(_00914_));
 sky130_fd_sc_hd__o211a_1 _24087_ (.A1(_00568_),
    .A2(_00577_),
    .B1(_00912_),
    .C1(_00914_),
    .X(_00915_));
 sky130_fd_sc_hd__o211ai_4 _24088_ (.A1(_00568_),
    .A2(_00577_),
    .B1(_00912_),
    .C1(_00914_),
    .Y(_00916_));
 sky130_fd_sc_hd__o22a_1 _24089_ (.A1(_00572_),
    .A2(_00631_),
    .B1(_00911_),
    .B2(_00913_),
    .X(_00917_));
 sky130_fd_sc_hd__o22ai_2 _24090_ (.A1(_00572_),
    .A2(_00631_),
    .B1(_00911_),
    .B2(_00913_),
    .Y(_00918_));
 sky130_fd_sc_hd__a2bb2oi_1 _24091_ (.A1_N(_00616_),
    .A2_N(_00622_),
    .B1(_00916_),
    .B2(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__o22ai_1 _24092_ (.A1(_00616_),
    .A2(_00622_),
    .B1(_00915_),
    .B2(_00917_),
    .Y(_00920_));
 sky130_fd_sc_hd__o211a_1 _24093_ (.A1(_00618_),
    .A2(_00623_),
    .B1(_00916_),
    .C1(_00918_),
    .X(_00922_));
 sky130_fd_sc_hd__o211ai_2 _24094_ (.A1(_00618_),
    .A2(_00623_),
    .B1(_00916_),
    .C1(_00918_),
    .Y(_00923_));
 sky130_fd_sc_hd__nor2_1 _24095_ (.A(_00919_),
    .B(_00922_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand2_1 _24096_ (.A(_00920_),
    .B(_00923_),
    .Y(_00925_));
 sky130_fd_sc_hd__and4_1 _24097_ (.A(_00298_),
    .B(_00300_),
    .C(_00627_),
    .D(_00628_),
    .X(_00926_));
 sky130_fd_sc_hd__a21boi_2 _24098_ (.A1(_00300_),
    .A2(_00628_),
    .B1_N(_00627_),
    .Y(_00927_));
 sky130_fd_sc_hd__a21oi_1 _24099_ (.A1(_00309_),
    .A2(_00926_),
    .B1(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__xor2_1 _24100_ (.A(_00925_),
    .B(_00928_),
    .X(net105));
 sky130_fd_sc_hd__a31o_1 _24101_ (.A1(_00705_),
    .A2(_00706_),
    .A3(_00708_),
    .B1(_00714_),
    .X(_00929_));
 sky130_fd_sc_hd__inv_2 _24102_ (.A(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__o22ai_4 _24103_ (.A1(_00733_),
    .A2(_00886_),
    .B1(_00727_),
    .B2(_00729_),
    .Y(_00932_));
 sky130_fd_sc_hd__o31a_1 _24104_ (.A1(_00727_),
    .A2(_00729_),
    .A3(_00889_),
    .B1(_00892_),
    .X(_00933_));
 sky130_fd_sc_hd__or3_1 _24105_ (.A(net54),
    .B(_04266_),
    .C(_04412_),
    .X(_00934_));
 sky130_fd_sc_hd__or3b_2 _24106_ (.A(_04069_),
    .B(net56),
    .C_N(net54),
    .X(_00935_));
 sky130_fd_sc_hd__o31a_1 _24107_ (.A1(net54),
    .A2(_04266_),
    .A3(_04412_),
    .B1(_00935_),
    .X(_00936_));
 sky130_fd_sc_hd__nand2_1 _24108_ (.A(_00703_),
    .B(_00706_),
    .Y(_00937_));
 sky130_fd_sc_hd__a32o_1 _24109_ (.A1(net220),
    .A2(net186),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net10),
    .X(_00938_));
 sky130_fd_sc_hd__a31oi_1 _24110_ (.A1(_00692_),
    .A2(_00693_),
    .A3(_00694_),
    .B1(_00688_),
    .Y(_00939_));
 sky130_fd_sc_hd__a21oi_1 _24111_ (.A1(_00689_),
    .A2(_00695_),
    .B1(_00696_),
    .Y(_00940_));
 sky130_fd_sc_hd__a32o_1 _24112_ (.A1(net184),
    .A2(net213),
    .A3(net239),
    .B1(_07308_),
    .B2(net11),
    .X(_00941_));
 sky130_fd_sc_hd__nand3_2 _24113_ (.A(_05290_),
    .B(_05292_),
    .C(net240),
    .Y(_00943_));
 sky130_fd_sc_hd__or3_1 _24114_ (.A(net51),
    .B(_04190_),
    .C(_04135_),
    .X(_00944_));
 sky130_fd_sc_hd__nor2_1 _24115_ (.A(_04113_),
    .B(_07226_),
    .Y(_00945_));
 sky130_fd_sc_hd__o311a_1 _24116_ (.A1(net11),
    .A2(_04557_),
    .A3(net208),
    .B1(net269),
    .C1(net209),
    .X(_00946_));
 sky130_fd_sc_hd__a31oi_2 _24117_ (.A1(net209),
    .A2(_05074_),
    .A3(net269),
    .B1(_00945_),
    .Y(_00947_));
 sky130_fd_sc_hd__o211ai_4 _24118_ (.A1(_04135_),
    .A2(_06866_),
    .B1(_00943_),
    .C1(_00947_),
    .Y(_00948_));
 sky130_fd_sc_hd__a21oi_1 _24119_ (.A1(_00943_),
    .A2(_00944_),
    .B1(_00947_),
    .Y(_00949_));
 sky130_fd_sc_hd__o2bb2ai_2 _24120_ (.A1_N(_00943_),
    .A2_N(_00944_),
    .B1(_00945_),
    .B2(_00946_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand2_1 _24121_ (.A(_00941_),
    .B(_00948_),
    .Y(_00951_));
 sky130_fd_sc_hd__a21oi_1 _24122_ (.A1(_00941_),
    .A2(_00948_),
    .B1(_00949_),
    .Y(_00952_));
 sky130_fd_sc_hd__a21oi_2 _24123_ (.A1(_00948_),
    .A2(_00950_),
    .B1(_00941_),
    .Y(_00954_));
 sky130_fd_sc_hd__a21o_1 _24124_ (.A1(_00948_),
    .A2(_00950_),
    .B1(_00941_),
    .X(_00955_));
 sky130_fd_sc_hd__and3_1 _24125_ (.A(_00941_),
    .B(_00948_),
    .C(_00950_),
    .X(_00956_));
 sky130_fd_sc_hd__nand3_1 _24126_ (.A(_00941_),
    .B(_00948_),
    .C(_00950_),
    .Y(_00957_));
 sky130_fd_sc_hd__o22ai_2 _24127_ (.A1(_00696_),
    .A2(_00939_),
    .B1(_00949_),
    .B2(_00951_),
    .Y(_00958_));
 sky130_fd_sc_hd__nor2_1 _24128_ (.A(_00954_),
    .B(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__a21boi_1 _24129_ (.A1(_00955_),
    .A2(_00957_),
    .B1_N(_00940_),
    .Y(_00960_));
 sky130_fd_sc_hd__o21ai_1 _24130_ (.A1(_00954_),
    .A2(_00956_),
    .B1(_00940_),
    .Y(_00961_));
 sky130_fd_sc_hd__o21bai_2 _24131_ (.A1(_00959_),
    .A2(_00960_),
    .B1_N(_00938_),
    .Y(_00962_));
 sky130_fd_sc_hd__o211ai_2 _24132_ (.A1(_00958_),
    .A2(_00954_),
    .B1(_00938_),
    .C1(_00961_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _24133_ (.A(_00962_),
    .B(_00963_),
    .Y(_00965_));
 sky130_fd_sc_hd__a21oi_4 _24134_ (.A1(_00703_),
    .A2(_00706_),
    .B1(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__a21oi_2 _24135_ (.A1(_00962_),
    .A2(_00963_),
    .B1(_00937_),
    .Y(_00967_));
 sky130_fd_sc_hd__a31o_1 _24136_ (.A1(_00703_),
    .A2(_00706_),
    .A3(_00965_),
    .B1(_00936_),
    .X(_00968_));
 sky130_fd_sc_hd__a211oi_4 _24137_ (.A1(_00934_),
    .A2(_00935_),
    .B1(_00966_),
    .C1(_00967_),
    .Y(_00969_));
 sky130_fd_sc_hd__o221a_1 _24138_ (.A1(_04069_),
    .A2(_08007_),
    .B1(_00966_),
    .B2(_00967_),
    .C1(_00934_),
    .X(_00970_));
 sky130_fd_sc_hd__o21ai_1 _24139_ (.A1(_00966_),
    .A2(_00967_),
    .B1(_00936_),
    .Y(_00971_));
 sky130_fd_sc_hd__o21ai_1 _24140_ (.A1(_00966_),
    .A2(_00968_),
    .B1(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__o31a_1 _24141_ (.A1(_00654_),
    .A2(_00656_),
    .A3(_00660_),
    .B1(_00665_),
    .X(_00973_));
 sky130_fd_sc_hd__nand2_1 _24142_ (.A(_00662_),
    .B(_00665_),
    .Y(_00974_));
 sky130_fd_sc_hd__a32oi_4 _24143_ (.A1(_00818_),
    .A2(_00832_),
    .A3(_00834_),
    .B1(_00848_),
    .B2(_00849_),
    .Y(_00976_));
 sky130_fd_sc_hd__o21ai_2 _24144_ (.A1(_00850_),
    .A2(_00835_),
    .B1(_00837_),
    .Y(_00977_));
 sky130_fd_sc_hd__a21o_1 _24145_ (.A1(_00652_),
    .A2(_00653_),
    .B1(_00649_),
    .X(_00978_));
 sky130_fd_sc_hd__o21ai_1 _24146_ (.A1(_00840_),
    .A2(_00842_),
    .B1(_00838_),
    .Y(_00979_));
 sky130_fd_sc_hd__a21oi_1 _24147_ (.A1(_00840_),
    .A2(_00842_),
    .B1(_00838_),
    .Y(_00980_));
 sky130_fd_sc_hd__o311a_1 _24148_ (.A1(net233),
    .A2(_04787_),
    .A3(_05551_),
    .B1(net273),
    .C1(net178),
    .X(_00981_));
 sky130_fd_sc_hd__and3_1 _24149_ (.A(_04190_),
    .B(net49),
    .C(net15),
    .X(_00982_));
 sky130_fd_sc_hd__a31o_1 _24150_ (.A1(net178),
    .A2(_05553_),
    .A3(net273),
    .B1(_00982_),
    .X(_00983_));
 sky130_fd_sc_hd__nor2_1 _24151_ (.A(_04168_),
    .B(_05766_),
    .Y(_00984_));
 sky130_fd_sc_hd__a31oi_2 _24152_ (.A1(net202),
    .A2(net173),
    .A3(_05762_),
    .B1(_00984_),
    .Y(_00985_));
 sky130_fd_sc_hd__nor2_1 _24153_ (.A(_04157_),
    .B(_06030_),
    .Y(_00987_));
 sky130_fd_sc_hd__a221oi_2 _24154_ (.A1(_03957_),
    .A2(_05926_),
    .B1(_05553_),
    .B2(net16),
    .C1(_06028_),
    .Y(_00988_));
 sky130_fd_sc_hd__a211o_1 _24155_ (.A1(_05553_),
    .A2(net16),
    .B1(_06028_),
    .C1(net204),
    .X(_00989_));
 sky130_fd_sc_hd__o211ai_4 _24156_ (.A1(_04157_),
    .A2(_06030_),
    .B1(_00985_),
    .C1(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__o21ba_1 _24157_ (.A1(_00987_),
    .A2(_00988_),
    .B1_N(_00985_),
    .X(_00991_));
 sky130_fd_sc_hd__o21bai_2 _24158_ (.A1(_00987_),
    .A2(_00988_),
    .B1_N(_00985_),
    .Y(_00992_));
 sky130_fd_sc_hd__o211a_1 _24159_ (.A1(_00981_),
    .A2(_00982_),
    .B1(_00990_),
    .C1(_00992_),
    .X(_00993_));
 sky130_fd_sc_hd__o211ai_2 _24160_ (.A1(_00981_),
    .A2(_00982_),
    .B1(_00990_),
    .C1(_00992_),
    .Y(_00994_));
 sky130_fd_sc_hd__a21oi_1 _24161_ (.A1(_00990_),
    .A2(_00992_),
    .B1(_00983_),
    .Y(_00995_));
 sky130_fd_sc_hd__a21o_1 _24162_ (.A1(_00990_),
    .A2(_00992_),
    .B1(_00983_),
    .X(_00996_));
 sky130_fd_sc_hd__o211ai_4 _24163_ (.A1(_00846_),
    .A2(_00980_),
    .B1(_00994_),
    .C1(_00996_),
    .Y(_00998_));
 sky130_fd_sc_hd__inv_2 _24164_ (.A(_00998_),
    .Y(_00999_));
 sky130_fd_sc_hd__o2bb2ai_4 _24165_ (.A1_N(_00845_),
    .A2_N(_00979_),
    .B1(_00993_),
    .B2(_00995_),
    .Y(_01000_));
 sky130_fd_sc_hd__o21a_1 _24166_ (.A1(_00649_),
    .A2(_00656_),
    .B1(_01000_),
    .X(_01001_));
 sky130_fd_sc_hd__o21ai_1 _24167_ (.A1(_00649_),
    .A2(_00656_),
    .B1(_01000_),
    .Y(_01002_));
 sky130_fd_sc_hd__o211a_2 _24168_ (.A1(_00649_),
    .A2(_00656_),
    .B1(_00998_),
    .C1(_01000_),
    .X(_01003_));
 sky130_fd_sc_hd__a21oi_2 _24169_ (.A1(_00998_),
    .A2(_01000_),
    .B1(_00978_),
    .Y(_01004_));
 sky130_fd_sc_hd__a21o_1 _24170_ (.A1(_00998_),
    .A2(_01000_),
    .B1(_00978_),
    .X(_01005_));
 sky130_fd_sc_hd__nand2_1 _24171_ (.A(_00977_),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__o211ai_4 _24172_ (.A1(_00999_),
    .A2(_01002_),
    .B1(_01005_),
    .C1(_00977_),
    .Y(_01007_));
 sky130_fd_sc_hd__a21o_1 _24173_ (.A1(_00662_),
    .A2(_00665_),
    .B1(_01007_),
    .X(_01009_));
 sky130_fd_sc_hd__o22ai_4 _24174_ (.A1(_00835_),
    .A2(_00976_),
    .B1(_01003_),
    .B2(_01004_),
    .Y(_01010_));
 sky130_fd_sc_hd__inv_2 _24175_ (.A(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__o221ai_2 _24176_ (.A1(_00835_),
    .A2(_00976_),
    .B1(_01003_),
    .B2(_01004_),
    .C1(_00973_),
    .Y(_01012_));
 sky130_fd_sc_hd__o311a_1 _24177_ (.A1(_00654_),
    .A2(_00656_),
    .A3(_00660_),
    .B1(_00665_),
    .C1(_01007_),
    .X(_01013_));
 sky130_fd_sc_hd__nand2_1 _24178_ (.A(_00974_),
    .B(_01010_),
    .Y(_01014_));
 sky130_fd_sc_hd__o21ai_1 _24179_ (.A1(_01003_),
    .A2(_01006_),
    .B1(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__o211ai_2 _24180_ (.A1(_01003_),
    .A2(_01006_),
    .B1(_01012_),
    .C1(_01014_),
    .Y(_01016_));
 sky130_fd_sc_hd__a21o_1 _24181_ (.A1(_01007_),
    .A2(_01010_),
    .B1(_00974_),
    .X(_01017_));
 sky130_fd_sc_hd__o211ai_2 _24182_ (.A1(_01003_),
    .A2(_01006_),
    .B1(_01010_),
    .C1(_00974_),
    .Y(_01018_));
 sky130_fd_sc_hd__a21boi_2 _24183_ (.A1(_00672_),
    .A2(_00675_),
    .B1_N(_00674_),
    .Y(_01020_));
 sky130_fd_sc_hd__a2bb2oi_1 _24184_ (.A1_N(_00673_),
    .A2_N(_00678_),
    .B1(_01009_),
    .B2(_01016_),
    .Y(_01021_));
 sky130_fd_sc_hd__o211ai_4 _24185_ (.A1(_00673_),
    .A2(_00678_),
    .B1(_01017_),
    .C1(_01018_),
    .Y(_01022_));
 sky130_fd_sc_hd__o211a_1 _24186_ (.A1(_00973_),
    .A2(_01007_),
    .B1(_01020_),
    .C1(_01016_),
    .X(_01023_));
 sky130_fd_sc_hd__o211ai_2 _24187_ (.A1(_00973_),
    .A2(_01007_),
    .B1(_01020_),
    .C1(_01016_),
    .Y(_01024_));
 sky130_fd_sc_hd__o2111ai_2 _24188_ (.A1(_00966_),
    .A2(_00968_),
    .B1(_00971_),
    .C1(_01022_),
    .D1(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__o22ai_2 _24189_ (.A1(_00969_),
    .A2(_00970_),
    .B1(_01021_),
    .B2(_01023_),
    .Y(_01026_));
 sky130_fd_sc_hd__a21o_1 _24190_ (.A1(_01022_),
    .A2(_01024_),
    .B1(_00972_),
    .X(_01027_));
 sky130_fd_sc_hd__o211ai_1 _24191_ (.A1(_00969_),
    .A2(_00970_),
    .B1(_01022_),
    .C1(_01024_),
    .Y(_01028_));
 sky130_fd_sc_hd__a21boi_1 _24192_ (.A1(_00863_),
    .A2(_00868_),
    .B1_N(_00865_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand3_2 _24193_ (.A(_01027_),
    .B(_01028_),
    .C(_01029_),
    .Y(_01031_));
 sky130_fd_sc_hd__o211a_2 _24194_ (.A1(_00864_),
    .A2(_00872_),
    .B1(_01025_),
    .C1(_01026_),
    .X(_01032_));
 sky130_fd_sc_hd__o211ai_2 _24195_ (.A1(_00864_),
    .A2(_00872_),
    .B1(_01025_),
    .C1(_01026_),
    .Y(_01033_));
 sky130_fd_sc_hd__o32a_1 _24196_ (.A1(_00637_),
    .A2(_00676_),
    .A3(_00680_),
    .B1(_00713_),
    .B2(_00714_),
    .X(_01034_));
 sky130_fd_sc_hd__o21a_1 _24197_ (.A1(_00684_),
    .A2(_00715_),
    .B1(_00683_),
    .X(_01035_));
 sky130_fd_sc_hd__a21oi_1 _24198_ (.A1(_01031_),
    .A2(_01033_),
    .B1(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__o2bb2ai_2 _24199_ (.A1_N(_01031_),
    .A2_N(_01033_),
    .B1(_01034_),
    .B2(_00682_),
    .Y(_01037_));
 sky130_fd_sc_hd__nand2_2 _24200_ (.A(_01031_),
    .B(_01035_),
    .Y(_01038_));
 sky130_fd_sc_hd__and3_2 _24201_ (.A(_01031_),
    .B(_01033_),
    .C(_01035_),
    .X(_01039_));
 sky130_fd_sc_hd__o21ai_2 _24202_ (.A1(_01032_),
    .A2(_01038_),
    .B1(_01037_),
    .Y(_01040_));
 sky130_fd_sc_hd__o31a_1 _24203_ (.A1(_00738_),
    .A2(_00769_),
    .A3(_00770_),
    .B1(_00737_),
    .X(_01042_));
 sky130_fd_sc_hd__a31o_1 _24204_ (.A1(_00757_),
    .A2(_00759_),
    .A3(_00762_),
    .B1(_12099_),
    .X(_01043_));
 sky130_fd_sc_hd__o21ai_1 _24205_ (.A1(_10540_),
    .A2(net135),
    .B1(_00755_),
    .Y(_01044_));
 sky130_fd_sc_hd__a21oi_1 _24206_ (.A1(_00753_),
    .A2(net133),
    .B1(_00754_),
    .Y(_01045_));
 sky130_fd_sc_hd__o211a_1 _24207_ (.A1(_00742_),
    .A2(_08878_),
    .B1(_08882_),
    .C1(_09298_),
    .X(_01046_));
 sky130_fd_sc_hd__o21ai_1 _24208_ (.A1(_08878_),
    .A2(_00742_),
    .B1(_00748_),
    .Y(_01047_));
 sky130_fd_sc_hd__o41a_1 _24209_ (.A1(_03286_),
    .A2(net25),
    .A3(_08207_),
    .A4(_00742_),
    .B1(_00748_),
    .X(_01048_));
 sky130_fd_sc_hd__o41ai_4 _24210_ (.A1(net8),
    .A2(net267),
    .A3(_06508_),
    .A4(net244),
    .B1(_08657_),
    .Y(_01049_));
 sky130_fd_sc_hd__o32a_1 _24211_ (.A1(_04059_),
    .A2(_04266_),
    .A3(net57),
    .B1(_04131_),
    .B2(_01049_),
    .X(_01050_));
 sky130_fd_sc_hd__o22ai_4 _24212_ (.A1(_04059_),
    .A2(_08660_),
    .B1(_04131_),
    .B2(_01049_),
    .Y(_01051_));
 sky130_fd_sc_hd__a31oi_4 _24213_ (.A1(net319),
    .A2(net161),
    .A3(net33),
    .B1(_01051_),
    .Y(_01053_));
 sky130_fd_sc_hd__nand2_1 _24214_ (.A(_08878_),
    .B(_01050_),
    .Y(_01054_));
 sky130_fd_sc_hd__o2111a_2 _24215_ (.A1(net166),
    .A2(net24),
    .B1(net33),
    .C1(net319),
    .D1(_01051_),
    .X(_01055_));
 sky130_fd_sc_hd__nand2_1 _24216_ (.A(net156),
    .B(_01051_),
    .Y(_01056_));
 sky130_fd_sc_hd__o22a_1 _24217_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_01051_),
    .B2(net156),
    .X(_01057_));
 sky130_fd_sc_hd__a22o_1 _24218_ (.A1(_08882_),
    .A2(_09298_),
    .B1(_01050_),
    .B2(_08878_),
    .X(_01058_));
 sky130_fd_sc_hd__o21ai_2 _24219_ (.A1(_01053_),
    .A2(_01055_),
    .B1(net146),
    .Y(_01059_));
 sky130_fd_sc_hd__o22ai_4 _24220_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_01053_),
    .B2(_01055_),
    .Y(_01060_));
 sky130_fd_sc_hd__nand3_2 _24221_ (.A(_01056_),
    .B(net146),
    .C(_01054_),
    .Y(_01061_));
 sky130_fd_sc_hd__a22oi_4 _24222_ (.A1(_00744_),
    .A2(_00748_),
    .B1(_01060_),
    .B2(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__o211ai_4 _24223_ (.A1(net146),
    .A2(_01053_),
    .B1(_01047_),
    .C1(_01059_),
    .Y(_01064_));
 sky130_fd_sc_hd__a2bb2oi_2 _24224_ (.A1_N(_00746_),
    .A2_N(_01046_),
    .B1(_01058_),
    .B2(_01059_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand3_2 _24225_ (.A(_01048_),
    .B(_01060_),
    .C(_01061_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand4_4 _24226_ (.A(net138),
    .B(net134),
    .C(_01064_),
    .D(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__o22ai_4 _24227_ (.A1(_10540_),
    .A2(net135),
    .B1(_01062_),
    .B2(_01065_),
    .Y(_01068_));
 sky130_fd_sc_hd__o21ai_1 _24228_ (.A1(_01062_),
    .A2(_01065_),
    .B1(net133),
    .Y(_01069_));
 sky130_fd_sc_hd__o211ai_1 _24229_ (.A1(_10540_),
    .A2(net135),
    .B1(_01064_),
    .C1(_01066_),
    .Y(_01070_));
 sky130_fd_sc_hd__o211a_1 _24230_ (.A1(_00754_),
    .A2(_00758_),
    .B1(_01067_),
    .C1(_01068_),
    .X(_01071_));
 sky130_fd_sc_hd__o211ai_4 _24231_ (.A1(_00754_),
    .A2(_00758_),
    .B1(_01067_),
    .C1(_01068_),
    .Y(_01072_));
 sky130_fd_sc_hd__a22oi_2 _24232_ (.A1(_00753_),
    .A2(_01044_),
    .B1(_01067_),
    .B2(_01068_),
    .Y(_01073_));
 sky130_fd_sc_hd__nand3_2 _24233_ (.A(_01045_),
    .B(_01069_),
    .C(_01070_),
    .Y(_01075_));
 sky130_fd_sc_hd__o311a_2 _24234_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_01072_),
    .C1(_01075_),
    .X(_01076_));
 sky130_fd_sc_hd__o211ai_4 _24235_ (.A1(_11042_),
    .A2(_11742_),
    .B1(_01072_),
    .C1(_01075_),
    .Y(_01077_));
 sky130_fd_sc_hd__a21oi_1 _24236_ (.A1(_01072_),
    .A2(_01075_),
    .B1(_12099_),
    .Y(_01078_));
 sky130_fd_sc_hd__o21ai_1 _24237_ (.A1(_01071_),
    .A2(_01073_),
    .B1(net132),
    .Y(_01079_));
 sky130_fd_sc_hd__o211ai_4 _24238_ (.A1(_00764_),
    .A2(_00768_),
    .B1(_01077_),
    .C1(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__o2bb2ai_4 _24239_ (.A1_N(_00766_),
    .A2_N(_01043_),
    .B1(_01076_),
    .B2(_01078_),
    .Y(_01081_));
 sky130_fd_sc_hd__o2111a_1 _24240_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_01080_),
    .D1(_01081_),
    .X(_01082_));
 sky130_fd_sc_hd__o2111ai_4 _24241_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_01080_),
    .D1(_01081_),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_1 _24242_ (.A1(_01080_),
    .A2(_01081_),
    .B1(_00736_),
    .Y(_01084_));
 sky130_fd_sc_hd__a22o_1 _24243_ (.A1(_00364_),
    .A2(_00367_),
    .B1(_01080_),
    .B2(_01081_),
    .X(_01086_));
 sky130_fd_sc_hd__o211a_1 _24244_ (.A1(_00775_),
    .A2(_00779_),
    .B1(_01083_),
    .C1(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__o211ai_4 _24245_ (.A1(_00775_),
    .A2(_00779_),
    .B1(_01083_),
    .C1(_01086_),
    .Y(_01088_));
 sky130_fd_sc_hd__o22ai_4 _24246_ (.A1(_00776_),
    .A2(_01042_),
    .B1(_01082_),
    .B2(_01084_),
    .Y(_01089_));
 sky130_fd_sc_hd__o21ai_2 _24247_ (.A1(_00810_),
    .A2(_00814_),
    .B1(_00860_),
    .Y(_01090_));
 sky130_fd_sc_hd__o211ai_2 _24248_ (.A1(net176),
    .A2(_07074_),
    .B1(net242),
    .C1(_07072_),
    .Y(_01091_));
 sky130_fd_sc_hd__or3_1 _24249_ (.A(net45),
    .B(_04212_),
    .C(_04102_),
    .X(_01092_));
 sky130_fd_sc_hd__o211ai_2 _24250_ (.A1(net176),
    .A2(_06759_),
    .B1(_05225_),
    .C1(net191),
    .Y(_01093_));
 sky130_fd_sc_hd__or3_1 _24251_ (.A(net46),
    .B(_04201_),
    .C(_04124_),
    .X(_01094_));
 sky130_fd_sc_hd__and4_1 _24252_ (.A(_01091_),
    .B(_01092_),
    .C(_01093_),
    .D(_01094_),
    .X(_01095_));
 sky130_fd_sc_hd__o2111ai_1 _24253_ (.A1(_04212_),
    .A2(_04989_),
    .B1(_01091_),
    .C1(_01093_),
    .D1(_01094_),
    .Y(_01097_));
 sky130_fd_sc_hd__a22oi_2 _24254_ (.A1(_01091_),
    .A2(_01092_),
    .B1(_01093_),
    .B2(_01094_),
    .Y(_01098_));
 sky130_fd_sc_hd__a32o_1 _24255_ (.A1(net197),
    .A2(_06452_),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net18),
    .X(_01099_));
 sky130_fd_sc_hd__o21bai_1 _24256_ (.A1(_01095_),
    .A2(_01098_),
    .B1_N(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2b_1 _24257_ (.A_N(_01098_),
    .B(_01099_),
    .Y(_01101_));
 sky130_fd_sc_hd__o21ai_4 _24258_ (.A1(_01095_),
    .A2(_01101_),
    .B1(_01100_),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_1 _24259_ (.A(_04245_),
    .B(_04483_),
    .Y(_01103_));
 sky130_fd_sc_hd__o211ai_1 _24260_ (.A1(net169),
    .A2(_07765_),
    .B1(_04480_),
    .C1(_07771_),
    .Y(_01104_));
 sky130_fd_sc_hd__a31oi_4 _24261_ (.A1(_07771_),
    .A2(_04480_),
    .A3(net166),
    .B1(_01103_),
    .Y(_01105_));
 sky130_fd_sc_hd__o211ai_4 _24262_ (.A1(net169),
    .A2(net268),
    .B1(_04267_),
    .C1(net164),
    .Y(_01106_));
 sky130_fd_sc_hd__or3b_2 _24263_ (.A(net41),
    .B(_04256_),
    .C_N(net40),
    .X(_01108_));
 sky130_fd_sc_hd__o221a_1 _24264_ (.A1(_04256_),
    .A2(_04270_),
    .B1(_04483_),
    .B2(_04245_),
    .C1(_01104_),
    .X(_01109_));
 sky130_fd_sc_hd__o211a_1 _24265_ (.A1(_04256_),
    .A2(_04270_),
    .B1(_01106_),
    .C1(_01105_),
    .X(_01110_));
 sky130_fd_sc_hd__o21ai_1 _24266_ (.A1(_04268_),
    .A2(_08209_),
    .B1(_01109_),
    .Y(_01111_));
 sky130_fd_sc_hd__a21oi_4 _24267_ (.A1(_01106_),
    .A2(_01108_),
    .B1(_01105_),
    .Y(_01112_));
 sky130_fd_sc_hd__a21o_1 _24268_ (.A1(_01106_),
    .A2(_01108_),
    .B1(_01105_),
    .X(_01113_));
 sky130_fd_sc_hd__o32a_2 _24269_ (.A1(_04896_),
    .A2(_07498_),
    .A3(_07502_),
    .B1(_04898_),
    .B2(_04223_),
    .X(_01114_));
 sky130_fd_sc_hd__a32o_1 _24270_ (.A1(_07499_),
    .A2(_07503_),
    .A3(_04895_),
    .B1(_04897_),
    .B2(net21),
    .X(_01115_));
 sky130_fd_sc_hd__o21ai_4 _24271_ (.A1(_01110_),
    .A2(_01112_),
    .B1(_01114_),
    .Y(_01116_));
 sky130_fd_sc_hd__a31o_1 _24272_ (.A1(_01105_),
    .A2(_01106_),
    .A3(_01108_),
    .B1(_01114_),
    .X(_01117_));
 sky130_fd_sc_hd__a211oi_4 _24273_ (.A1(_01109_),
    .A2(_01106_),
    .B1(_01114_),
    .C1(_01112_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand3_2 _24274_ (.A(_01111_),
    .B(_01113_),
    .C(_01115_),
    .Y(_01120_));
 sky130_fd_sc_hd__o31a_2 _24275_ (.A1(_00819_),
    .A2(_00820_),
    .A3(_00829_),
    .B1(_00831_),
    .X(_01121_));
 sky130_fd_sc_hd__a21oi_4 _24276_ (.A1(_01116_),
    .A2(_01120_),
    .B1(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand2_1 _24277_ (.A(_01121_),
    .B(_01116_),
    .Y(_01123_));
 sky130_fd_sc_hd__o211a_1 _24278_ (.A1(_01112_),
    .A2(_01117_),
    .B1(_01116_),
    .C1(_01121_),
    .X(_01124_));
 sky130_fd_sc_hd__o211ai_2 _24279_ (.A1(_01112_),
    .A2(_01117_),
    .B1(_01121_),
    .C1(_01116_),
    .Y(_01125_));
 sky130_fd_sc_hd__o21ai_2 _24280_ (.A1(_01122_),
    .A2(_01124_),
    .B1(_01102_),
    .Y(_01126_));
 sky130_fd_sc_hd__a31o_1 _24281_ (.A1(_01116_),
    .A2(_01120_),
    .A3(_01121_),
    .B1(_01102_),
    .X(_01127_));
 sky130_fd_sc_hd__o21ai_1 _24282_ (.A1(_01122_),
    .A2(_01127_),
    .B1(_01126_),
    .Y(_01128_));
 sky130_fd_sc_hd__o21a_1 _24283_ (.A1(_01122_),
    .A2(_01127_),
    .B1(_01126_),
    .X(_01130_));
 sky130_fd_sc_hd__o31ai_4 _24284_ (.A1(_00803_),
    .A2(_00356_),
    .A3(_00801_),
    .B1(_00406_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand2_2 _24285_ (.A(_00797_),
    .B(_00804_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_2 _24286_ (.A(net319),
    .B(_04218_),
    .Y(_01133_));
 sky130_fd_sc_hd__or3b_1 _24287_ (.A(net40),
    .B(net319),
    .C_N(net39),
    .X(_01134_));
 sky130_fd_sc_hd__a21oi_2 _24288_ (.A1(net150),
    .A2(_08668_),
    .B1(_04216_),
    .Y(_01135_));
 sky130_fd_sc_hd__o21ai_1 _24289_ (.A1(net159),
    .A2(_08666_),
    .B1(net281),
    .Y(_01136_));
 sky130_fd_sc_hd__o211ai_2 _24290_ (.A1(net169),
    .A2(net268),
    .B1(net319),
    .C1(_03704_),
    .Y(_01137_));
 sky130_fd_sc_hd__a31oi_4 _24291_ (.A1(net319),
    .A2(net161),
    .A3(_03704_),
    .B1(_00790_),
    .Y(_01138_));
 sky130_fd_sc_hd__o211ai_4 _24292_ (.A1(net319),
    .A2(_03737_),
    .B1(_01137_),
    .C1(_00795_),
    .Y(_01139_));
 sky130_fd_sc_hd__a22oi_4 _24293_ (.A1(_00795_),
    .A2(_01138_),
    .B1(_01136_),
    .B2(_01134_),
    .Y(_01141_));
 sky130_fd_sc_hd__a221oi_2 _24294_ (.A1(net25),
    .A2(_04217_),
    .B1(_08670_),
    .B2(net281),
    .C1(_01139_),
    .Y(_01142_));
 sky130_fd_sc_hd__a221o_1 _24295_ (.A1(net25),
    .A2(_04217_),
    .B1(_08670_),
    .B2(net281),
    .C1(_01139_),
    .X(_01143_));
 sky130_fd_sc_hd__o31ai_2 _24296_ (.A1(_01133_),
    .A2(_01135_),
    .A3(_01139_),
    .B1(_00355_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand3b_2 _24297_ (.A_N(_01141_),
    .B(_01143_),
    .C(_00355_),
    .Y(_01145_));
 sky130_fd_sc_hd__o22ai_4 _24298_ (.A1(_00037_),
    .A2(_00352_),
    .B1(_01141_),
    .B2(_01142_),
    .Y(_01146_));
 sky130_fd_sc_hd__o21a_1 _24299_ (.A1(_01141_),
    .A2(_01144_),
    .B1(_01146_),
    .X(_01147_));
 sky130_fd_sc_hd__a21o_1 _24300_ (.A1(_01145_),
    .A2(_01146_),
    .B1(_01132_),
    .X(_01148_));
 sky130_fd_sc_hd__o211ai_4 _24301_ (.A1(_01141_),
    .A2(_01144_),
    .B1(_01146_),
    .C1(_01132_),
    .Y(_01149_));
 sky130_fd_sc_hd__o211a_1 _24302_ (.A1(_01132_),
    .A2(_01147_),
    .B1(_00806_),
    .C1(_01131_),
    .X(_01150_));
 sky130_fd_sc_hd__o211ai_4 _24303_ (.A1(_01132_),
    .A2(_01147_),
    .B1(_00806_),
    .C1(_01131_),
    .Y(_01152_));
 sky130_fd_sc_hd__a22oi_2 _24304_ (.A1(_00806_),
    .A2(_01131_),
    .B1(_01148_),
    .B2(_01149_),
    .Y(_01153_));
 sky130_fd_sc_hd__a22o_1 _24305_ (.A1(_00806_),
    .A2(_01131_),
    .B1(_01148_),
    .B2(_01149_),
    .X(_01154_));
 sky130_fd_sc_hd__o21ai_1 _24306_ (.A1(_01150_),
    .A2(_01153_),
    .B1(_01130_),
    .Y(_01155_));
 sky130_fd_sc_hd__nand3_1 _24307_ (.A(_01154_),
    .B(_01128_),
    .C(_01152_),
    .Y(_01156_));
 sky130_fd_sc_hd__and3_2 _24308_ (.A(_01130_),
    .B(_01152_),
    .C(_01154_),
    .X(_01157_));
 sky130_fd_sc_hd__o2111ai_4 _24309_ (.A1(_01127_),
    .A2(_01122_),
    .B1(_01126_),
    .C1(_01152_),
    .D1(_01154_),
    .Y(_01158_));
 sky130_fd_sc_hd__o21ai_2 _24310_ (.A1(_01150_),
    .A2(_01153_),
    .B1(_01128_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _24311_ (.A(_01159_),
    .B(net130),
    .Y(_01160_));
 sky130_fd_sc_hd__nand3_4 _24312_ (.A(_01159_),
    .B(net130),
    .C(_01158_),
    .Y(_01161_));
 sky130_fd_sc_hd__o211ai_4 _24313_ (.A1(_00360_),
    .A2(_11741_),
    .B1(_01156_),
    .C1(_01155_),
    .Y(_01163_));
 sky130_fd_sc_hd__a22oi_4 _24314_ (.A1(_00817_),
    .A2(_00860_),
    .B1(_01161_),
    .B2(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__o2111a_1 _24315_ (.A1(_00810_),
    .A2(_00814_),
    .B1(_00860_),
    .C1(_01161_),
    .D1(_01163_),
    .X(_01165_));
 sky130_fd_sc_hd__o211a_1 _24316_ (.A1(_00816_),
    .A2(_00859_),
    .B1(_01161_),
    .C1(_01163_),
    .X(_01166_));
 sky130_fd_sc_hd__o221ai_4 _24317_ (.A1(_00816_),
    .A2(_00859_),
    .B1(_01160_),
    .B2(_01157_),
    .C1(_01163_),
    .Y(_01167_));
 sky130_fd_sc_hd__a21oi_2 _24318_ (.A1(_01161_),
    .A2(_01163_),
    .B1(_01090_),
    .Y(_01168_));
 sky130_fd_sc_hd__a21o_1 _24319_ (.A1(_01161_),
    .A2(_01163_),
    .B1(_01090_),
    .X(_01169_));
 sky130_fd_sc_hd__o211ai_4 _24320_ (.A1(_01166_),
    .A2(_01168_),
    .B1(_01088_),
    .C1(_01089_),
    .Y(_01170_));
 sky130_fd_sc_hd__o2bb2ai_2 _24321_ (.A1_N(_01088_),
    .A2_N(_01089_),
    .B1(_01164_),
    .B2(_01165_),
    .Y(_01171_));
 sky130_fd_sc_hd__o2bb2a_1 _24322_ (.A1_N(_01088_),
    .A2_N(_01089_),
    .B1(_01166_),
    .B2(_01168_),
    .X(_01172_));
 sky130_fd_sc_hd__o2bb2ai_2 _24323_ (.A1_N(_01088_),
    .A2_N(_01089_),
    .B1(_01166_),
    .B2(_01168_),
    .Y(_01174_));
 sky130_fd_sc_hd__o211ai_4 _24324_ (.A1(_01164_),
    .A2(_01165_),
    .B1(_01088_),
    .C1(_01089_),
    .Y(_01175_));
 sky130_fd_sc_hd__a31oi_4 _24325_ (.A1(_00783_),
    .A2(_00876_),
    .A3(_00879_),
    .B1(_00784_),
    .Y(_01176_));
 sky130_fd_sc_hd__a31o_1 _24326_ (.A1(_00783_),
    .A2(_00876_),
    .A3(_00879_),
    .B1(_00784_),
    .X(_01177_));
 sky130_fd_sc_hd__a21oi_4 _24327_ (.A1(_01174_),
    .A2(_01175_),
    .B1(_01176_),
    .Y(_01178_));
 sky130_fd_sc_hd__o2111ai_4 _24328_ (.A1(_00784_),
    .A2(_00880_),
    .B1(_01170_),
    .C1(_01171_),
    .D1(_00783_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand2_1 _24329_ (.A(_01176_),
    .B(_01175_),
    .Y(_01180_));
 sky130_fd_sc_hd__a21oi_1 _24330_ (.A1(_01170_),
    .A2(_01171_),
    .B1(_01177_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand3_4 _24331_ (.A(_01176_),
    .B(_01175_),
    .C(_01174_),
    .Y(_01182_));
 sky130_fd_sc_hd__o211ai_1 _24332_ (.A1(_01038_),
    .A2(_01032_),
    .B1(_01037_),
    .C1(_01182_),
    .Y(_01183_));
 sky130_fd_sc_hd__o2111ai_4 _24333_ (.A1(_01038_),
    .A2(_01032_),
    .B1(_01037_),
    .C1(_01179_),
    .D1(_01182_),
    .Y(_01185_));
 sky130_fd_sc_hd__o22ai_4 _24334_ (.A1(_01036_),
    .A2(_01039_),
    .B1(_01178_),
    .B2(_01181_),
    .Y(_01186_));
 sky130_fd_sc_hd__o21ai_1 _24335_ (.A1(_01178_),
    .A2(_01183_),
    .B1(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__o2111a_2 _24336_ (.A1(_00735_),
    .A2(_00887_),
    .B1(_00932_),
    .C1(_01185_),
    .D1(_01186_),
    .X(_01188_));
 sky130_fd_sc_hd__o2111ai_1 _24337_ (.A1(_00735_),
    .A2(_00887_),
    .B1(_00932_),
    .C1(_01185_),
    .D1(_01186_),
    .Y(_01189_));
 sky130_fd_sc_hd__a22oi_2 _24338_ (.A1(_00890_),
    .A2(_00932_),
    .B1(_01185_),
    .B2(_01186_),
    .Y(_01190_));
 sky130_fd_sc_hd__a22o_1 _24339_ (.A1(_00890_),
    .A2(_00932_),
    .B1(_01185_),
    .B2(_01186_),
    .X(_01191_));
 sky130_fd_sc_hd__a32o_1 _24340_ (.A1(_00717_),
    .A2(_00718_),
    .A3(_00722_),
    .B1(_00724_),
    .B2(_00585_),
    .X(_01192_));
 sky130_fd_sc_hd__nand3b_1 _24341_ (.A_N(_01192_),
    .B(_01191_),
    .C(_01189_),
    .Y(_01193_));
 sky130_fd_sc_hd__o21ai_1 _24342_ (.A1(_01188_),
    .A2(_01190_),
    .B1(_01192_),
    .Y(_01194_));
 sky130_fd_sc_hd__o21bai_2 _24343_ (.A1(_01188_),
    .A2(_01190_),
    .B1_N(_01192_),
    .Y(_01196_));
 sky130_fd_sc_hd__a21boi_2 _24344_ (.A1(_00933_),
    .A2(_01187_),
    .B1_N(_01192_),
    .Y(_01197_));
 sky130_fd_sc_hd__nand3_1 _24345_ (.A(_01189_),
    .B(_01191_),
    .C(_01192_),
    .Y(_01198_));
 sky130_fd_sc_hd__o211ai_4 _24346_ (.A1(_00898_),
    .A2(_00906_),
    .B1(_01193_),
    .C1(_01194_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand3_4 _24347_ (.A(_01196_),
    .B(_01198_),
    .C(_00907_),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _24348_ (.A(_01199_),
    .B(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__a21o_1 _24349_ (.A1(_01199_),
    .A2(_01200_),
    .B1(_00929_),
    .X(_01202_));
 sky130_fd_sc_hd__and3_1 _24350_ (.A(_00929_),
    .B(_01199_),
    .C(_01200_),
    .X(_01203_));
 sky130_fd_sc_hd__o211ai_4 _24351_ (.A1(_00710_),
    .A2(_00714_),
    .B1(_01199_),
    .C1(_01200_),
    .Y(_01204_));
 sky130_fd_sc_hd__o211a_1 _24352_ (.A1(_00573_),
    .A2(_00543_),
    .B1(_00569_),
    .C1(_00912_),
    .X(_01205_));
 sky130_fd_sc_hd__o21ai_1 _24353_ (.A1(_00632_),
    .A2(_00913_),
    .B1(_00912_),
    .Y(_01207_));
 sky130_fd_sc_hd__a21oi_1 _24354_ (.A1(_01202_),
    .A2(_01204_),
    .B1(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__o2bb2ai_1 _24355_ (.A1_N(_01202_),
    .A2_N(_01204_),
    .B1(_01205_),
    .B2(_00913_),
    .Y(_01209_));
 sky130_fd_sc_hd__a22oi_1 _24356_ (.A1(_01201_),
    .A2(_00930_),
    .B1(_00916_),
    .B2(_00912_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_1 _24357_ (.A(_01207_),
    .B(_01202_),
    .Y(_01211_));
 sky130_fd_sc_hd__a21oi_2 _24358_ (.A1(_01204_),
    .A2(_01210_),
    .B1(_01208_),
    .Y(_01212_));
 sky130_fd_sc_hd__o21ai_1 _24359_ (.A1(_00925_),
    .A2(_00928_),
    .B1(_00923_),
    .Y(_01213_));
 sky130_fd_sc_hd__xor2_1 _24360_ (.A(_01212_),
    .B(_01213_),
    .X(net106));
 sky130_fd_sc_hd__a31o_1 _24361_ (.A1(_00937_),
    .A2(_00962_),
    .A3(_00963_),
    .B1(_00969_),
    .X(_01214_));
 sky130_fd_sc_hd__inv_2 _24362_ (.A(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__a21o_1 _24363_ (.A1(_01031_),
    .A2(_01035_),
    .B1(_01032_),
    .X(_01217_));
 sky130_fd_sc_hd__o22ai_2 _24364_ (.A1(_01172_),
    .A2(_01180_),
    .B1(_01178_),
    .B2(_01040_),
    .Y(_01218_));
 sky130_fd_sc_hd__a21boi_2 _24365_ (.A1(_01081_),
    .A2(_00736_),
    .B1_N(_01080_),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_1 _24366_ (.A(_01080_),
    .B(_01083_),
    .Y(_01220_));
 sky130_fd_sc_hd__o21ai_1 _24367_ (.A1(net132),
    .A2(_01073_),
    .B1(_01072_),
    .Y(_01221_));
 sky130_fd_sc_hd__or3_2 _24368_ (.A(net57),
    .B(_04266_),
    .C(_04069_),
    .X(_01222_));
 sky130_fd_sc_hd__o31ai_2 _24369_ (.A1(net262),
    .A2(net244),
    .A3(_04407_),
    .B1(_08657_),
    .Y(_01223_));
 sky130_fd_sc_hd__nand4_2 _24370_ (.A(_04266_),
    .B(net225),
    .C(net57),
    .D(_04409_),
    .Y(_01224_));
 sky130_fd_sc_hd__o22ai_4 _24371_ (.A1(_04069_),
    .A2(_08660_),
    .B1(_04410_),
    .B2(_01223_),
    .Y(_01225_));
 sky130_fd_sc_hd__a21oi_4 _24372_ (.A1(_08876_),
    .A2(net319),
    .B1(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__nand3_1 _24373_ (.A(_08878_),
    .B(_01222_),
    .C(_01224_),
    .Y(_01228_));
 sky130_fd_sc_hd__a21oi_2 _24374_ (.A1(_01222_),
    .A2(_01224_),
    .B1(_08878_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand3_2 _24375_ (.A(_01225_),
    .B(net159),
    .C(net33),
    .Y(_01230_));
 sky130_fd_sc_hd__o22a_1 _24376_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_01225_),
    .B2(net156),
    .X(_01231_));
 sky130_fd_sc_hd__a31o_1 _24377_ (.A1(_08878_),
    .A2(_01222_),
    .A3(_01224_),
    .B1(net146),
    .X(_01232_));
 sky130_fd_sc_hd__a21o_1 _24378_ (.A1(_01228_),
    .A2(_01230_),
    .B1(_09300_),
    .X(_01233_));
 sky130_fd_sc_hd__o22ai_2 _24379_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_01226_),
    .B2(_01229_),
    .Y(_01234_));
 sky130_fd_sc_hd__o2111ai_4 _24380_ (.A1(_04495_),
    .A2(net150),
    .B1(_08882_),
    .C1(_01228_),
    .D1(_01230_),
    .Y(_01235_));
 sky130_fd_sc_hd__a21oi_1 _24381_ (.A1(_09300_),
    .A2(_01054_),
    .B1(_01055_),
    .Y(_01236_));
 sky130_fd_sc_hd__o211ai_1 _24382_ (.A1(_01050_),
    .A2(_08878_),
    .B1(_01235_),
    .C1(_01234_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand3_2 _24383_ (.A(_01234_),
    .B(_01235_),
    .C(_01236_),
    .Y(_01239_));
 sky130_fd_sc_hd__a21oi_1 _24384_ (.A1(_01234_),
    .A2(_01235_),
    .B1(_01236_),
    .Y(_01240_));
 sky130_fd_sc_hd__o221ai_4 _24385_ (.A1(_01055_),
    .A2(_01057_),
    .B1(_01226_),
    .B2(net146),
    .C1(_01233_),
    .Y(_01241_));
 sky130_fd_sc_hd__a21oi_1 _24386_ (.A1(_01239_),
    .A2(_01241_),
    .B1(net133),
    .Y(_01242_));
 sky130_fd_sc_hd__a22o_1 _24387_ (.A1(net138),
    .A2(net134),
    .B1(_01239_),
    .B2(_01241_),
    .X(_01243_));
 sky130_fd_sc_hd__o211a_2 _24388_ (.A1(_01057_),
    .A2(_01237_),
    .B1(_01241_),
    .C1(net133),
    .X(_01244_));
 sky130_fd_sc_hd__nand3_2 _24389_ (.A(net133),
    .B(_01239_),
    .C(_01241_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand2_1 _24390_ (.A(_01243_),
    .B(_01245_),
    .Y(_01246_));
 sky130_fd_sc_hd__o21ai_1 _24391_ (.A1(_10546_),
    .A2(_01065_),
    .B1(_01064_),
    .Y(_01247_));
 sky130_fd_sc_hd__a32o_1 _24392_ (.A1(_01048_),
    .A2(_01060_),
    .A3(_01061_),
    .B1(_01064_),
    .B2(_10546_),
    .X(_01248_));
 sky130_fd_sc_hd__a21oi_1 _24393_ (.A1(_01243_),
    .A2(_01245_),
    .B1(_01247_),
    .Y(_01250_));
 sky130_fd_sc_hd__o21ai_2 _24394_ (.A1(_01242_),
    .A2(_01244_),
    .B1(_01248_),
    .Y(_01251_));
 sky130_fd_sc_hd__nand2_1 _24395_ (.A(_01243_),
    .B(_01247_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor3_2 _24396_ (.A(_01242_),
    .B(_01248_),
    .C(_01244_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand3_1 _24397_ (.A(_01243_),
    .B(_01245_),
    .C(_01247_),
    .Y(_01254_));
 sky130_fd_sc_hd__a21oi_1 _24398_ (.A1(_01251_),
    .A2(_01254_),
    .B1(_12099_),
    .Y(_01255_));
 sky130_fd_sc_hd__o21ai_2 _24399_ (.A1(_01250_),
    .A2(_01253_),
    .B1(net132),
    .Y(_01256_));
 sky130_fd_sc_hd__a21oi_2 _24400_ (.A1(_01246_),
    .A2(_01248_),
    .B1(net132),
    .Y(_01257_));
 sky130_fd_sc_hd__o221ai_4 _24401_ (.A1(_11042_),
    .A2(_11742_),
    .B1(_01244_),
    .B2(_01252_),
    .C1(_01251_),
    .Y(_01258_));
 sky130_fd_sc_hd__a221oi_2 _24402_ (.A1(_01072_),
    .A2(_01077_),
    .B1(_01254_),
    .B2(_01257_),
    .C1(_01255_),
    .Y(_01259_));
 sky130_fd_sc_hd__o211ai_4 _24403_ (.A1(_01071_),
    .A2(_01076_),
    .B1(_01256_),
    .C1(_01258_),
    .Y(_01261_));
 sky130_fd_sc_hd__a21oi_2 _24404_ (.A1(_01256_),
    .A2(_01258_),
    .B1(_01221_),
    .Y(_01262_));
 sky130_fd_sc_hd__a21o_1 _24405_ (.A1(_01256_),
    .A2(_01258_),
    .B1(_01221_),
    .X(_01263_));
 sky130_fd_sc_hd__o22ai_2 _24406_ (.A1(net130),
    .A2(_00366_),
    .B1(_01259_),
    .B2(_01262_),
    .Y(_01264_));
 sky130_fd_sc_hd__o2111ai_4 _24407_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_01261_),
    .D1(_01263_),
    .Y(_01265_));
 sky130_fd_sc_hd__o211ai_2 _24408_ (.A1(net130),
    .A2(_00366_),
    .B1(_01261_),
    .C1(_01263_),
    .Y(_01266_));
 sky130_fd_sc_hd__o21ai_2 _24409_ (.A1(_01259_),
    .A2(_01262_),
    .B1(_00736_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_1 _24410_ (.A(_01264_),
    .B(_01265_),
    .Y(_01268_));
 sky130_fd_sc_hd__and3_1 _24411_ (.A(_01220_),
    .B(_01264_),
    .C(_01265_),
    .X(_01269_));
 sky130_fd_sc_hd__nand3_2 _24412_ (.A(_01220_),
    .B(_01264_),
    .C(_01265_),
    .Y(_01270_));
 sky130_fd_sc_hd__and3_1 _24413_ (.A(_01267_),
    .B(_01219_),
    .C(_01266_),
    .X(_01272_));
 sky130_fd_sc_hd__nand3_4 _24414_ (.A(_01267_),
    .B(_01219_),
    .C(_01266_),
    .Y(_01273_));
 sky130_fd_sc_hd__a32o_2 _24415_ (.A1(_00806_),
    .A2(_01131_),
    .A3(_01148_),
    .B1(_01154_),
    .B2(_01130_),
    .X(_01274_));
 sky130_fd_sc_hd__a21oi_1 _24416_ (.A1(_01111_),
    .A2(_01115_),
    .B1(_01112_),
    .Y(_01275_));
 sky130_fd_sc_hd__and3_1 _24417_ (.A(_04102_),
    .B(net22),
    .C(net42),
    .X(_01276_));
 sky130_fd_sc_hd__o311a_1 _24418_ (.A1(net233),
    .A2(_05927_),
    .A3(_07767_),
    .B1(_07771_),
    .C1(_04895_),
    .X(_01277_));
 sky130_fd_sc_hd__a31oi_2 _24419_ (.A1(_07771_),
    .A2(_04895_),
    .A3(net166),
    .B1(_01276_),
    .Y(_01278_));
 sky130_fd_sc_hd__a31o_1 _24420_ (.A1(_07771_),
    .A2(_04895_),
    .A3(net166),
    .B1(_01276_),
    .X(_01279_));
 sky130_fd_sc_hd__o211ai_2 _24421_ (.A1(net169),
    .A2(net268),
    .B1(_04480_),
    .C1(net164),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_1 _24422_ (.A(_04256_),
    .B(_04483_),
    .Y(_01281_));
 sky130_fd_sc_hd__or3b_1 _24423_ (.A(net42),
    .B(_04256_),
    .C_N(net41),
    .X(_01283_));
 sky130_fd_sc_hd__a31oi_4 _24424_ (.A1(net164),
    .A2(net161),
    .A3(_04480_),
    .B1(_01281_),
    .Y(_01284_));
 sky130_fd_sc_hd__a21oi_1 _24425_ (.A1(net150),
    .A2(_08668_),
    .B1(_04268_),
    .Y(_01285_));
 sky130_fd_sc_hd__o21ai_2 _24426_ (.A1(_08664_),
    .A2(_08666_),
    .B1(_04267_),
    .Y(_01286_));
 sky130_fd_sc_hd__nor2_1 _24427_ (.A(net319),
    .B(_04270_),
    .Y(_01287_));
 sky130_fd_sc_hd__or3b_4 _24428_ (.A(net41),
    .B(net319),
    .C_N(net40),
    .X(_01288_));
 sky130_fd_sc_hd__a21oi_1 _24429_ (.A1(_08670_),
    .A2(_04267_),
    .B1(_01287_),
    .Y(_01289_));
 sky130_fd_sc_hd__a22oi_4 _24430_ (.A1(_01280_),
    .A2(_01283_),
    .B1(_01286_),
    .B2(_01288_),
    .Y(_01290_));
 sky130_fd_sc_hd__o21bai_1 _24431_ (.A1(_01285_),
    .A2(_01287_),
    .B1_N(_01284_),
    .Y(_01291_));
 sky130_fd_sc_hd__o211a_1 _24432_ (.A1(net319),
    .A2(_04270_),
    .B1(_01284_),
    .C1(_01286_),
    .X(_01292_));
 sky130_fd_sc_hd__o211ai_2 _24433_ (.A1(net319),
    .A2(_04270_),
    .B1(_01284_),
    .C1(_01286_),
    .Y(_01294_));
 sky130_fd_sc_hd__o21ai_1 _24434_ (.A1(_01290_),
    .A2(_01292_),
    .B1(_01278_),
    .Y(_01295_));
 sky130_fd_sc_hd__o21ai_1 _24435_ (.A1(_01284_),
    .A2(_01289_),
    .B1(_01279_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand3_1 _24436_ (.A(_01291_),
    .B(_01294_),
    .C(_01278_),
    .Y(_01297_));
 sky130_fd_sc_hd__o22ai_2 _24437_ (.A1(_01276_),
    .A2(_01277_),
    .B1(_01290_),
    .B2(_01292_),
    .Y(_01298_));
 sky130_fd_sc_hd__a2bb2oi_1 _24438_ (.A1_N(_01112_),
    .A2_N(_01119_),
    .B1(_01297_),
    .B2(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__o221ai_4 _24439_ (.A1(_01112_),
    .A2(_01119_),
    .B1(_01292_),
    .B2(_01296_),
    .C1(_01295_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand3_2 _24440_ (.A(_01298_),
    .B(_01275_),
    .C(_01297_),
    .Y(_01301_));
 sky130_fd_sc_hd__nor2_1 _24441_ (.A(_04201_),
    .B(_05465_),
    .Y(_01302_));
 sky130_fd_sc_hd__o311a_1 _24442_ (.A1(net244),
    .A2(net241),
    .A3(_06759_),
    .B1(_05462_),
    .C1(net191),
    .X(_01303_));
 sky130_fd_sc_hd__o32a_1 _24443_ (.A1(_05463_),
    .A2(_06756_),
    .A3(net190),
    .B1(_05465_),
    .B2(_04201_),
    .X(_01305_));
 sky130_fd_sc_hd__nor2_1 _24444_ (.A(_04212_),
    .B(_05229_),
    .Y(_01306_));
 sky130_fd_sc_hd__a31oi_2 _24445_ (.A1(_07072_),
    .A2(net170),
    .A3(_05225_),
    .B1(_01306_),
    .Y(_01307_));
 sky130_fd_sc_hd__and3_1 _24446_ (.A(_04124_),
    .B(net21),
    .C(net43),
    .X(_01308_));
 sky130_fd_sc_hd__a31oi_4 _24447_ (.A1(_07499_),
    .A2(_07503_),
    .A3(net242),
    .B1(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__nor2_1 _24448_ (.A(_01307_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__o221a_1 _24449_ (.A1(_04212_),
    .A2(_05229_),
    .B1(_07079_),
    .B2(_05226_),
    .C1(_01309_),
    .X(_01311_));
 sky130_fd_sc_hd__nand2_1 _24450_ (.A(_01307_),
    .B(_01309_),
    .Y(_01312_));
 sky130_fd_sc_hd__o22ai_1 _24451_ (.A1(_01302_),
    .A2(_01303_),
    .B1(_01310_),
    .B2(_01311_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand3b_1 _24452_ (.A_N(_01310_),
    .B(_01312_),
    .C(_01305_),
    .Y(_01314_));
 sky130_fd_sc_hd__nand2_2 _24453_ (.A(_01313_),
    .B(_01314_),
    .Y(_01316_));
 sky130_fd_sc_hd__a21o_1 _24454_ (.A1(_01300_),
    .A2(_01301_),
    .B1(_01316_),
    .X(_01317_));
 sky130_fd_sc_hd__nand3_4 _24455_ (.A(_01300_),
    .B(_01301_),
    .C(_01316_),
    .Y(_01318_));
 sky130_fd_sc_hd__a31oi_4 _24456_ (.A1(net319),
    .A2(net161),
    .A3(net281),
    .B1(_01133_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand2_1 _24457_ (.A(_01139_),
    .B(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand3b_2 _24458_ (.A_N(_01319_),
    .B(_01138_),
    .C(_00795_),
    .Y(_01321_));
 sky130_fd_sc_hd__o2111ai_4 _24459_ (.A1(_03714_),
    .A2(net150),
    .B1(_00791_),
    .C1(_00795_),
    .D1(_01319_),
    .Y(_01322_));
 sky130_fd_sc_hd__a31o_1 _24460_ (.A1(_00791_),
    .A2(_00795_),
    .A3(_01137_),
    .B1(_01319_),
    .X(_01323_));
 sky130_fd_sc_hd__a2bb2o_4 _24461_ (.A1_N(_00037_),
    .A2_N(_00352_),
    .B1(_01322_),
    .B2(_01323_),
    .X(_01324_));
 sky130_fd_sc_hd__nand4_4 _24462_ (.A(_00038_),
    .B(_00353_),
    .C(_01322_),
    .D(_01323_),
    .Y(_01325_));
 sky130_fd_sc_hd__a21oi_1 _24463_ (.A1(_01324_),
    .A2(_01325_),
    .B1(_01141_),
    .Y(_01327_));
 sky130_fd_sc_hd__and3_2 _24464_ (.A(_01324_),
    .B(_01325_),
    .C(_01141_),
    .X(_01328_));
 sky130_fd_sc_hd__o2111ai_4 _24465_ (.A1(_01133_),
    .A2(_01135_),
    .B1(_01139_),
    .C1(_01324_),
    .D1(_01325_),
    .Y(_01329_));
 sky130_fd_sc_hd__a21oi_4 _24466_ (.A1(_01145_),
    .A2(_01149_),
    .B1(_01327_),
    .Y(_01330_));
 sky130_fd_sc_hd__and4_2 _24467_ (.A(_00356_),
    .B(_00795_),
    .C(_01320_),
    .D(_01321_),
    .X(_01331_));
 sky130_fd_sc_hd__nand4_4 _24468_ (.A(_00356_),
    .B(_00795_),
    .C(_01320_),
    .D(_01321_),
    .Y(_01332_));
 sky130_fd_sc_hd__a31o_1 _24469_ (.A1(_01141_),
    .A2(_01324_),
    .A3(_01325_),
    .B1(_01331_),
    .X(_01333_));
 sky130_fd_sc_hd__o21a_1 _24470_ (.A1(_00796_),
    .A2(_01324_),
    .B1(_01329_),
    .X(_01334_));
 sky130_fd_sc_hd__a211o_1 _24471_ (.A1(_01317_),
    .A2(_01318_),
    .B1(_01330_),
    .C1(_01333_),
    .X(_01335_));
 sky130_fd_sc_hd__o211ai_2 _24472_ (.A1(_01330_),
    .A2(_01333_),
    .B1(_01317_),
    .C1(_01318_),
    .Y(_01336_));
 sky130_fd_sc_hd__and3_2 _24473_ (.A(_01317_),
    .B(_01318_),
    .C(_01334_),
    .X(_01338_));
 sky130_fd_sc_hd__nand4_2 _24474_ (.A(_01317_),
    .B(_01318_),
    .C(_01329_),
    .D(_01332_),
    .Y(_01339_));
 sky130_fd_sc_hd__o2bb2ai_1 _24475_ (.A1_N(_01317_),
    .A2_N(_01318_),
    .B1(_01330_),
    .B2(_01333_),
    .Y(_01340_));
 sky130_fd_sc_hd__o2111ai_4 _24476_ (.A1(_01330_),
    .A2(_01339_),
    .B1(_01340_),
    .C1(_00361_),
    .D1(_11740_),
    .Y(_01341_));
 sky130_fd_sc_hd__inv_2 _24477_ (.A(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__o211ai_4 _24478_ (.A1(_00360_),
    .A2(_11741_),
    .B1(_01336_),
    .C1(_01335_),
    .Y(_01343_));
 sky130_fd_sc_hd__a21boi_2 _24479_ (.A1(_01341_),
    .A2(_01343_),
    .B1_N(_01274_),
    .Y(_01344_));
 sky130_fd_sc_hd__o2111a_2 _24480_ (.A1(_01128_),
    .A2(_01153_),
    .B1(_01341_),
    .C1(_01343_),
    .D1(_01152_),
    .X(_01345_));
 sky130_fd_sc_hd__and2_1 _24481_ (.A(_01274_),
    .B(_01343_),
    .X(_01346_));
 sky130_fd_sc_hd__and3_1 _24482_ (.A(_01274_),
    .B(_01341_),
    .C(_01343_),
    .X(_01347_));
 sky130_fd_sc_hd__a21oi_2 _24483_ (.A1(_01341_),
    .A2(_01343_),
    .B1(_01274_),
    .Y(_01349_));
 sky130_fd_sc_hd__o211ai_2 _24484_ (.A1(_01347_),
    .A2(_01349_),
    .B1(_01270_),
    .C1(_01273_),
    .Y(_01350_));
 sky130_fd_sc_hd__o2bb2ai_2 _24485_ (.A1_N(_01270_),
    .A2_N(_01273_),
    .B1(_01344_),
    .B2(_01345_),
    .Y(_01351_));
 sky130_fd_sc_hd__o2bb2ai_2 _24486_ (.A1_N(_01270_),
    .A2_N(_01273_),
    .B1(_01347_),
    .B2(_01349_),
    .Y(_01352_));
 sky130_fd_sc_hd__o211ai_2 _24487_ (.A1(_01344_),
    .A2(_01345_),
    .B1(_01270_),
    .C1(_01273_),
    .Y(_01353_));
 sky130_fd_sc_hd__a31o_1 _24488_ (.A1(_01089_),
    .A2(_01167_),
    .A3(_01169_),
    .B1(_01087_),
    .X(_01354_));
 sky130_fd_sc_hd__a31oi_2 _24489_ (.A1(_01089_),
    .A2(_01167_),
    .A3(_01169_),
    .B1(_01087_),
    .Y(_01355_));
 sky130_fd_sc_hd__and3_1 _24490_ (.A(_01350_),
    .B(_01351_),
    .C(_01355_),
    .X(_01356_));
 sky130_fd_sc_hd__nand3_4 _24491_ (.A(_01350_),
    .B(_01351_),
    .C(_01355_),
    .Y(_01357_));
 sky130_fd_sc_hd__and3_1 _24492_ (.A(_01354_),
    .B(_01353_),
    .C(_01352_),
    .X(_01358_));
 sky130_fd_sc_hd__nand3_4 _24493_ (.A(_01354_),
    .B(_01353_),
    .C(_01352_),
    .Y(_01360_));
 sky130_fd_sc_hd__a21oi_2 _24494_ (.A1(_00983_),
    .A2(_00990_),
    .B1(_00991_),
    .Y(_01361_));
 sky130_fd_sc_hd__a21o_1 _24495_ (.A1(_01097_),
    .A2(_01099_),
    .B1(_01098_),
    .X(_01362_));
 sky130_fd_sc_hd__a32o_1 _24496_ (.A1(net176),
    .A2(_05933_),
    .A3(net273),
    .B1(_06326_),
    .B2(net16),
    .X(_01363_));
 sky130_fd_sc_hd__or3b_2 _24497_ (.A(net49),
    .B(_04168_),
    .C_N(net48),
    .X(_01364_));
 sky130_fd_sc_hd__o211ai_4 _24498_ (.A1(_05927_),
    .A2(_06220_),
    .B1(net274),
    .C1(net202),
    .Y(_01365_));
 sky130_fd_sc_hd__or3b_4 _24499_ (.A(net48),
    .B(_04179_),
    .C_N(net47),
    .X(_01366_));
 sky130_fd_sc_hd__o211ai_4 _24500_ (.A1(net176),
    .A2(_06451_),
    .B1(_05762_),
    .C1(net197),
    .Y(_01367_));
 sky130_fd_sc_hd__o2111a_1 _24501_ (.A1(_04168_),
    .A2(_06030_),
    .B1(_01365_),
    .C1(_01366_),
    .D1(_01367_),
    .X(_01368_));
 sky130_fd_sc_hd__o2111ai_4 _24502_ (.A1(_04168_),
    .A2(_06030_),
    .B1(_01365_),
    .C1(_01366_),
    .D1(_01367_),
    .Y(_01369_));
 sky130_fd_sc_hd__a22oi_4 _24503_ (.A1(_01364_),
    .A2(_01365_),
    .B1(_01366_),
    .B2(_01367_),
    .Y(_01371_));
 sky130_fd_sc_hd__a22o_1 _24504_ (.A1(_01364_),
    .A2(_01365_),
    .B1(_01366_),
    .B2(_01367_),
    .X(_01372_));
 sky130_fd_sc_hd__o21bai_4 _24505_ (.A1(_01368_),
    .A2(_01371_),
    .B1_N(_01363_),
    .Y(_01373_));
 sky130_fd_sc_hd__and3_1 _24506_ (.A(_01363_),
    .B(_01369_),
    .C(_01372_),
    .X(_01374_));
 sky130_fd_sc_hd__nand3_2 _24507_ (.A(_01363_),
    .B(_01369_),
    .C(_01372_),
    .Y(_01375_));
 sky130_fd_sc_hd__a21oi_4 _24508_ (.A1(_01373_),
    .A2(_01375_),
    .B1(_01362_),
    .Y(_01376_));
 sky130_fd_sc_hd__and3_1 _24509_ (.A(_01362_),
    .B(_01373_),
    .C(_01375_),
    .X(_01377_));
 sky130_fd_sc_hd__nand3_1 _24510_ (.A(_01362_),
    .B(_01373_),
    .C(_01375_),
    .Y(_01378_));
 sky130_fd_sc_hd__a31o_1 _24511_ (.A1(_01362_),
    .A2(_01373_),
    .A3(_01375_),
    .B1(_01361_),
    .X(_01379_));
 sky130_fd_sc_hd__o21ai_1 _24512_ (.A1(_01376_),
    .A2(_01377_),
    .B1(_01361_),
    .Y(_01380_));
 sky130_fd_sc_hd__nand3b_1 _24513_ (.A_N(_01376_),
    .B(_01378_),
    .C(_01361_),
    .Y(_01382_));
 sky130_fd_sc_hd__o22ai_2 _24514_ (.A1(_00991_),
    .A2(_00993_),
    .B1(_01376_),
    .B2(_01377_),
    .Y(_01383_));
 sky130_fd_sc_hd__o22ai_2 _24515_ (.A1(_01119_),
    .A2(_01123_),
    .B1(_01102_),
    .B2(_01122_),
    .Y(_01384_));
 sky130_fd_sc_hd__o2111ai_4 _24516_ (.A1(_01102_),
    .A2(_01122_),
    .B1(_01125_),
    .C1(_01382_),
    .D1(_01383_),
    .Y(_01385_));
 sky130_fd_sc_hd__o211ai_4 _24517_ (.A1(_01376_),
    .A2(_01379_),
    .B1(_01380_),
    .C1(_01384_),
    .Y(_01386_));
 sky130_fd_sc_hd__inv_2 _24518_ (.A(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__a21o_1 _24519_ (.A1(_00978_),
    .A2(_01000_),
    .B1(_00999_),
    .X(_01388_));
 sky130_fd_sc_hd__a21oi_2 _24520_ (.A1(_01385_),
    .A2(_01386_),
    .B1(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__a21o_1 _24521_ (.A1(_01385_),
    .A2(_01386_),
    .B1(_01388_),
    .X(_01390_));
 sky130_fd_sc_hd__o211a_2 _24522_ (.A1(_00999_),
    .A2(_01001_),
    .B1(_01385_),
    .C1(_01386_),
    .X(_01391_));
 sky130_fd_sc_hd__o211ai_4 _24523_ (.A1(_00999_),
    .A2(_01001_),
    .B1(_01385_),
    .C1(_01386_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand3_4 _24524_ (.A(_01015_),
    .B(_01390_),
    .C(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__o22ai_4 _24525_ (.A1(_01011_),
    .A2(_01013_),
    .B1(_01389_),
    .B2(_01391_),
    .Y(_01395_));
 sky130_fd_sc_hd__o2bb2a_2 _24526_ (.A1_N(_04560_),
    .A2_N(net238),
    .B1(_08007_),
    .B2(_04080_),
    .X(_01396_));
 sky130_fd_sc_hd__a32o_1 _24527_ (.A1(net220),
    .A2(net186),
    .A3(net238),
    .B1(_08006_),
    .B2(net10),
    .X(_01397_));
 sky130_fd_sc_hd__a2bb2o_2 _24528_ (.A1_N(_00958_),
    .A2_N(_00954_),
    .B1(_00938_),
    .B2(_00961_),
    .X(_01398_));
 sky130_fd_sc_hd__a32o_1 _24529_ (.A1(net184),
    .A2(net213),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net11),
    .X(_01399_));
 sky130_fd_sc_hd__a32o_1 _24530_ (.A1(net209),
    .A2(_05074_),
    .A3(net239),
    .B1(_07308_),
    .B2(net13),
    .X(_01400_));
 sky130_fd_sc_hd__or3b_1 _24531_ (.A(_04135_),
    .B(net52),
    .C_N(net51),
    .X(_01401_));
 sky130_fd_sc_hd__nand3_4 _24532_ (.A(_05290_),
    .B(_05292_),
    .C(net269),
    .Y(_01402_));
 sky130_fd_sc_hd__or3_2 _24533_ (.A(net51),
    .B(_04190_),
    .C(_04146_),
    .X(_01404_));
 sky130_fd_sc_hd__o211ai_4 _24534_ (.A1(net184),
    .A2(_05551_),
    .B1(net240),
    .C1(net178),
    .Y(_01405_));
 sky130_fd_sc_hd__a22oi_4 _24535_ (.A1(_01401_),
    .A2(_01402_),
    .B1(_01404_),
    .B2(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__a22o_1 _24536_ (.A1(_01401_),
    .A2(_01402_),
    .B1(_01404_),
    .B2(_01405_),
    .X(_01407_));
 sky130_fd_sc_hd__o2111a_1 _24537_ (.A1(_04135_),
    .A2(_07226_),
    .B1(_01402_),
    .C1(_01404_),
    .D1(_01405_),
    .X(_01408_));
 sky130_fd_sc_hd__o2111ai_4 _24538_ (.A1(_04135_),
    .A2(_07226_),
    .B1(_01402_),
    .C1(_01404_),
    .D1(_01405_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand3_1 _24539_ (.A(_01400_),
    .B(_01407_),
    .C(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__o21bai_1 _24540_ (.A1(_01406_),
    .A2(_01408_),
    .B1_N(_01400_),
    .Y(_01411_));
 sky130_fd_sc_hd__o21ai_1 _24541_ (.A1(_01406_),
    .A2(_01408_),
    .B1(_01400_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand3b_1 _24542_ (.A_N(_01400_),
    .B(_01407_),
    .C(_01409_),
    .Y(_01413_));
 sky130_fd_sc_hd__nand3_1 _24543_ (.A(_01412_),
    .B(_01413_),
    .C(_00952_),
    .Y(_01415_));
 sky130_fd_sc_hd__nand3b_2 _24544_ (.A_N(_00952_),
    .B(_01410_),
    .C(_01411_),
    .Y(_01416_));
 sky130_fd_sc_hd__a21o_1 _24545_ (.A1(_01415_),
    .A2(_01416_),
    .B1(_01399_),
    .X(_01417_));
 sky130_fd_sc_hd__nand3_2 _24546_ (.A(_01399_),
    .B(_01415_),
    .C(_01416_),
    .Y(_01418_));
 sky130_fd_sc_hd__a21o_1 _24547_ (.A1(_01417_),
    .A2(_01418_),
    .B1(_01398_),
    .X(_01419_));
 sky130_fd_sc_hd__and3_1 _24548_ (.A(_01398_),
    .B(_01417_),
    .C(_01418_),
    .X(_01420_));
 sky130_fd_sc_hd__nand3_4 _24549_ (.A(_01398_),
    .B(_01417_),
    .C(_01418_),
    .Y(_01421_));
 sky130_fd_sc_hd__a21oi_1 _24550_ (.A1(_01419_),
    .A2(_01421_),
    .B1(_01397_),
    .Y(_01422_));
 sky130_fd_sc_hd__nand3_2 _24551_ (.A(_01397_),
    .B(_01419_),
    .C(_01421_),
    .Y(_01423_));
 sky130_fd_sc_hd__inv_2 _24552_ (.A(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__and3_1 _24553_ (.A(_01419_),
    .B(_01421_),
    .C(_01396_),
    .X(_01426_));
 sky130_fd_sc_hd__a21oi_2 _24554_ (.A1(_01419_),
    .A2(_01421_),
    .B1(_01396_),
    .Y(_01427_));
 sky130_fd_sc_hd__o211ai_2 _24555_ (.A1(_01422_),
    .A2(_01424_),
    .B1(_01394_),
    .C1(_01395_),
    .Y(_01428_));
 sky130_fd_sc_hd__o2bb2ai_1 _24556_ (.A1_N(_01394_),
    .A2_N(_01395_),
    .B1(_01426_),
    .B2(_01427_),
    .Y(_01429_));
 sky130_fd_sc_hd__o2bb2ai_1 _24557_ (.A1_N(_01394_),
    .A2_N(_01395_),
    .B1(_01422_),
    .B2(_01424_),
    .Y(_01430_));
 sky130_fd_sc_hd__o21ai_2 _24558_ (.A1(_01426_),
    .A2(_01427_),
    .B1(_01395_),
    .Y(_01431_));
 sky130_fd_sc_hd__o211ai_2 _24559_ (.A1(_01426_),
    .A2(_01427_),
    .B1(_01394_),
    .C1(_01395_),
    .Y(_01432_));
 sky130_fd_sc_hd__o2bb2ai_1 _24560_ (.A1_N(_01090_),
    .A2_N(_01163_),
    .B1(_01160_),
    .B2(_01157_),
    .Y(_01433_));
 sky130_fd_sc_hd__a21boi_1 _24561_ (.A1(_01090_),
    .A2(_01163_),
    .B1_N(_01161_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand3_2 _24562_ (.A(_01428_),
    .B(_01429_),
    .C(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__and3_2 _24563_ (.A(_01430_),
    .B(_01432_),
    .C(_01433_),
    .X(_01437_));
 sky130_fd_sc_hd__nand3_2 _24564_ (.A(_01430_),
    .B(_01432_),
    .C(_01433_),
    .Y(_01438_));
 sky130_fd_sc_hd__o211a_1 _24565_ (.A1(_00966_),
    .A2(_00968_),
    .B1(_00971_),
    .C1(_01024_),
    .X(_01439_));
 sky130_fd_sc_hd__o21ai_1 _24566_ (.A1(_00972_),
    .A2(_01023_),
    .B1(_01022_),
    .Y(_01440_));
 sky130_fd_sc_hd__o31a_1 _24567_ (.A1(_00969_),
    .A2(_00970_),
    .A3(_01023_),
    .B1(_01022_),
    .X(_01441_));
 sky130_fd_sc_hd__a21oi_1 _24568_ (.A1(_01435_),
    .A2(_01438_),
    .B1(_01440_),
    .Y(_01442_));
 sky130_fd_sc_hd__a21o_1 _24569_ (.A1(_01435_),
    .A2(_01438_),
    .B1(_01440_),
    .X(_01443_));
 sky130_fd_sc_hd__a31o_1 _24570_ (.A1(_01428_),
    .A2(_01429_),
    .A3(_01434_),
    .B1(_01441_),
    .X(_01444_));
 sky130_fd_sc_hd__and3_2 _24571_ (.A(_01435_),
    .B(_01438_),
    .C(_01440_),
    .X(_01445_));
 sky130_fd_sc_hd__o211ai_1 _24572_ (.A1(_01021_),
    .A2(_01439_),
    .B1(_01438_),
    .C1(_01435_),
    .Y(_01446_));
 sky130_fd_sc_hd__and3_1 _24573_ (.A(_01435_),
    .B(_01438_),
    .C(_01441_),
    .X(_01448_));
 sky130_fd_sc_hd__o2bb2a_1 _24574_ (.A1_N(_01435_),
    .A2_N(_01438_),
    .B1(_01439_),
    .B2(_01021_),
    .X(_01449_));
 sky130_fd_sc_hd__o21ai_2 _24575_ (.A1(_01437_),
    .A2(_01444_),
    .B1(_01443_),
    .Y(_01450_));
 sky130_fd_sc_hd__o2bb2ai_2 _24576_ (.A1_N(_01357_),
    .A2_N(_01360_),
    .B1(_01442_),
    .B2(_01445_),
    .Y(_01451_));
 sky130_fd_sc_hd__and3_1 _24577_ (.A(_01357_),
    .B(_01443_),
    .C(_01446_),
    .X(_01452_));
 sky130_fd_sc_hd__o2111ai_4 _24578_ (.A1(_01437_),
    .A2(_01444_),
    .B1(_01443_),
    .C1(_01357_),
    .D1(_01360_),
    .Y(_01453_));
 sky130_fd_sc_hd__o211ai_2 _24579_ (.A1(_01442_),
    .A2(_01445_),
    .B1(_01357_),
    .C1(_01360_),
    .Y(_01454_));
 sky130_fd_sc_hd__o2bb2ai_1 _24580_ (.A1_N(_01357_),
    .A2_N(_01360_),
    .B1(_01448_),
    .B2(_01449_),
    .Y(_01455_));
 sky130_fd_sc_hd__nand3_2 _24581_ (.A(_01218_),
    .B(_01451_),
    .C(_01453_),
    .Y(_01456_));
 sky130_fd_sc_hd__o2111ai_4 _24582_ (.A1(_01040_),
    .A2(_01178_),
    .B1(_01182_),
    .C1(_01454_),
    .D1(_01455_),
    .Y(_01457_));
 sky130_fd_sc_hd__o211ai_4 _24583_ (.A1(_01032_),
    .A2(_01039_),
    .B1(_01456_),
    .C1(_01457_),
    .Y(_01459_));
 sky130_fd_sc_hd__a21o_2 _24584_ (.A1(_01456_),
    .A2(_01457_),
    .B1(_01217_),
    .X(_01460_));
 sky130_fd_sc_hd__nor2_1 _24585_ (.A(_01192_),
    .B(_01188_),
    .Y(_01461_));
 sky130_fd_sc_hd__a41o_1 _24586_ (.A1(_00890_),
    .A2(_00932_),
    .A3(_01185_),
    .A4(_01186_),
    .B1(_01192_),
    .X(_01462_));
 sky130_fd_sc_hd__o211a_1 _24587_ (.A1(_01188_),
    .A2(_01197_),
    .B1(_01459_),
    .C1(_01460_),
    .X(_01463_));
 sky130_fd_sc_hd__o211ai_4 _24588_ (.A1(_01188_),
    .A2(_01197_),
    .B1(_01459_),
    .C1(_01460_),
    .Y(_01464_));
 sky130_fd_sc_hd__a22oi_4 _24589_ (.A1(_01459_),
    .A2(_01460_),
    .B1(_01462_),
    .B2(_01191_),
    .Y(_01465_));
 sky130_fd_sc_hd__o2bb2ai_1 _24590_ (.A1_N(_01459_),
    .A2_N(_01460_),
    .B1(_01461_),
    .B2(_01190_),
    .Y(_01466_));
 sky130_fd_sc_hd__o21ai_1 _24591_ (.A1(_00966_),
    .A2(_00969_),
    .B1(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__o21ai_2 _24592_ (.A1(_01463_),
    .A2(_01465_),
    .B1(_01214_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand3_1 _24593_ (.A(_01466_),
    .B(_01215_),
    .C(_01464_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand4_2 _24594_ (.A(_01200_),
    .B(_01204_),
    .C(_01468_),
    .D(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__a22oi_2 _24595_ (.A1(_01200_),
    .A2(_01204_),
    .B1(_01468_),
    .B2(_01470_),
    .Y(_01472_));
 sky130_fd_sc_hd__a22o_1 _24596_ (.A1(_01200_),
    .A2(_01204_),
    .B1(_01468_),
    .B2(_01470_),
    .X(_01473_));
 sky130_fd_sc_hd__nand2_1 _24597_ (.A(_01471_),
    .B(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__o2111a_1 _24598_ (.A1(_01203_),
    .A2(_01211_),
    .B1(_01209_),
    .C1(_00920_),
    .D1(_00923_),
    .X(_01475_));
 sky130_fd_sc_hd__nand3_2 _24599_ (.A(_00307_),
    .B(_00926_),
    .C(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__o22ai_2 _24600_ (.A1(_01203_),
    .A2(_01211_),
    .B1(_00923_),
    .B2(_01208_),
    .Y(_01477_));
 sky130_fd_sc_hd__a31oi_4 _24601_ (.A1(_00924_),
    .A2(_01212_),
    .A3(_00927_),
    .B1(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_4 _24602_ (.A(_01476_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__nand4_4 _24603_ (.A(_12394_),
    .B(_01476_),
    .C(_01478_),
    .D(_12398_),
    .Y(_01481_));
 sky130_fd_sc_hd__and4b_4 _24604_ (.A_N(_00302_),
    .B(_00303_),
    .C(_00926_),
    .D(_01475_),
    .X(_01482_));
 sky130_fd_sc_hd__o22a_1 _24605_ (.A1(_01479_),
    .A2(_01482_),
    .B1(_01481_),
    .B2(_12401_),
    .X(_01483_));
 sky130_fd_sc_hd__o22ai_2 _24606_ (.A1(_01479_),
    .A2(_01482_),
    .B1(_01481_),
    .B2(_12401_),
    .Y(_01484_));
 sky130_fd_sc_hd__xor2_1 _24607_ (.A(_01474_),
    .B(_01484_),
    .X(net107));
 sky130_fd_sc_hd__a32o_1 _24608_ (.A1(_01218_),
    .A2(_01451_),
    .A3(_01453_),
    .B1(_01457_),
    .B2(_01217_),
    .X(_01485_));
 sky130_fd_sc_hd__a32oi_2 _24609_ (.A1(_01218_),
    .A2(_01451_),
    .A3(_01453_),
    .B1(_01457_),
    .B2(_01217_),
    .Y(_01486_));
 sky130_fd_sc_hd__a31o_1 _24610_ (.A1(_01430_),
    .A2(_01432_),
    .A3(_01433_),
    .B1(_01445_),
    .X(_01487_));
 sky130_fd_sc_hd__and3_2 _24611_ (.A(_04102_),
    .B(net24),
    .C(net42),
    .X(_01488_));
 sky130_fd_sc_hd__o311a_1 _24612_ (.A1(net176),
    .A2(_07074_),
    .A3(net268),
    .B1(_04895_),
    .C1(net164),
    .X(_01489_));
 sky130_fd_sc_hd__a31oi_4 _24613_ (.A1(net164),
    .A2(_08208_),
    .A3(_04895_),
    .B1(_01488_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _24614_ (.A(_04267_),
    .B(_08664_),
    .Y(_01492_));
 sky130_fd_sc_hd__a31oi_4 _24615_ (.A1(net319),
    .A2(net162),
    .A3(_04267_),
    .B1(_01287_),
    .Y(_01493_));
 sky130_fd_sc_hd__a21oi_1 _24616_ (.A1(_08665_),
    .A2(_08668_),
    .B1(_04481_),
    .Y(_01494_));
 sky130_fd_sc_hd__o21ai_4 _24617_ (.A1(_08664_),
    .A2(_08666_),
    .B1(_04480_),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_1 _24618_ (.A(net319),
    .B(_04483_),
    .Y(_01496_));
 sky130_fd_sc_hd__or3b_4 _24619_ (.A(net42),
    .B(net319),
    .C_N(net41),
    .X(_01497_));
 sky130_fd_sc_hd__a21oi_1 _24620_ (.A1(_08670_),
    .A2(_04480_),
    .B1(_01496_),
    .Y(_01498_));
 sky130_fd_sc_hd__a22oi_4 _24621_ (.A1(_01288_),
    .A2(_01492_),
    .B1(_01495_),
    .B2(_01497_),
    .Y(_01499_));
 sky130_fd_sc_hd__o21bai_1 _24622_ (.A1(_01494_),
    .A2(_01496_),
    .B1_N(_01493_),
    .Y(_01500_));
 sky130_fd_sc_hd__o211a_1 _24623_ (.A1(net319),
    .A2(_04483_),
    .B1(_01493_),
    .C1(_01495_),
    .X(_01502_));
 sky130_fd_sc_hd__o2111ai_4 _24624_ (.A1(_04268_),
    .A2(_08665_),
    .B1(_01288_),
    .C1(_01495_),
    .D1(_01497_),
    .Y(_01503_));
 sky130_fd_sc_hd__o21ai_2 _24625_ (.A1(_01499_),
    .A2(_01502_),
    .B1(_01491_),
    .Y(_01504_));
 sky130_fd_sc_hd__a31oi_2 _24626_ (.A1(_01495_),
    .A2(_01497_),
    .A3(_01493_),
    .B1(_01491_),
    .Y(_01505_));
 sky130_fd_sc_hd__a31o_1 _24627_ (.A1(_01495_),
    .A2(_01497_),
    .A3(_01493_),
    .B1(_01491_),
    .X(_01506_));
 sky130_fd_sc_hd__o22ai_4 _24628_ (.A1(_01488_),
    .A2(_01489_),
    .B1(_01499_),
    .B2(_01502_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand3_2 _24629_ (.A(_01500_),
    .B(_01503_),
    .C(_01491_),
    .Y(_01508_));
 sky130_fd_sc_hd__a31o_1 _24630_ (.A1(_01286_),
    .A2(_01288_),
    .A3(_01284_),
    .B1(_01278_),
    .X(_01509_));
 sky130_fd_sc_hd__o21ai_1 _24631_ (.A1(_01284_),
    .A2(_01289_),
    .B1(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__a21oi_2 _24632_ (.A1(_01279_),
    .A2(_01294_),
    .B1(_01290_),
    .Y(_01511_));
 sky130_fd_sc_hd__a21oi_2 _24633_ (.A1(_01507_),
    .A2(_01508_),
    .B1(_01511_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand3_4 _24634_ (.A(_01504_),
    .B(_01506_),
    .C(_01510_),
    .Y(_01514_));
 sky130_fd_sc_hd__nand3_4 _24635_ (.A(_01507_),
    .B(_01508_),
    .C(_01511_),
    .Y(_01515_));
 sky130_fd_sc_hd__o22a_1 _24636_ (.A1(_04212_),
    .A2(_05465_),
    .B1(_07079_),
    .B2(_05463_),
    .X(_01516_));
 sky130_fd_sc_hd__a32o_1 _24637_ (.A1(_07072_),
    .A2(net170),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net20),
    .X(_01517_));
 sky130_fd_sc_hd__nor2_1 _24638_ (.A(_04223_),
    .B(_05229_),
    .Y(_01518_));
 sky130_fd_sc_hd__a31oi_2 _24639_ (.A1(_07499_),
    .A2(_07503_),
    .A3(_05225_),
    .B1(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__or3_1 _24640_ (.A(net45),
    .B(_04245_),
    .C(_04102_),
    .X(_01520_));
 sky130_fd_sc_hd__o211ai_2 _24641_ (.A1(net170),
    .A2(_07765_),
    .B1(net242),
    .C1(_07771_),
    .Y(_01521_));
 sky130_fd_sc_hd__a21oi_1 _24642_ (.A1(_01520_),
    .A2(_01521_),
    .B1(_01519_),
    .Y(_01522_));
 sky130_fd_sc_hd__a21o_1 _24643_ (.A1(_01520_),
    .A2(_01521_),
    .B1(_01519_),
    .X(_01524_));
 sky130_fd_sc_hd__nand3_2 _24644_ (.A(_01519_),
    .B(_01520_),
    .C(_01521_),
    .Y(_01525_));
 sky130_fd_sc_hd__a21oi_1 _24645_ (.A1(_01524_),
    .A2(_01525_),
    .B1(_01517_),
    .Y(_01526_));
 sky130_fd_sc_hd__and3_1 _24646_ (.A(_01517_),
    .B(_01524_),
    .C(_01525_),
    .X(_01527_));
 sky130_fd_sc_hd__nand3_1 _24647_ (.A(_01524_),
    .B(_01525_),
    .C(_01516_),
    .Y(_01528_));
 sky130_fd_sc_hd__a21o_1 _24648_ (.A1(_01524_),
    .A2(_01525_),
    .B1(_01516_),
    .X(_01529_));
 sky130_fd_sc_hd__nand2_2 _24649_ (.A(_01528_),
    .B(_01529_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand3_4 _24650_ (.A(_01514_),
    .B(_01515_),
    .C(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__o2bb2ai_4 _24651_ (.A1_N(_01514_),
    .A2_N(_01515_),
    .B1(_01526_),
    .B2(_01527_),
    .Y(_01532_));
 sky130_fd_sc_hd__o2111a_2 _24652_ (.A1(_00796_),
    .A2(_01324_),
    .B1(_01329_),
    .C1(_01531_),
    .D1(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__o2111ai_4 _24653_ (.A1(_00796_),
    .A2(_01324_),
    .B1(_01329_),
    .C1(_01531_),
    .D1(_01532_),
    .Y(_01535_));
 sky130_fd_sc_hd__a22oi_4 _24654_ (.A1(_01329_),
    .A2(_01332_),
    .B1(_01531_),
    .B2(_01532_),
    .Y(_01536_));
 sky130_fd_sc_hd__a22o_1 _24655_ (.A1(_01329_),
    .A2(_01332_),
    .B1(_01531_),
    .B2(_01532_),
    .X(_01537_));
 sky130_fd_sc_hd__o22ai_4 _24656_ (.A1(_00360_),
    .A2(_11741_),
    .B1(_01536_),
    .B2(_01533_),
    .Y(_01538_));
 sky130_fd_sc_hd__nand3_2 _24657_ (.A(_01537_),
    .B(net130),
    .C(_01535_),
    .Y(_01539_));
 sky130_fd_sc_hd__a211oi_2 _24658_ (.A1(_01538_),
    .A2(_01539_),
    .B1(_01330_),
    .C1(_01338_),
    .Y(_01540_));
 sky130_fd_sc_hd__a211o_1 _24659_ (.A1(_01538_),
    .A2(_01539_),
    .B1(_01330_),
    .C1(_01338_),
    .X(_01541_));
 sky130_fd_sc_hd__o211a_1 _24660_ (.A1(_01330_),
    .A2(_01338_),
    .B1(_01538_),
    .C1(_01539_),
    .X(_01542_));
 sky130_fd_sc_hd__o211ai_2 _24661_ (.A1(_01330_),
    .A2(_01338_),
    .B1(_01538_),
    .C1(_01539_),
    .Y(_01543_));
 sky130_fd_sc_hd__nor2_1 _24662_ (.A(_01540_),
    .B(_01542_),
    .Y(_01544_));
 sky130_fd_sc_hd__nand2_2 _24663_ (.A(_01541_),
    .B(_01543_),
    .Y(_01546_));
 sky130_fd_sc_hd__o22ai_2 _24664_ (.A1(_01252_),
    .A2(_01244_),
    .B1(net132),
    .B2(_01250_),
    .Y(_01547_));
 sky130_fd_sc_hd__a21oi_1 _24665_ (.A1(net133),
    .A2(_01239_),
    .B1(_01240_),
    .Y(_01548_));
 sky130_fd_sc_hd__a21o_1 _24666_ (.A1(net133),
    .A2(_01239_),
    .B1(_01240_),
    .X(_01549_));
 sky130_fd_sc_hd__or3_2 _24667_ (.A(net57),
    .B(_04266_),
    .C(_04080_),
    .X(_01550_));
 sky130_fd_sc_hd__nand3_4 _24668_ (.A(net220),
    .B(net186),
    .C(_08657_),
    .Y(_01551_));
 sky130_fd_sc_hd__a21oi_4 _24669_ (.A1(_01550_),
    .A2(_01551_),
    .B1(_08878_),
    .Y(_01552_));
 sky130_fd_sc_hd__a21o_1 _24670_ (.A1(_01550_),
    .A2(_01551_),
    .B1(_08878_),
    .X(_01553_));
 sky130_fd_sc_hd__o311a_2 _24671_ (.A1(_04080_),
    .A2(net57),
    .A3(_04266_),
    .B1(_01551_),
    .C1(_08878_),
    .X(_01554_));
 sky130_fd_sc_hd__nand3_2 _24672_ (.A(_08878_),
    .B(_01550_),
    .C(_01551_),
    .Y(_01555_));
 sky130_fd_sc_hd__o21ai_1 _24673_ (.A1(_01552_),
    .A2(_01554_),
    .B1(net146),
    .Y(_01557_));
 sky130_fd_sc_hd__o22ai_4 _24674_ (.A1(_08881_),
    .A2(_09297_),
    .B1(_01552_),
    .B2(_01554_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand3_2 _24675_ (.A(_01553_),
    .B(_01555_),
    .C(net146),
    .Y(_01559_));
 sky130_fd_sc_hd__a21oi_2 _24676_ (.A1(net156),
    .A2(_01225_),
    .B1(_09300_),
    .Y(_01560_));
 sky130_fd_sc_hd__a22oi_2 _24677_ (.A1(_01230_),
    .A2(_01232_),
    .B1(_01558_),
    .B2(_01559_),
    .Y(_01561_));
 sky130_fd_sc_hd__o221ai_4 _24678_ (.A1(_01229_),
    .A2(_01231_),
    .B1(_01554_),
    .B2(net146),
    .C1(_01557_),
    .Y(_01562_));
 sky130_fd_sc_hd__o211a_2 _24679_ (.A1(_01226_),
    .A2(_01560_),
    .B1(_01559_),
    .C1(_01558_),
    .X(_01563_));
 sky130_fd_sc_hd__o211ai_4 _24680_ (.A1(_01226_),
    .A2(_01560_),
    .B1(_01559_),
    .C1(_01558_),
    .Y(_01564_));
 sky130_fd_sc_hd__o22ai_4 _24681_ (.A1(_10540_),
    .A2(net135),
    .B1(_01561_),
    .B2(_01563_),
    .Y(_01565_));
 sky130_fd_sc_hd__nand4_1 _24682_ (.A(net138),
    .B(net134),
    .C(_01562_),
    .D(_01564_),
    .Y(_01566_));
 sky130_fd_sc_hd__a21o_1 _24683_ (.A1(_01562_),
    .A2(_01564_),
    .B1(_10546_),
    .X(_01568_));
 sky130_fd_sc_hd__o211ai_1 _24684_ (.A1(_10540_),
    .A2(net135),
    .B1(_01562_),
    .C1(_01564_),
    .Y(_01569_));
 sky130_fd_sc_hd__a21oi_1 _24685_ (.A1(_01565_),
    .A2(_01566_),
    .B1(_01549_),
    .Y(_01570_));
 sky130_fd_sc_hd__nand3_2 _24686_ (.A(_01568_),
    .B(_01569_),
    .C(_01548_),
    .Y(_01571_));
 sky130_fd_sc_hd__a32oi_4 _24687_ (.A1(net133),
    .A2(_01562_),
    .A3(_01564_),
    .B1(_01241_),
    .B2(_01245_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand3_2 _24688_ (.A(_01549_),
    .B(_01565_),
    .C(_01566_),
    .Y(_01573_));
 sky130_fd_sc_hd__a21oi_1 _24689_ (.A1(_01571_),
    .A2(_01573_),
    .B1(_12099_),
    .Y(_01574_));
 sky130_fd_sc_hd__a21o_1 _24690_ (.A1(_01571_),
    .A2(_01573_),
    .B1(_12099_),
    .X(_01575_));
 sky130_fd_sc_hd__o311a_1 _24691_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_01571_),
    .C1(_01573_),
    .X(_01576_));
 sky130_fd_sc_hd__o211ai_4 _24692_ (.A1(_11742_),
    .A2(_11042_),
    .B1(_01573_),
    .C1(_01571_),
    .Y(_01577_));
 sky130_fd_sc_hd__a21oi_2 _24693_ (.A1(_01575_),
    .A2(_01577_),
    .B1(_01547_),
    .Y(_01579_));
 sky130_fd_sc_hd__o21bai_4 _24694_ (.A1(_01574_),
    .A2(_01576_),
    .B1_N(_01547_),
    .Y(_01580_));
 sky130_fd_sc_hd__o211a_1 _24695_ (.A1(_01253_),
    .A2(_01257_),
    .B1(_01575_),
    .C1(_01577_),
    .X(_01581_));
 sky130_fd_sc_hd__o211ai_4 _24696_ (.A1(_01253_),
    .A2(_01257_),
    .B1(_01575_),
    .C1(_01577_),
    .Y(_01582_));
 sky130_fd_sc_hd__o22ai_4 _24697_ (.A1(net130),
    .A2(_00366_),
    .B1(_01579_),
    .B2(_01581_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _24698_ (.A(_01580_),
    .B(_00736_),
    .Y(_01584_));
 sky130_fd_sc_hd__and3_1 _24699_ (.A(_01580_),
    .B(_01582_),
    .C(_00736_),
    .X(_01585_));
 sky130_fd_sc_hd__o2111ai_4 _24700_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_01580_),
    .D1(_01582_),
    .Y(_01586_));
 sky130_fd_sc_hd__o21ai_4 _24701_ (.A1(_00737_),
    .A2(_01262_),
    .B1(_01261_),
    .Y(_01587_));
 sky130_fd_sc_hd__a21oi_4 _24702_ (.A1(_01583_),
    .A2(_01586_),
    .B1(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__a21o_1 _24703_ (.A1(_01583_),
    .A2(_01586_),
    .B1(_01587_),
    .X(_01590_));
 sky130_fd_sc_hd__nand2_2 _24704_ (.A(_01587_),
    .B(_01583_),
    .Y(_01591_));
 sky130_fd_sc_hd__o211a_1 _24705_ (.A1(_01581_),
    .A2(_01584_),
    .B1(_01583_),
    .C1(_01587_),
    .X(_01592_));
 sky130_fd_sc_hd__a31o_1 _24706_ (.A1(_00736_),
    .A2(_01580_),
    .A3(_01582_),
    .B1(_01591_),
    .X(_01593_));
 sky130_fd_sc_hd__o22ai_4 _24707_ (.A1(_01540_),
    .A2(_01542_),
    .B1(_01588_),
    .B2(_01592_),
    .Y(_01594_));
 sky130_fd_sc_hd__o211ai_4 _24708_ (.A1(_01585_),
    .A2(_01591_),
    .B1(_01590_),
    .C1(_01544_),
    .Y(_01595_));
 sky130_fd_sc_hd__o22a_1 _24709_ (.A1(_01347_),
    .A2(_01349_),
    .B1(_01219_),
    .B2(_01268_),
    .X(_01596_));
 sky130_fd_sc_hd__o21a_1 _24710_ (.A1(_01344_),
    .A2(_01345_),
    .B1(_01273_),
    .X(_01597_));
 sky130_fd_sc_hd__o21ai_1 _24711_ (.A1(_01344_),
    .A2(_01345_),
    .B1(_01273_),
    .Y(_01598_));
 sky130_fd_sc_hd__o21ai_1 _24712_ (.A1(_01219_),
    .A2(_01268_),
    .B1(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__a21oi_2 _24713_ (.A1(_01594_),
    .A2(_01595_),
    .B1(_01599_),
    .Y(_01601_));
 sky130_fd_sc_hd__o2bb2ai_1 _24714_ (.A1_N(_01594_),
    .A2_N(_01595_),
    .B1(_01596_),
    .B2(_01272_),
    .Y(_01602_));
 sky130_fd_sc_hd__o211a_2 _24715_ (.A1(_01269_),
    .A2(_01597_),
    .B1(_01595_),
    .C1(_01594_),
    .X(_01603_));
 sky130_fd_sc_hd__o211ai_1 _24716_ (.A1(_01269_),
    .A2(_01597_),
    .B1(_01595_),
    .C1(_01594_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _24717_ (.A(_01386_),
    .B(_01393_),
    .Y(_01605_));
 sky130_fd_sc_hd__a21oi_1 _24718_ (.A1(_01363_),
    .A2(_01369_),
    .B1(_01371_),
    .Y(_01606_));
 sky130_fd_sc_hd__and3_1 _24719_ (.A(net202),
    .B(net173),
    .C(net273),
    .X(_01607_));
 sky130_fd_sc_hd__and3_1 _24720_ (.A(_04190_),
    .B(net49),
    .C(net17),
    .X(_01608_));
 sky130_fd_sc_hd__a31o_1 _24721_ (.A1(net202),
    .A2(net173),
    .A3(net273),
    .B1(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__or3b_1 _24722_ (.A(net48),
    .B(_04201_),
    .C_N(net47),
    .X(_01610_));
 sky130_fd_sc_hd__o211ai_2 _24723_ (.A1(net176),
    .A2(_06759_),
    .B1(_05762_),
    .C1(net191),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_1 _24724_ (.A(_04179_),
    .B(_06030_),
    .Y(_01613_));
 sky130_fd_sc_hd__o311a_1 _24725_ (.A1(net244),
    .A2(net241),
    .A3(_06451_),
    .B1(net274),
    .C1(net197),
    .X(_01614_));
 sky130_fd_sc_hd__a31oi_1 _24726_ (.A1(net197),
    .A2(_06452_),
    .A3(net274),
    .B1(_01613_),
    .Y(_01615_));
 sky130_fd_sc_hd__o2bb2a_2 _24727_ (.A1_N(_01610_),
    .A2_N(_01612_),
    .B1(_01613_),
    .B2(_01614_),
    .X(_01616_));
 sky130_fd_sc_hd__o2bb2ai_1 _24728_ (.A1_N(_01610_),
    .A2_N(_01612_),
    .B1(_01613_),
    .B2(_01614_),
    .Y(_01617_));
 sky130_fd_sc_hd__o211ai_2 _24729_ (.A1(_04201_),
    .A2(_05766_),
    .B1(_01612_),
    .C1(_01615_),
    .Y(_01618_));
 sky130_fd_sc_hd__a21oi_1 _24730_ (.A1(_01617_),
    .A2(_01618_),
    .B1(_01609_),
    .Y(_01619_));
 sky130_fd_sc_hd__a21o_1 _24731_ (.A1(_01617_),
    .A2(_01618_),
    .B1(_01609_),
    .X(_01620_));
 sky130_fd_sc_hd__o211a_2 _24732_ (.A1(_01607_),
    .A2(_01608_),
    .B1(_01617_),
    .C1(_01618_),
    .X(_01621_));
 sky130_fd_sc_hd__o211ai_1 _24733_ (.A1(_01607_),
    .A2(_01608_),
    .B1(_01617_),
    .C1(_01618_),
    .Y(_01623_));
 sky130_fd_sc_hd__o2bb2ai_1 _24734_ (.A1_N(_01307_),
    .A2_N(_01309_),
    .B1(_01302_),
    .B2(_01303_),
    .Y(_01624_));
 sky130_fd_sc_hd__o21ai_1 _24735_ (.A1(_01307_),
    .A2(_01309_),
    .B1(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__o221a_1 _24736_ (.A1(_01307_),
    .A2(_01309_),
    .B1(_01619_),
    .B2(_01621_),
    .C1(_01624_),
    .X(_01626_));
 sky130_fd_sc_hd__o21bai_2 _24737_ (.A1(_01619_),
    .A2(_01621_),
    .B1_N(_01625_),
    .Y(_01627_));
 sky130_fd_sc_hd__nand3_2 _24738_ (.A(_01620_),
    .B(_01623_),
    .C(_01625_),
    .Y(_01628_));
 sky130_fd_sc_hd__a21boi_1 _24739_ (.A1(_01627_),
    .A2(_01628_),
    .B1_N(_01606_),
    .Y(_01629_));
 sky130_fd_sc_hd__a221o_1 _24740_ (.A1(_01363_),
    .A2(_01369_),
    .B1(_01627_),
    .B2(_01628_),
    .C1(_01371_),
    .X(_01630_));
 sky130_fd_sc_hd__o211a_1 _24741_ (.A1(_01371_),
    .A2(_01374_),
    .B1(_01627_),
    .C1(_01628_),
    .X(_01631_));
 sky130_fd_sc_hd__o211ai_1 _24742_ (.A1(_01371_),
    .A2(_01374_),
    .B1(_01627_),
    .C1(_01628_),
    .Y(_01632_));
 sky130_fd_sc_hd__a21o_1 _24743_ (.A1(_01301_),
    .A2(_01316_),
    .B1(_01299_),
    .X(_01634_));
 sky130_fd_sc_hd__o211ai_4 _24744_ (.A1(_01629_),
    .A2(_01631_),
    .B1(_01300_),
    .C1(_01318_),
    .Y(_01635_));
 sky130_fd_sc_hd__nand3_2 _24745_ (.A(_01630_),
    .B(_01632_),
    .C(_01634_),
    .Y(_01636_));
 sky130_fd_sc_hd__and3_1 _24746_ (.A(_00992_),
    .B(_00994_),
    .C(_01378_),
    .X(_01637_));
 sky130_fd_sc_hd__o21ai_2 _24747_ (.A1(_01361_),
    .A2(_01376_),
    .B1(_01378_),
    .Y(_01638_));
 sky130_fd_sc_hd__nand3_2 _24748_ (.A(_01635_),
    .B(_01636_),
    .C(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__o2bb2ai_4 _24749_ (.A1_N(_01635_),
    .A2_N(_01636_),
    .B1(_01637_),
    .B2(_01376_),
    .Y(_01640_));
 sky130_fd_sc_hd__o211a_2 _24750_ (.A1(_01387_),
    .A2(_01391_),
    .B1(_01639_),
    .C1(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__o211ai_2 _24751_ (.A1(_01387_),
    .A2(_01391_),
    .B1(_01639_),
    .C1(_01640_),
    .Y(_01642_));
 sky130_fd_sc_hd__o2bb2a_2 _24752_ (.A1_N(_04792_),
    .A2_N(net238),
    .B1(_08007_),
    .B2(_04091_),
    .X(_01643_));
 sky130_fd_sc_hd__and3b_1 _24753_ (.A_N(net54),
    .B(net53),
    .C(net13),
    .X(_01645_));
 sky130_fd_sc_hd__o311a_1 _24754_ (.A1(net11),
    .A2(_04557_),
    .A3(_05073_),
    .B1(_07642_),
    .C1(net209),
    .X(_01646_));
 sky130_fd_sc_hd__a21oi_2 _24755_ (.A1(net13),
    .A2(_07643_),
    .B1(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__a21oi_2 _24756_ (.A1(_01400_),
    .A2(_01409_),
    .B1(_01406_),
    .Y(_01648_));
 sky130_fd_sc_hd__a21o_1 _24757_ (.A1(_01400_),
    .A2(_01409_),
    .B1(_01406_),
    .X(_01649_));
 sky130_fd_sc_hd__a32o_1 _24758_ (.A1(_05290_),
    .A2(_05292_),
    .A3(net239),
    .B1(_07308_),
    .B2(net14),
    .X(_01650_));
 sky130_fd_sc_hd__nor2_1 _24759_ (.A(_04157_),
    .B(_06866_),
    .Y(_01651_));
 sky130_fd_sc_hd__a211oi_2 _24760_ (.A1(_05553_),
    .A2(net16),
    .B1(_06864_),
    .C1(net204),
    .Y(_01652_));
 sky130_fd_sc_hd__o221ai_4 _24761_ (.A1(net233),
    .A2(_05927_),
    .B1(_04157_),
    .B2(net207),
    .C1(net240),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _24762_ (.A(_04146_),
    .B(_07226_),
    .Y(_01654_));
 sky130_fd_sc_hd__or3b_1 _24763_ (.A(_04146_),
    .B(net52),
    .C_N(net51),
    .X(_01656_));
 sky130_fd_sc_hd__a211oi_4 _24764_ (.A1(_04788_),
    .A2(_05550_),
    .B1(_07224_),
    .C1(_05548_),
    .Y(_01657_));
 sky130_fd_sc_hd__o211ai_2 _24765_ (.A1(_04789_),
    .A2(_05551_),
    .B1(net269),
    .C1(net178),
    .Y(_01658_));
 sky130_fd_sc_hd__o22a_1 _24766_ (.A1(_01651_),
    .A2(_01652_),
    .B1(_01654_),
    .B2(_01657_),
    .X(_01659_));
 sky130_fd_sc_hd__o22ai_4 _24767_ (.A1(_01651_),
    .A2(_01652_),
    .B1(_01654_),
    .B2(_01657_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand4b_4 _24768_ (.A_N(_01651_),
    .B(_01653_),
    .C(_01656_),
    .D(_01658_),
    .Y(_01661_));
 sky130_fd_sc_hd__a21o_1 _24769_ (.A1(_01660_),
    .A2(_01661_),
    .B1(_01650_),
    .X(_01662_));
 sky130_fd_sc_hd__nand3_1 _24770_ (.A(_01650_),
    .B(_01660_),
    .C(_01661_),
    .Y(_01663_));
 sky130_fd_sc_hd__a21bo_1 _24771_ (.A1(_01660_),
    .A2(_01661_),
    .B1_N(_01650_),
    .X(_01664_));
 sky130_fd_sc_hd__nand3b_2 _24772_ (.A_N(_01650_),
    .B(_01660_),
    .C(_01661_),
    .Y(_01665_));
 sky130_fd_sc_hd__nand3_1 _24773_ (.A(_01649_),
    .B(_01662_),
    .C(_01663_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand3_1 _24774_ (.A(_01664_),
    .B(_01665_),
    .C(_01648_),
    .Y(_01668_));
 sky130_fd_sc_hd__nand3_1 _24775_ (.A(_01662_),
    .B(_01663_),
    .C(_01648_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand3_1 _24776_ (.A(_01649_),
    .B(_01664_),
    .C(_01665_),
    .Y(_01670_));
 sky130_fd_sc_hd__o211ai_2 _24777_ (.A1(_01645_),
    .A2(_01646_),
    .B1(_01669_),
    .C1(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__nand3_1 _24778_ (.A(_01667_),
    .B(_01668_),
    .C(_01647_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand2_1 _24779_ (.A(_01399_),
    .B(_01415_),
    .Y(_01673_));
 sky130_fd_sc_hd__a22oi_2 _24780_ (.A1(_01671_),
    .A2(_01672_),
    .B1(_01673_),
    .B2(_01416_),
    .Y(_01674_));
 sky130_fd_sc_hd__and4_1 _24781_ (.A(_01416_),
    .B(_01671_),
    .C(_01672_),
    .D(_01673_),
    .X(_01675_));
 sky130_fd_sc_hd__nor2_2 _24782_ (.A(_01674_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__xnor2_4 _24783_ (.A(_01643_),
    .B(_01676_),
    .Y(_01678_));
 sky130_fd_sc_hd__xor2_1 _24784_ (.A(_01643_),
    .B(_01676_),
    .X(_01679_));
 sky130_fd_sc_hd__a21oi_2 _24785_ (.A1(_01639_),
    .A2(_01640_),
    .B1(_01605_),
    .Y(_01680_));
 sky130_fd_sc_hd__a21o_1 _24786_ (.A1(_01639_),
    .A2(_01640_),
    .B1(_01605_),
    .X(_01681_));
 sky130_fd_sc_hd__nand3_1 _24787_ (.A(_01678_),
    .B(_01681_),
    .C(_01642_),
    .Y(_01682_));
 sky130_fd_sc_hd__o21ai_1 _24788_ (.A1(_01641_),
    .A2(_01680_),
    .B1(_01679_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand3_2 _24789_ (.A(_01642_),
    .B(_01679_),
    .C(_01681_),
    .Y(_01684_));
 sky130_fd_sc_hd__o21ai_2 _24790_ (.A1(_01641_),
    .A2(_01680_),
    .B1(_01678_),
    .Y(_01685_));
 sky130_fd_sc_hd__a21oi_2 _24791_ (.A1(_01274_),
    .A2(_01343_),
    .B1(_01342_),
    .Y(_01686_));
 sky130_fd_sc_hd__nand3_2 _24792_ (.A(_01684_),
    .B(_01685_),
    .C(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__o211ai_4 _24793_ (.A1(_01342_),
    .A2(_01346_),
    .B1(_01682_),
    .C1(_01683_),
    .Y(_01689_));
 sky130_fd_sc_hd__o41a_1 _24794_ (.A1(_01011_),
    .A2(_01013_),
    .A3(_01389_),
    .A4(_01391_),
    .B1(_01431_),
    .X(_01690_));
 sky130_fd_sc_hd__a22o_1 _24795_ (.A1(_01394_),
    .A2(_01431_),
    .B1(_01687_),
    .B2(_01689_),
    .X(_01691_));
 sky130_fd_sc_hd__nand4_2 _24796_ (.A(_01394_),
    .B(_01431_),
    .C(_01687_),
    .D(_01689_),
    .Y(_01692_));
 sky130_fd_sc_hd__a21bo_1 _24797_ (.A1(_01687_),
    .A2(_01689_),
    .B1_N(_01690_),
    .X(_01693_));
 sky130_fd_sc_hd__nand3b_1 _24798_ (.A_N(_01690_),
    .B(_01689_),
    .C(_01687_),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _24799_ (.A(_01691_),
    .B(_01692_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand4_2 _24800_ (.A(_01602_),
    .B(_01604_),
    .C(_01691_),
    .D(_01692_),
    .Y(_01696_));
 sky130_fd_sc_hd__o21ai_2 _24801_ (.A1(_01601_),
    .A2(_01603_),
    .B1(_01695_),
    .Y(_01697_));
 sky130_fd_sc_hd__o211ai_1 _24802_ (.A1(_01601_),
    .A2(_01603_),
    .B1(_01691_),
    .C1(_01692_),
    .Y(_01698_));
 sky130_fd_sc_hd__a21oi_1 _24803_ (.A1(_01691_),
    .A2(_01692_),
    .B1(_01601_),
    .Y(_01700_));
 sky130_fd_sc_hd__a211o_1 _24804_ (.A1(_01691_),
    .A2(_01692_),
    .B1(_01601_),
    .C1(_01603_),
    .X(_01701_));
 sky130_fd_sc_hd__a2bb2oi_1 _24805_ (.A1_N(_01358_),
    .A2_N(_01452_),
    .B1(_01696_),
    .B2(_01697_),
    .Y(_01702_));
 sky130_fd_sc_hd__o211ai_2 _24806_ (.A1(_01358_),
    .A2(_01452_),
    .B1(_01698_),
    .C1(_01701_),
    .Y(_01703_));
 sky130_fd_sc_hd__o2111a_1 _24807_ (.A1(_01450_),
    .A2(_01356_),
    .B1(_01360_),
    .C1(_01696_),
    .D1(_01697_),
    .X(_01704_));
 sky130_fd_sc_hd__o2111ai_4 _24808_ (.A1(_01450_),
    .A2(_01356_),
    .B1(_01360_),
    .C1(_01696_),
    .D1(_01697_),
    .Y(_01705_));
 sky130_fd_sc_hd__o21bai_1 _24809_ (.A1(_01702_),
    .A2(_01704_),
    .B1_N(_01487_),
    .Y(_01706_));
 sky130_fd_sc_hd__o211ai_2 _24810_ (.A1(_01437_),
    .A2(_01445_),
    .B1(_01703_),
    .C1(_01705_),
    .Y(_01707_));
 sky130_fd_sc_hd__o22ai_1 _24811_ (.A1(_01437_),
    .A2(_01445_),
    .B1(_01702_),
    .B2(_01704_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand4_1 _24812_ (.A(_01438_),
    .B(_01446_),
    .C(_01703_),
    .D(_01705_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand3_2 _24813_ (.A(_01706_),
    .B(_01707_),
    .C(_01485_),
    .Y(_01711_));
 sky130_fd_sc_hd__nand3_2 _24814_ (.A(_01486_),
    .B(_01708_),
    .C(_01709_),
    .Y(_01712_));
 sky130_fd_sc_hd__and2_1 _24815_ (.A(_01397_),
    .B(_01419_),
    .X(_01713_));
 sky130_fd_sc_hd__a31o_1 _24816_ (.A1(_01398_),
    .A2(_01417_),
    .A3(_01418_),
    .B1(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__o2bb2ai_2 _24817_ (.A1_N(_01711_),
    .A2_N(_01712_),
    .B1(_01713_),
    .B2(_01420_),
    .Y(_01715_));
 sky130_fd_sc_hd__nand4_4 _24818_ (.A(_01421_),
    .B(_01423_),
    .C(_01711_),
    .D(_01712_),
    .Y(_01716_));
 sky130_fd_sc_hd__a22oi_1 _24819_ (.A1(_01464_),
    .A2(_01467_),
    .B1(_01715_),
    .B2(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__a22o_1 _24820_ (.A1(_01464_),
    .A2(_01467_),
    .B1(_01715_),
    .B2(_01716_),
    .X(_01718_));
 sky130_fd_sc_hd__o2111ai_4 _24821_ (.A1(_01215_),
    .A2(_01465_),
    .B1(_01715_),
    .C1(_01716_),
    .D1(_01464_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _24822_ (.A(_01718_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__o21ai_1 _24823_ (.A1(_01472_),
    .A2(_01483_),
    .B1(_01471_),
    .Y(_01722_));
 sky130_fd_sc_hd__xor2_1 _24824_ (.A(_01720_),
    .B(_01722_),
    .X(net108));
 sky130_fd_sc_hd__nand4_2 _24825_ (.A(_01471_),
    .B(_01473_),
    .C(_01718_),
    .D(_01719_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21oi_2 _24826_ (.A1(_01719_),
    .A2(_01472_),
    .B1(_01717_),
    .Y(_01724_));
 sky130_fd_sc_hd__o21a_1 _24827_ (.A1(_01484_),
    .A2(_01723_),
    .B1(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__a32o_1 _24828_ (.A1(_01485_),
    .A2(_01706_),
    .A3(_01707_),
    .B1(_01712_),
    .B2(_01714_),
    .X(_01726_));
 sky130_fd_sc_hd__a21o_1 _24829_ (.A1(_01705_),
    .A2(_01487_),
    .B1(_01702_),
    .X(_01727_));
 sky130_fd_sc_hd__a21oi_1 _24830_ (.A1(_01705_),
    .A2(_01487_),
    .B1(_01702_),
    .Y(_01728_));
 sky130_fd_sc_hd__o2bb2ai_4 _24831_ (.A1_N(_01572_),
    .A2_N(_01565_),
    .B1(net132),
    .B2(_01570_),
    .Y(_01729_));
 sky130_fd_sc_hd__o21a_1 _24832_ (.A1(net140),
    .A2(net136),
    .B1(_01562_),
    .X(_01730_));
 sky130_fd_sc_hd__nand2_1 _24833_ (.A(net133),
    .B(_01564_),
    .Y(_01732_));
 sky130_fd_sc_hd__a21o_1 _24834_ (.A1(net144),
    .A2(_01555_),
    .B1(_01552_),
    .X(_01733_));
 sky130_fd_sc_hd__a21oi_2 _24835_ (.A1(net144),
    .A2(_01555_),
    .B1(_01552_),
    .Y(_01734_));
 sky130_fd_sc_hd__nor2_1 _24836_ (.A(_04091_),
    .B(_08660_),
    .Y(_01735_));
 sky130_fd_sc_hd__or3_2 _24837_ (.A(net57),
    .B(_04266_),
    .C(_04091_),
    .X(_01736_));
 sky130_fd_sc_hd__o211ai_4 _24838_ (.A1(net233),
    .A2(_04787_),
    .B1(_08657_),
    .C1(net213),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_1 _24839_ (.A(net149),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__o311a_2 _24840_ (.A1(_04091_),
    .A2(net57),
    .A3(_04266_),
    .B1(_01737_),
    .C1(net149),
    .X(_01739_));
 sky130_fd_sc_hd__a21oi_4 _24841_ (.A1(_01736_),
    .A2(_01737_),
    .B1(net149),
    .Y(_01740_));
 sky130_fd_sc_hd__a21o_1 _24842_ (.A1(_01736_),
    .A2(_01737_),
    .B1(net149),
    .X(_01741_));
 sky130_fd_sc_hd__o22a_1 _24843_ (.A1(net237),
    .A2(_09297_),
    .B1(_01735_),
    .B2(_01738_),
    .X(_01743_));
 sky130_fd_sc_hd__a31o_1 _24844_ (.A1(net149),
    .A2(_01736_),
    .A3(_01737_),
    .B1(net145),
    .X(_01744_));
 sky130_fd_sc_hd__o21ai_2 _24845_ (.A1(_01739_),
    .A2(_01740_),
    .B1(net145),
    .Y(_01745_));
 sky130_fd_sc_hd__o22ai_4 _24846_ (.A1(net237),
    .A2(_09297_),
    .B1(_01739_),
    .B2(_01740_),
    .Y(_01746_));
 sky130_fd_sc_hd__o211ai_4 _24847_ (.A1(_01735_),
    .A2(_01738_),
    .B1(net145),
    .C1(_01741_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand3_4 _24848_ (.A(_01745_),
    .B(_01733_),
    .C(_01744_),
    .Y(_01748_));
 sky130_fd_sc_hd__and3_2 _24849_ (.A(_01734_),
    .B(_01746_),
    .C(_01747_),
    .X(_01749_));
 sky130_fd_sc_hd__nand3_2 _24850_ (.A(_01734_),
    .B(_01746_),
    .C(_01747_),
    .Y(_01750_));
 sky130_fd_sc_hd__a21oi_2 _24851_ (.A1(_01748_),
    .A2(_01750_),
    .B1(net133),
    .Y(_01751_));
 sky130_fd_sc_hd__a31o_1 _24852_ (.A1(_01745_),
    .A2(_01733_),
    .A3(_01744_),
    .B1(_10546_),
    .X(_01752_));
 sky130_fd_sc_hd__o211ai_2 _24853_ (.A1(net140),
    .A2(net136),
    .B1(_01748_),
    .C1(_01750_),
    .Y(_01754_));
 sky130_fd_sc_hd__a21o_1 _24854_ (.A1(_01748_),
    .A2(_01750_),
    .B1(_10546_),
    .X(_01755_));
 sky130_fd_sc_hd__o2bb2ai_4 _24855_ (.A1_N(_01562_),
    .A2_N(_01732_),
    .B1(_01749_),
    .B2(_01752_),
    .Y(_01756_));
 sky130_fd_sc_hd__o211ai_4 _24856_ (.A1(_01563_),
    .A2(_01730_),
    .B1(_01754_),
    .C1(_01755_),
    .Y(_01757_));
 sky130_fd_sc_hd__o21ai_1 _24857_ (.A1(_01751_),
    .A2(_01756_),
    .B1(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__and3_2 _24858_ (.A(_01758_),
    .B(net143),
    .C(_11743_),
    .X(_01759_));
 sky130_fd_sc_hd__nand2_1 _24859_ (.A(_01758_),
    .B(net132),
    .Y(_01760_));
 sky130_fd_sc_hd__o221ai_4 _24860_ (.A1(net141),
    .A2(_11742_),
    .B1(_01751_),
    .B2(_01756_),
    .C1(_01757_),
    .Y(_01761_));
 sky130_fd_sc_hd__a21oi_4 _24861_ (.A1(_01760_),
    .A2(_01761_),
    .B1(_01729_),
    .Y(_01762_));
 sky130_fd_sc_hd__a21o_1 _24862_ (.A1(_01760_),
    .A2(_01761_),
    .B1(_01729_),
    .X(_01763_));
 sky130_fd_sc_hd__nand2_2 _24863_ (.A(_01729_),
    .B(_01761_),
    .Y(_01765_));
 sky130_fd_sc_hd__a21oi_1 _24864_ (.A1(net132),
    .A2(_01758_),
    .B1(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__a31o_1 _24865_ (.A1(net143),
    .A2(_11743_),
    .A3(_01758_),
    .B1(_01765_),
    .X(_01767_));
 sky130_fd_sc_hd__o21ai_1 _24866_ (.A1(_01762_),
    .A2(_01766_),
    .B1(_00737_),
    .Y(_01768_));
 sky130_fd_sc_hd__o2111ai_4 _24867_ (.A1(_01765_),
    .A2(_01759_),
    .B1(_00367_),
    .C1(_00364_),
    .D1(_01763_),
    .Y(_01769_));
 sky130_fd_sc_hd__o221ai_4 _24868_ (.A1(net130),
    .A2(_00366_),
    .B1(_01759_),
    .B2(_01765_),
    .C1(_01763_),
    .Y(_01770_));
 sky130_fd_sc_hd__o21ai_2 _24869_ (.A1(_01762_),
    .A2(_01766_),
    .B1(_00736_),
    .Y(_01771_));
 sky130_fd_sc_hd__o21ai_1 _24870_ (.A1(_00737_),
    .A2(_01579_),
    .B1(_01582_),
    .Y(_01772_));
 sky130_fd_sc_hd__a21oi_2 _24871_ (.A1(_01580_),
    .A2(_00736_),
    .B1(_01581_),
    .Y(_01773_));
 sky130_fd_sc_hd__o2111a_1 _24872_ (.A1(_00737_),
    .A2(_01579_),
    .B1(_01582_),
    .C1(_01770_),
    .D1(_01771_),
    .X(_01774_));
 sky130_fd_sc_hd__nand3_2 _24873_ (.A(_01770_),
    .B(_01771_),
    .C(_01773_),
    .Y(_01776_));
 sky130_fd_sc_hd__nand3_4 _24874_ (.A(_01768_),
    .B(_01769_),
    .C(_01772_),
    .Y(_01777_));
 sky130_fd_sc_hd__a31o_1 _24875_ (.A1(_01332_),
    .A2(_01531_),
    .A3(_01532_),
    .B1(_01328_),
    .X(_01778_));
 sky130_fd_sc_hd__nor2_1 _24876_ (.A(_04223_),
    .B(_05465_),
    .Y(_01779_));
 sky130_fd_sc_hd__o311a_1 _24877_ (.A1(net244),
    .A2(net241),
    .A3(_07501_),
    .B1(_05462_),
    .C1(_07499_),
    .X(_01780_));
 sky130_fd_sc_hd__a31o_1 _24878_ (.A1(_07499_),
    .A2(_07503_),
    .A3(_05462_),
    .B1(_01779_),
    .X(_01781_));
 sky130_fd_sc_hd__or3_1 _24879_ (.A(net46),
    .B(_04245_),
    .C(_04124_),
    .X(_01782_));
 sky130_fd_sc_hd__o211ai_4 _24880_ (.A1(net170),
    .A2(_07765_),
    .B1(_05225_),
    .C1(_07771_),
    .Y(_01783_));
 sky130_fd_sc_hd__or3_2 _24881_ (.A(net45),
    .B(_04256_),
    .C(_04102_),
    .X(_01784_));
 sky130_fd_sc_hd__nand3_2 _24882_ (.A(net164),
    .B(_08208_),
    .C(net242),
    .Y(_01785_));
 sky130_fd_sc_hd__a22oi_2 _24883_ (.A1(_01782_),
    .A2(_01783_),
    .B1(_01784_),
    .B2(_01785_),
    .Y(_01787_));
 sky130_fd_sc_hd__a22o_1 _24884_ (.A1(_01782_),
    .A2(_01783_),
    .B1(_01784_),
    .B2(_01785_),
    .X(_01788_));
 sky130_fd_sc_hd__o2111a_1 _24885_ (.A1(_04245_),
    .A2(_05229_),
    .B1(_01783_),
    .C1(_01784_),
    .D1(_01785_),
    .X(_01789_));
 sky130_fd_sc_hd__o2111ai_4 _24886_ (.A1(_04245_),
    .A2(_05229_),
    .B1(_01783_),
    .C1(_01784_),
    .D1(_01785_),
    .Y(_01790_));
 sky130_fd_sc_hd__o211ai_2 _24887_ (.A1(_01779_),
    .A2(_01780_),
    .B1(_01788_),
    .C1(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__a21o_1 _24888_ (.A1(_01788_),
    .A2(_01790_),
    .B1(_01781_),
    .X(_01792_));
 sky130_fd_sc_hd__o21ai_1 _24889_ (.A1(_01787_),
    .A2(_01789_),
    .B1(_01781_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand3b_1 _24890_ (.A_N(_01781_),
    .B(_01788_),
    .C(_01790_),
    .Y(_01794_));
 sky130_fd_sc_hd__nand2_1 _24891_ (.A(_01793_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__nand2_1 _24892_ (.A(_01791_),
    .B(_01792_),
    .Y(_01796_));
 sky130_fd_sc_hd__and3_1 _24893_ (.A(_04102_),
    .B(net25),
    .C(net42),
    .X(_01798_));
 sky130_fd_sc_hd__a21oi_1 _24894_ (.A1(_08665_),
    .A2(_08668_),
    .B1(_04896_),
    .Y(_01799_));
 sky130_fd_sc_hd__a21oi_1 _24895_ (.A1(_08670_),
    .A2(_04895_),
    .B1(_01798_),
    .Y(_01800_));
 sky130_fd_sc_hd__o311a_2 _24896_ (.A1(net25),
    .A2(_04481_),
    .A3(_08207_),
    .B1(_01497_),
    .C1(_01493_),
    .X(_01801_));
 sky130_fd_sc_hd__o221ai_2 _24897_ (.A1(net319),
    .A2(_04483_),
    .B1(net150),
    .B2(_04481_),
    .C1(_01493_),
    .Y(_01802_));
 sky130_fd_sc_hd__o2111ai_2 _24898_ (.A1(_04481_),
    .A2(_08665_),
    .B1(_01493_),
    .C1(_01497_),
    .D1(_01800_),
    .Y(_01803_));
 sky130_fd_sc_hd__o21ai_1 _24899_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01802_),
    .Y(_01804_));
 sky130_fd_sc_hd__nand2_1 _24900_ (.A(_01800_),
    .B(_01802_),
    .Y(_01805_));
 sky130_fd_sc_hd__o21ai_2 _24901_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01801_),
    .Y(_01806_));
 sky130_fd_sc_hd__o21ai_2 _24902_ (.A1(_01493_),
    .A2(_01498_),
    .B1(_01491_),
    .Y(_01807_));
 sky130_fd_sc_hd__a22oi_4 _24903_ (.A1(_01803_),
    .A2(_01804_),
    .B1(_01807_),
    .B2(_01503_),
    .Y(_01809_));
 sky130_fd_sc_hd__nand4_1 _24904_ (.A(_01500_),
    .B(_01506_),
    .C(_01805_),
    .D(_01806_),
    .Y(_01810_));
 sky130_fd_sc_hd__a2bb2oi_4 _24905_ (.A1_N(_01499_),
    .A2_N(_01505_),
    .B1(_01805_),
    .B2(_01806_),
    .Y(_01811_));
 sky130_fd_sc_hd__nor3_2 _24906_ (.A(_01811_),
    .B(_01796_),
    .C(_01809_),
    .Y(_01812_));
 sky130_fd_sc_hd__a211o_2 _24907_ (.A1(_01793_),
    .A2(_01794_),
    .B1(_01809_),
    .C1(_01811_),
    .X(_01813_));
 sky130_fd_sc_hd__o2bb2a_1 _24908_ (.A1_N(_01791_),
    .A2_N(_01792_),
    .B1(_01809_),
    .B2(_01811_),
    .X(_01814_));
 sky130_fd_sc_hd__o21ai_2 _24909_ (.A1(_01809_),
    .A2(_01811_),
    .B1(_01796_),
    .Y(_01815_));
 sky130_fd_sc_hd__o211ai_4 _24910_ (.A1(_00796_),
    .A2(_01324_),
    .B1(_01813_),
    .C1(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__o21ai_2 _24911_ (.A1(_01812_),
    .A2(_01814_),
    .B1(_01331_),
    .Y(_01817_));
 sky130_fd_sc_hd__o2bb2ai_4 _24912_ (.A1_N(_01816_),
    .A2_N(_01817_),
    .B1(_11741_),
    .B2(_00360_),
    .Y(_01818_));
 sky130_fd_sc_hd__inv_2 _24913_ (.A(_01818_),
    .Y(_01820_));
 sky130_fd_sc_hd__o2111ai_4 _24914_ (.A1(_13066_),
    .A2(_00357_),
    .B1(_11740_),
    .C1(_01816_),
    .D1(_01817_),
    .Y(_01821_));
 sky130_fd_sc_hd__inv_2 _24915_ (.A(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21o_1 _24916_ (.A1(_01818_),
    .A2(_01821_),
    .B1(_01778_),
    .X(_01823_));
 sky130_fd_sc_hd__inv_2 _24917_ (.A(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__o21ai_4 _24918_ (.A1(_01328_),
    .A2(_01533_),
    .B1(_01818_),
    .Y(_01825_));
 sky130_fd_sc_hd__and3_1 _24919_ (.A(_01778_),
    .B(_01818_),
    .C(_01821_),
    .X(_01826_));
 sky130_fd_sc_hd__o22a_1 _24920_ (.A1(_01328_),
    .A2(_01533_),
    .B1(_01820_),
    .B2(_01822_),
    .X(_01827_));
 sky130_fd_sc_hd__and4_1 _24921_ (.A(_01329_),
    .B(_01535_),
    .C(_01818_),
    .D(_01821_),
    .X(_01828_));
 sky130_fd_sc_hd__o21ai_4 _24922_ (.A1(_01822_),
    .A2(_01825_),
    .B1(_01823_),
    .Y(_01829_));
 sky130_fd_sc_hd__o2bb2ai_1 _24923_ (.A1_N(_01776_),
    .A2_N(_01777_),
    .B1(_01824_),
    .B2(_01826_),
    .Y(_01831_));
 sky130_fd_sc_hd__o2111ai_2 _24924_ (.A1(_01822_),
    .A2(_01825_),
    .B1(_01823_),
    .C1(_01776_),
    .D1(_01777_),
    .Y(_01832_));
 sky130_fd_sc_hd__nand3_1 _24925_ (.A(_01776_),
    .B(_01777_),
    .C(_01829_),
    .Y(_01833_));
 sky130_fd_sc_hd__o2bb2ai_2 _24926_ (.A1_N(_01776_),
    .A2_N(_01777_),
    .B1(_01827_),
    .B2(_01828_),
    .Y(_01834_));
 sky130_fd_sc_hd__nand2_1 _24927_ (.A(_01831_),
    .B(_01832_),
    .Y(_01835_));
 sky130_fd_sc_hd__o22a_1 _24928_ (.A1(_01585_),
    .A2(_01591_),
    .B1(_01588_),
    .B2(_01546_),
    .X(_01836_));
 sky130_fd_sc_hd__o22ai_1 _24929_ (.A1(_01585_),
    .A2(_01591_),
    .B1(_01588_),
    .B2(_01546_),
    .Y(_01837_));
 sky130_fd_sc_hd__and3_1 _24930_ (.A(_01836_),
    .B(_01834_),
    .C(_01833_),
    .X(_01838_));
 sky130_fd_sc_hd__o2111ai_4 _24931_ (.A1(_01546_),
    .A2(_01588_),
    .B1(_01593_),
    .C1(_01833_),
    .D1(_01834_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand3_1 _24932_ (.A(_01831_),
    .B(_01832_),
    .C(_01837_),
    .Y(_01840_));
 sky130_fd_sc_hd__nand2_1 _24933_ (.A(_01839_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o31a_1 _24934_ (.A1(_00364_),
    .A2(_01533_),
    .A3(_01536_),
    .B1(_01543_),
    .X(_01842_));
 sky130_fd_sc_hd__a31o_1 _24935_ (.A1(net130),
    .A2(_01535_),
    .A3(_01537_),
    .B1(_01542_),
    .X(_01843_));
 sky130_fd_sc_hd__o2bb2a_2 _24936_ (.A1_N(_05076_),
    .A2_N(net238),
    .B1(_08007_),
    .B2(_04113_),
    .X(_01844_));
 sky130_fd_sc_hd__and3b_1 _24937_ (.A_N(net54),
    .B(net53),
    .C(net14),
    .X(_01845_));
 sky130_fd_sc_hd__and3_1 _24938_ (.A(_05290_),
    .B(_05292_),
    .C(_07642_),
    .X(_01846_));
 sky130_fd_sc_hd__a31o_1 _24939_ (.A1(_05290_),
    .A2(_05292_),
    .A3(_07642_),
    .B1(_01845_),
    .X(_01847_));
 sky130_fd_sc_hd__a32oi_2 _24940_ (.A1(net178),
    .A2(_05553_),
    .A3(net239),
    .B1(_07308_),
    .B2(net15),
    .Y(_01848_));
 sky130_fd_sc_hd__a32o_1 _24941_ (.A1(net178),
    .A2(_05553_),
    .A3(net239),
    .B1(_07308_),
    .B2(net15),
    .X(_01849_));
 sky130_fd_sc_hd__nor2_1 _24942_ (.A(_04168_),
    .B(_06866_),
    .Y(_01850_));
 sky130_fd_sc_hd__o311a_2 _24943_ (.A1(_05551_),
    .A2(_05925_),
    .A3(_06220_),
    .B1(_06863_),
    .C1(_06219_),
    .X(_01852_));
 sky130_fd_sc_hd__a31oi_2 _24944_ (.A1(net202),
    .A2(net173),
    .A3(net240),
    .B1(_01850_),
    .Y(_01853_));
 sky130_fd_sc_hd__or3b_2 _24945_ (.A(_04157_),
    .B(net52),
    .C_N(net51),
    .X(_01854_));
 sky130_fd_sc_hd__o31ai_2 _24946_ (.A1(net204),
    .A2(_07224_),
    .A3(_05932_),
    .B1(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__o21ai_4 _24947_ (.A1(_01850_),
    .A2(_01852_),
    .B1(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__o211a_1 _24948_ (.A1(_05935_),
    .A2(_07224_),
    .B1(_01853_),
    .C1(_01854_),
    .X(_01857_));
 sky130_fd_sc_hd__o211ai_4 _24949_ (.A1(_05935_),
    .A2(_07224_),
    .B1(_01853_),
    .C1(_01854_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand3_2 _24950_ (.A(_01849_),
    .B(_01856_),
    .C(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__a21o_1 _24951_ (.A1(_01856_),
    .A2(_01858_),
    .B1(_01849_),
    .X(_01860_));
 sky130_fd_sc_hd__a21o_1 _24952_ (.A1(_01856_),
    .A2(_01858_),
    .B1(_01848_),
    .X(_01861_));
 sky130_fd_sc_hd__nand3_1 _24953_ (.A(_01848_),
    .B(_01856_),
    .C(_01858_),
    .Y(_01863_));
 sky130_fd_sc_hd__a21o_1 _24954_ (.A1(_01650_),
    .A2(_01661_),
    .B1(_01659_),
    .X(_01864_));
 sky130_fd_sc_hd__a21oi_1 _24955_ (.A1(_01650_),
    .A2(_01661_),
    .B1(_01659_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand3_2 _24956_ (.A(_01864_),
    .B(_01860_),
    .C(_01859_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand3_2 _24957_ (.A(_01861_),
    .B(_01863_),
    .C(_01865_),
    .Y(_01867_));
 sky130_fd_sc_hd__a221o_2 _24958_ (.A1(net14),
    .A2(_07643_),
    .B1(_01866_),
    .B2(_01867_),
    .C1(_01846_),
    .X(_01868_));
 sky130_fd_sc_hd__o211ai_4 _24959_ (.A1(_01845_),
    .A2(_01846_),
    .B1(_01866_),
    .C1(_01867_),
    .Y(_01869_));
 sky130_fd_sc_hd__a32oi_4 _24960_ (.A1(_01648_),
    .A2(_01664_),
    .A3(_01665_),
    .B1(_01667_),
    .B2(_01647_),
    .Y(_01870_));
 sky130_fd_sc_hd__a21o_1 _24961_ (.A1(_01868_),
    .A2(_01869_),
    .B1(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__nand3_4 _24962_ (.A(_01868_),
    .B(_01869_),
    .C(_01870_),
    .Y(_01872_));
 sky130_fd_sc_hd__inv_2 _24963_ (.A(_01872_),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2_1 _24964_ (.A(_01871_),
    .B(_01872_),
    .Y(_01875_));
 sky130_fd_sc_hd__nor2_2 _24965_ (.A(_01844_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__a31o_1 _24966_ (.A1(_01868_),
    .A2(_01869_),
    .A3(_01870_),
    .B1(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__o21a_1 _24967_ (.A1(_01844_),
    .A2(_01875_),
    .B1(_01872_),
    .X(_01878_));
 sky130_fd_sc_hd__a21oi_2 _24968_ (.A1(_01871_),
    .A2(_01872_),
    .B1(_01844_),
    .Y(_01879_));
 sky130_fd_sc_hd__and3_1 _24969_ (.A(_01871_),
    .B(_01872_),
    .C(_01844_),
    .X(_01880_));
 sky130_fd_sc_hd__a21boi_2 _24970_ (.A1(_01871_),
    .A2(_01872_),
    .B1_N(_01844_),
    .Y(_01881_));
 sky130_fd_sc_hd__a21boi_4 _24971_ (.A1(_01635_),
    .A2(_01638_),
    .B1_N(_01636_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21oi_1 _24972_ (.A1(_01609_),
    .A2(_01618_),
    .B1(_01616_),
    .Y(_01883_));
 sky130_fd_sc_hd__a32o_1 _24973_ (.A1(net197),
    .A2(_06452_),
    .A3(net273),
    .B1(_06326_),
    .B2(net18),
    .X(_01885_));
 sky130_fd_sc_hd__or3b_1 _24974_ (.A(net48),
    .B(_04212_),
    .C_N(net47),
    .X(_01886_));
 sky130_fd_sc_hd__o211ai_4 _24975_ (.A1(net176),
    .A2(_07074_),
    .B1(_05762_),
    .C1(_07072_),
    .Y(_01887_));
 sky130_fd_sc_hd__nor2_1 _24976_ (.A(_04201_),
    .B(_06030_),
    .Y(_01888_));
 sky130_fd_sc_hd__or3b_1 _24977_ (.A(net49),
    .B(_04201_),
    .C_N(net48),
    .X(_01889_));
 sky130_fd_sc_hd__o311a_1 _24978_ (.A1(net244),
    .A2(net241),
    .A3(_06759_),
    .B1(net274),
    .C1(net192),
    .X(_01890_));
 sky130_fd_sc_hd__o211ai_2 _24979_ (.A1(net176),
    .A2(_06759_),
    .B1(net274),
    .C1(net192),
    .Y(_01891_));
 sky130_fd_sc_hd__o2bb2a_1 _24980_ (.A1_N(_01886_),
    .A2_N(_01887_),
    .B1(_01888_),
    .B2(_01890_),
    .X(_01892_));
 sky130_fd_sc_hd__o2bb2ai_2 _24981_ (.A1_N(_01886_),
    .A2_N(_01887_),
    .B1(_01888_),
    .B2(_01890_),
    .Y(_01893_));
 sky130_fd_sc_hd__o2111ai_4 _24982_ (.A1(_04212_),
    .A2(_05766_),
    .B1(_01887_),
    .C1(_01889_),
    .D1(_01891_),
    .Y(_01894_));
 sky130_fd_sc_hd__and3_1 _24983_ (.A(_01885_),
    .B(_01893_),
    .C(_01894_),
    .X(_01896_));
 sky130_fd_sc_hd__nand3_2 _24984_ (.A(_01885_),
    .B(_01893_),
    .C(_01894_),
    .Y(_01897_));
 sky130_fd_sc_hd__a21o_1 _24985_ (.A1(_01893_),
    .A2(_01894_),
    .B1(_01885_),
    .X(_01898_));
 sky130_fd_sc_hd__a21bo_1 _24986_ (.A1(_01893_),
    .A2(_01894_),
    .B1_N(_01885_),
    .X(_01899_));
 sky130_fd_sc_hd__nand3b_1 _24987_ (.A_N(_01885_),
    .B(_01893_),
    .C(_01894_),
    .Y(_01900_));
 sky130_fd_sc_hd__a21o_1 _24988_ (.A1(_01517_),
    .A2(_01525_),
    .B1(_01522_),
    .X(_01901_));
 sky130_fd_sc_hd__a21oi_1 _24989_ (.A1(_01517_),
    .A2(_01525_),
    .B1(_01522_),
    .Y(_01902_));
 sky130_fd_sc_hd__and3_1 _24990_ (.A(_01899_),
    .B(_01900_),
    .C(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__nand3_2 _24991_ (.A(_01899_),
    .B(_01900_),
    .C(_01902_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand3_4 _24992_ (.A(_01897_),
    .B(_01898_),
    .C(_01901_),
    .Y(_01905_));
 sky130_fd_sc_hd__inv_2 _24993_ (.A(_01905_),
    .Y(_01907_));
 sky130_fd_sc_hd__a21boi_4 _24994_ (.A1(_01904_),
    .A2(_01905_),
    .B1_N(_01883_),
    .Y(_01908_));
 sky130_fd_sc_hd__a21bo_1 _24995_ (.A1(_01904_),
    .A2(_01905_),
    .B1_N(_01883_),
    .X(_01909_));
 sky130_fd_sc_hd__o211a_2 _24996_ (.A1(_01616_),
    .A2(_01621_),
    .B1(_01904_),
    .C1(_01905_),
    .X(_01910_));
 sky130_fd_sc_hd__o211ai_1 _24997_ (.A1(_01616_),
    .A2(_01621_),
    .B1(_01904_),
    .C1(_01905_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_1 _24998_ (.A(_01909_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__a21oi_4 _24999_ (.A1(_01515_),
    .A2(_01530_),
    .B1(_01513_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor3_4 _25000_ (.A(_01908_),
    .B(_01910_),
    .C(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__a211o_1 _25001_ (.A1(_01514_),
    .A2(_01531_),
    .B1(_01908_),
    .C1(_01910_),
    .X(_01915_));
 sky130_fd_sc_hd__o21a_2 _25002_ (.A1(_01908_),
    .A2(_01910_),
    .B1(_01913_),
    .X(_01916_));
 sky130_fd_sc_hd__o21ai_1 _25003_ (.A1(_01908_),
    .A2(_01910_),
    .B1(_01913_),
    .Y(_01918_));
 sky130_fd_sc_hd__o21a_2 _25004_ (.A1(_01606_),
    .A2(_01626_),
    .B1(_01628_),
    .X(_01919_));
 sky130_fd_sc_hd__a21oi_2 _25005_ (.A1(_01912_),
    .A2(_01913_),
    .B1(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__a211o_1 _25006_ (.A1(_01912_),
    .A2(_01913_),
    .B1(_01919_),
    .C1(_01914_),
    .X(_01921_));
 sky130_fd_sc_hd__o21ai_1 _25007_ (.A1(_01914_),
    .A2(_01916_),
    .B1(_01919_),
    .Y(_01922_));
 sky130_fd_sc_hd__o21bai_4 _25008_ (.A1(_01914_),
    .A2(_01916_),
    .B1_N(_01919_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand3_2 _25009_ (.A(_01915_),
    .B(_01918_),
    .C(_01919_),
    .Y(_01924_));
 sky130_fd_sc_hd__a21oi_4 _25010_ (.A1(_01923_),
    .A2(_01924_),
    .B1(_01882_),
    .Y(_01925_));
 sky130_fd_sc_hd__a21o_1 _25011_ (.A1(_01923_),
    .A2(_01924_),
    .B1(_01882_),
    .X(_01926_));
 sky130_fd_sc_hd__a21boi_4 _25012_ (.A1(_01921_),
    .A2(_01922_),
    .B1_N(_01882_),
    .Y(_01927_));
 sky130_fd_sc_hd__nand3_2 _25013_ (.A(_01882_),
    .B(_01923_),
    .C(_01924_),
    .Y(_01929_));
 sky130_fd_sc_hd__o21a_1 _25014_ (.A1(_01876_),
    .A2(_01881_),
    .B1(_01926_),
    .X(_01930_));
 sky130_fd_sc_hd__o21ai_2 _25015_ (.A1(_01879_),
    .A2(_01880_),
    .B1(_01929_),
    .Y(_01931_));
 sky130_fd_sc_hd__o31a_1 _25016_ (.A1(_01876_),
    .A2(_01881_),
    .A3(_01927_),
    .B1(_01926_),
    .X(_01932_));
 sky130_fd_sc_hd__o211ai_2 _25017_ (.A1(_01876_),
    .A2(_01881_),
    .B1(_01926_),
    .C1(_01929_),
    .Y(_01933_));
 sky130_fd_sc_hd__o22ai_2 _25018_ (.A1(_01879_),
    .A2(_01880_),
    .B1(_01925_),
    .B2(_01927_),
    .Y(_01934_));
 sky130_fd_sc_hd__o22ai_2 _25019_ (.A1(_01876_),
    .A2(_01881_),
    .B1(_01925_),
    .B2(_01927_),
    .Y(_01935_));
 sky130_fd_sc_hd__and3_1 _25020_ (.A(_01934_),
    .B(_01842_),
    .C(_01933_),
    .X(_01936_));
 sky130_fd_sc_hd__nand3_2 _25021_ (.A(_01934_),
    .B(_01842_),
    .C(_01933_),
    .Y(_01937_));
 sky130_fd_sc_hd__o211ai_4 _25022_ (.A1(_01925_),
    .A2(_01931_),
    .B1(_01935_),
    .C1(_01843_),
    .Y(_01938_));
 sky130_fd_sc_hd__nor2_1 _25023_ (.A(_01641_),
    .B(_01678_),
    .Y(_01940_));
 sky130_fd_sc_hd__o2bb2ai_2 _25024_ (.A1_N(_01937_),
    .A2_N(_01938_),
    .B1(_01940_),
    .B2(_01680_),
    .Y(_01941_));
 sky130_fd_sc_hd__o2111ai_4 _25025_ (.A1(_01641_),
    .A2(_01678_),
    .B1(_01681_),
    .C1(_01937_),
    .D1(_01938_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _25026_ (.A(_01941_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__a22o_1 _25027_ (.A1(_01839_),
    .A2(_01840_),
    .B1(_01941_),
    .B2(_01942_),
    .X(_01944_));
 sky130_fd_sc_hd__nand3_1 _25028_ (.A(_01839_),
    .B(_01941_),
    .C(_01942_),
    .Y(_01945_));
 sky130_fd_sc_hd__nand3_1 _25029_ (.A(_01840_),
    .B(_01941_),
    .C(_01942_),
    .Y(_01946_));
 sky130_fd_sc_hd__nand3_1 _25030_ (.A(_01839_),
    .B(_01840_),
    .C(_01943_),
    .Y(_01947_));
 sky130_fd_sc_hd__nand3_1 _25031_ (.A(_01841_),
    .B(_01941_),
    .C(_01942_),
    .Y(_01948_));
 sky130_fd_sc_hd__a31oi_1 _25032_ (.A1(_01602_),
    .A2(_01693_),
    .A3(_01694_),
    .B1(_01603_),
    .Y(_01949_));
 sky130_fd_sc_hd__o221a_1 _25033_ (.A1(_01838_),
    .A2(_01946_),
    .B1(_01603_),
    .B2(_01700_),
    .C1(_01944_),
    .X(_01951_));
 sky130_fd_sc_hd__o221ai_2 _25034_ (.A1(_01838_),
    .A2(_01946_),
    .B1(_01603_),
    .B2(_01700_),
    .C1(_01944_),
    .Y(_01952_));
 sky130_fd_sc_hd__nand3_1 _25035_ (.A(_01947_),
    .B(_01948_),
    .C(_01949_),
    .Y(_01953_));
 sky130_fd_sc_hd__a32oi_2 _25036_ (.A1(_01684_),
    .A2(_01685_),
    .A3(_01686_),
    .B1(_01689_),
    .B2(_01690_),
    .Y(_01954_));
 sky130_fd_sc_hd__a32o_1 _25037_ (.A1(_01684_),
    .A2(_01685_),
    .A3(_01686_),
    .B1(_01689_),
    .B2(_01690_),
    .X(_01955_));
 sky130_fd_sc_hd__a21o_1 _25038_ (.A1(_01952_),
    .A2(_01953_),
    .B1(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__nand3_1 _25039_ (.A(_01952_),
    .B(_01953_),
    .C(_01955_),
    .Y(_01957_));
 sky130_fd_sc_hd__a21o_1 _25040_ (.A1(_01952_),
    .A2(_01953_),
    .B1(_01954_),
    .X(_01958_));
 sky130_fd_sc_hd__a31o_1 _25041_ (.A1(_01947_),
    .A2(_01948_),
    .A3(_01949_),
    .B1(_01955_),
    .X(_01959_));
 sky130_fd_sc_hd__o211a_1 _25042_ (.A1(_01951_),
    .A2(_01959_),
    .B1(_01958_),
    .C1(_01727_),
    .X(_01960_));
 sky130_fd_sc_hd__o211ai_1 _25043_ (.A1(_01951_),
    .A2(_01959_),
    .B1(_01958_),
    .C1(_01727_),
    .Y(_01962_));
 sky130_fd_sc_hd__nand3_1 _25044_ (.A(_01728_),
    .B(_01956_),
    .C(_01957_),
    .Y(_01963_));
 sky130_fd_sc_hd__o21bai_2 _25045_ (.A1(_01643_),
    .A2(_01675_),
    .B1_N(_01674_),
    .Y(_01964_));
 sky130_fd_sc_hd__a21o_1 _25046_ (.A1(_01962_),
    .A2(_01963_),
    .B1(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__nand3_1 _25047_ (.A(_01962_),
    .B(_01963_),
    .C(_01964_),
    .Y(_01966_));
 sky130_fd_sc_hd__a21o_1 _25048_ (.A1(_01965_),
    .A2(_01966_),
    .B1(_01726_),
    .X(_01967_));
 sky130_fd_sc_hd__inv_2 _25049_ (.A(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand3_1 _25050_ (.A(_01726_),
    .B(_01965_),
    .C(_01966_),
    .Y(_01969_));
 sky130_fd_sc_hd__nand2_1 _25051_ (.A(_01967_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__xor2_1 _25052_ (.A(_01725_),
    .B(_01970_),
    .X(net110));
 sky130_fd_sc_hd__a21o_1 _25053_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01960_),
    .X(_01972_));
 sky130_fd_sc_hd__a21oi_1 _25054_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01960_),
    .Y(_01973_));
 sky130_fd_sc_hd__a21o_1 _25055_ (.A1(_01953_),
    .A2(_01954_),
    .B1(_01951_),
    .X(_01974_));
 sky130_fd_sc_hd__o21a_1 _25056_ (.A1(_01680_),
    .A2(_01940_),
    .B1(_01938_),
    .X(_01975_));
 sky130_fd_sc_hd__nor2_1 _25057_ (.A(_01936_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__a31o_1 _25058_ (.A1(_01842_),
    .A2(_01933_),
    .A3(_01934_),
    .B1(_01975_),
    .X(_01977_));
 sky130_fd_sc_hd__o21ai_2 _25059_ (.A1(_01835_),
    .A2(_01836_),
    .B1(_01945_),
    .Y(_01978_));
 sky130_fd_sc_hd__and3_1 _25060_ (.A(_01329_),
    .B(_01535_),
    .C(_01821_),
    .X(_01979_));
 sky130_fd_sc_hd__a21o_1 _25061_ (.A1(_01778_),
    .A2(_01818_),
    .B1(_01822_),
    .X(_01980_));
 sky130_fd_sc_hd__a32oi_2 _25062_ (.A1(_05290_),
    .A2(_05292_),
    .A3(net238),
    .B1(_08006_),
    .B2(net14),
    .Y(_01981_));
 sky130_fd_sc_hd__a32o_1 _25063_ (.A1(_05290_),
    .A2(_05292_),
    .A3(net238),
    .B1(_08006_),
    .B2(net14),
    .X(_01983_));
 sky130_fd_sc_hd__o311a_1 _25064_ (.A1(net233),
    .A2(_04787_),
    .A3(_05551_),
    .B1(_07642_),
    .C1(net178),
    .X(_01984_));
 sky130_fd_sc_hd__and3b_1 _25065_ (.A_N(net54),
    .B(net53),
    .C(net15),
    .X(_01985_));
 sky130_fd_sc_hd__a31o_1 _25066_ (.A1(net178),
    .A2(_05553_),
    .A3(_07642_),
    .B1(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__o21ai_1 _25067_ (.A1(_01848_),
    .A2(_01857_),
    .B1(_01856_),
    .Y(_01987_));
 sky130_fd_sc_hd__a22oi_2 _25068_ (.A1(_05934_),
    .A2(net239),
    .B1(_07308_),
    .B2(net16),
    .Y(_01988_));
 sky130_fd_sc_hd__a32o_1 _25069_ (.A1(net176),
    .A2(_05933_),
    .A3(net239),
    .B1(_07308_),
    .B2(net16),
    .X(_01989_));
 sky130_fd_sc_hd__a32oi_4 _25070_ (.A1(net202),
    .A2(net173),
    .A3(net269),
    .B1(_07225_),
    .B2(net17),
    .Y(_01990_));
 sky130_fd_sc_hd__or3_1 _25071_ (.A(net51),
    .B(_04190_),
    .C(_04179_),
    .X(_01991_));
 sky130_fd_sc_hd__nand3_1 _25072_ (.A(net197),
    .B(_06452_),
    .C(net240),
    .Y(_01992_));
 sky130_fd_sc_hd__a21oi_1 _25073_ (.A1(_01991_),
    .A2(_01992_),
    .B1(_01990_),
    .Y(_01994_));
 sky130_fd_sc_hd__a21o_1 _25074_ (.A1(_01991_),
    .A2(_01992_),
    .B1(_01990_),
    .X(_01995_));
 sky130_fd_sc_hd__o311a_1 _25075_ (.A1(_04179_),
    .A2(_04190_),
    .A3(net51),
    .B1(_01992_),
    .C1(_01990_),
    .X(_01996_));
 sky130_fd_sc_hd__o221ai_2 _25076_ (.A1(_06454_),
    .A2(_06864_),
    .B1(_06866_),
    .B2(_04179_),
    .C1(_01990_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand3_1 _25077_ (.A(_01989_),
    .B(_01995_),
    .C(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__o21ai_1 _25078_ (.A1(_01994_),
    .A2(_01996_),
    .B1(_01988_),
    .Y(_01999_));
 sky130_fd_sc_hd__o21ai_1 _25079_ (.A1(_01994_),
    .A2(_01996_),
    .B1(_01989_),
    .Y(_02000_));
 sky130_fd_sc_hd__nand3_1 _25080_ (.A(_01988_),
    .B(_01995_),
    .C(_01997_),
    .Y(_02001_));
 sky130_fd_sc_hd__nand4_4 _25081_ (.A(_01856_),
    .B(_01859_),
    .C(_02000_),
    .D(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__nand3_2 _25082_ (.A(_01987_),
    .B(_01998_),
    .C(_01999_),
    .Y(_02003_));
 sky130_fd_sc_hd__a21oi_1 _25083_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_01986_),
    .Y(_02005_));
 sky130_fd_sc_hd__a21o_1 _25084_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_01986_),
    .X(_02006_));
 sky130_fd_sc_hd__o211a_1 _25085_ (.A1(_01984_),
    .A2(_01985_),
    .B1(_02002_),
    .C1(_02003_),
    .X(_02007_));
 sky130_fd_sc_hd__o211ai_1 _25086_ (.A1(_01984_),
    .A2(_01985_),
    .B1(_02002_),
    .C1(_02003_),
    .Y(_02008_));
 sky130_fd_sc_hd__a32o_1 _25087_ (.A1(_01859_),
    .A2(_01860_),
    .A3(_01864_),
    .B1(_01867_),
    .B2(_01847_),
    .X(_02009_));
 sky130_fd_sc_hd__a32oi_2 _25088_ (.A1(_01859_),
    .A2(_01860_),
    .A3(_01864_),
    .B1(_01867_),
    .B2(_01847_),
    .Y(_02010_));
 sky130_fd_sc_hd__a21oi_1 _25089_ (.A1(_02006_),
    .A2(_02008_),
    .B1(_02009_),
    .Y(_02011_));
 sky130_fd_sc_hd__o21ai_1 _25090_ (.A1(_02005_),
    .A2(_02007_),
    .B1(_02010_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor3_2 _25091_ (.A(_02005_),
    .B(_02007_),
    .C(_02010_),
    .Y(_02013_));
 sky130_fd_sc_hd__o21a_1 _25092_ (.A1(_02011_),
    .A2(_02013_),
    .B1(_01981_),
    .X(_02014_));
 sky130_fd_sc_hd__o21ai_1 _25093_ (.A1(_02011_),
    .A2(_02013_),
    .B1(_01981_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_1 _25094_ (.A(_01983_),
    .B(_02012_),
    .Y(_02017_));
 sky130_fd_sc_hd__nor2_1 _25095_ (.A(_02013_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__o21a_1 _25096_ (.A1(_02013_),
    .A2(_02017_),
    .B1(_02016_),
    .X(_02019_));
 sky130_fd_sc_hd__o21ai_1 _25097_ (.A1(_02013_),
    .A2(_02017_),
    .B1(_02016_),
    .Y(_02020_));
 sky130_fd_sc_hd__o31a_1 _25098_ (.A1(_01908_),
    .A2(_01910_),
    .A3(_01913_),
    .B1(_01919_),
    .X(_02021_));
 sky130_fd_sc_hd__o21ai_2 _25099_ (.A1(_01919_),
    .A2(_01916_),
    .B1(_01915_),
    .Y(_02022_));
 sky130_fd_sc_hd__a311oi_2 _25100_ (.A1(_01901_),
    .A2(_01898_),
    .A3(_01897_),
    .B1(_01616_),
    .C1(_01621_),
    .Y(_02023_));
 sky130_fd_sc_hd__o21a_1 _25101_ (.A1(_01616_),
    .A2(_01621_),
    .B1(_01904_),
    .X(_02024_));
 sky130_fd_sc_hd__a31o_1 _25102_ (.A1(_01899_),
    .A2(_01900_),
    .A3(_01902_),
    .B1(_02023_),
    .X(_02025_));
 sky130_fd_sc_hd__a21oi_2 _25103_ (.A1(_01791_),
    .A2(_01792_),
    .B1(_01811_),
    .Y(_02027_));
 sky130_fd_sc_hd__a21o_1 _25104_ (.A1(_01810_),
    .A2(_01795_),
    .B1(_01811_),
    .X(_02028_));
 sky130_fd_sc_hd__a21o_1 _25105_ (.A1(_01885_),
    .A2(_01894_),
    .B1(_01892_),
    .X(_02029_));
 sky130_fd_sc_hd__nor2_1 _25106_ (.A(_01781_),
    .B(_01787_),
    .Y(_02030_));
 sky130_fd_sc_hd__o21ai_1 _25107_ (.A1(_01779_),
    .A2(_01780_),
    .B1(_01790_),
    .Y(_02031_));
 sky130_fd_sc_hd__a21o_1 _25108_ (.A1(_01781_),
    .A2(_01790_),
    .B1(_01787_),
    .X(_02032_));
 sky130_fd_sc_hd__o311a_1 _25109_ (.A1(net244),
    .A2(net241),
    .A3(_06759_),
    .B1(net273),
    .C1(net192),
    .X(_02033_));
 sky130_fd_sc_hd__and3_1 _25110_ (.A(_04190_),
    .B(net19),
    .C(net49),
    .X(_02034_));
 sky130_fd_sc_hd__o2bb2a_2 _25111_ (.A1_N(net19),
    .A2_N(_06326_),
    .B1(_06764_),
    .B2(_06325_),
    .X(_02035_));
 sky130_fd_sc_hd__a31o_1 _25112_ (.A1(net192),
    .A2(_06762_),
    .A3(net273),
    .B1(_02034_),
    .X(_02036_));
 sky130_fd_sc_hd__or3b_2 _25113_ (.A(net49),
    .B(_04212_),
    .C_N(net48),
    .X(_02038_));
 sky130_fd_sc_hd__o221ai_4 _25114_ (.A1(net176),
    .A2(_07074_),
    .B1(_04212_),
    .B2(net190),
    .C1(net274),
    .Y(_02039_));
 sky130_fd_sc_hd__nor2_1 _25115_ (.A(_04223_),
    .B(_05766_),
    .Y(_02040_));
 sky130_fd_sc_hd__or3b_1 _25116_ (.A(net48),
    .B(_04223_),
    .C_N(net47),
    .X(_02041_));
 sky130_fd_sc_hd__a211oi_2 _25117_ (.A1(net204),
    .A2(_07500_),
    .B1(_05763_),
    .C1(_07498_),
    .Y(_02042_));
 sky130_fd_sc_hd__o211ai_2 _25118_ (.A1(net176),
    .A2(_07501_),
    .B1(_05762_),
    .C1(_07499_),
    .Y(_02043_));
 sky130_fd_sc_hd__o2bb2ai_4 _25119_ (.A1_N(_02038_),
    .A2_N(_02039_),
    .B1(_02040_),
    .B2(_02042_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand4_4 _25120_ (.A(_02038_),
    .B(_02039_),
    .C(_02041_),
    .D(_02043_),
    .Y(_02045_));
 sky130_fd_sc_hd__nand2_1 _25121_ (.A(_02044_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__a21oi_4 _25122_ (.A1(_02044_),
    .A2(_02045_),
    .B1(_02036_),
    .Y(_02047_));
 sky130_fd_sc_hd__a21o_1 _25123_ (.A1(_02044_),
    .A2(_02045_),
    .B1(_02036_),
    .X(_02049_));
 sky130_fd_sc_hd__o211a_1 _25124_ (.A1(_02033_),
    .A2(_02034_),
    .B1(_02044_),
    .C1(_02045_),
    .X(_02050_));
 sky130_fd_sc_hd__o211ai_2 _25125_ (.A1(_02033_),
    .A2(_02034_),
    .B1(_02044_),
    .C1(_02045_),
    .Y(_02051_));
 sky130_fd_sc_hd__o2bb2ai_2 _25126_ (.A1_N(_01788_),
    .A2_N(_02031_),
    .B1(_02035_),
    .B2(_02046_),
    .Y(_02052_));
 sky130_fd_sc_hd__nand3_2 _25127_ (.A(_02032_),
    .B(_02049_),
    .C(_02051_),
    .Y(_02053_));
 sky130_fd_sc_hd__o22ai_4 _25128_ (.A1(_01789_),
    .A2(_02030_),
    .B1(_02047_),
    .B2(_02050_),
    .Y(_02054_));
 sky130_fd_sc_hd__o221a_1 _25129_ (.A1(_01892_),
    .A2(_01896_),
    .B1(_02047_),
    .B2(_02052_),
    .C1(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__o221ai_4 _25130_ (.A1(_01892_),
    .A2(_01896_),
    .B1(_02047_),
    .B2(_02052_),
    .C1(_02054_),
    .Y(_02056_));
 sky130_fd_sc_hd__a21oi_2 _25131_ (.A1(_02053_),
    .A2(_02054_),
    .B1(_02029_),
    .Y(_02057_));
 sky130_fd_sc_hd__a21o_1 _25132_ (.A1(_02053_),
    .A2(_02054_),
    .B1(_02029_),
    .X(_02058_));
 sky130_fd_sc_hd__nand3_4 _25133_ (.A(_02058_),
    .B(_02028_),
    .C(_02056_),
    .Y(_02060_));
 sky130_fd_sc_hd__o22a_1 _25134_ (.A1(_01809_),
    .A2(_02027_),
    .B1(_02055_),
    .B2(_02057_),
    .X(_02061_));
 sky130_fd_sc_hd__o22ai_4 _25135_ (.A1(_01809_),
    .A2(_02027_),
    .B1(_02055_),
    .B2(_02057_),
    .Y(_02062_));
 sky130_fd_sc_hd__o21ai_2 _25136_ (.A1(_02025_),
    .A2(_02061_),
    .B1(_02060_),
    .Y(_02063_));
 sky130_fd_sc_hd__a2bb2oi_1 _25137_ (.A1_N(_01903_),
    .A2_N(_02023_),
    .B1(_02060_),
    .B2(_02062_),
    .Y(_02064_));
 sky130_fd_sc_hd__a2bb2o_2 _25138_ (.A1_N(_01903_),
    .A2_N(_02023_),
    .B1(_02060_),
    .B2(_02062_),
    .X(_02065_));
 sky130_fd_sc_hd__o211a_1 _25139_ (.A1(_01907_),
    .A2(_02024_),
    .B1(_02060_),
    .C1(_02062_),
    .X(_02066_));
 sky130_fd_sc_hd__o211ai_4 _25140_ (.A1(_01907_),
    .A2(_02024_),
    .B1(_02060_),
    .C1(_02062_),
    .Y(_02067_));
 sky130_fd_sc_hd__o22ai_4 _25141_ (.A1(_01916_),
    .A2(_02021_),
    .B1(_02064_),
    .B2(_02066_),
    .Y(_02068_));
 sky130_fd_sc_hd__o21ai_1 _25142_ (.A1(_01914_),
    .A2(_01920_),
    .B1(_02065_),
    .Y(_02069_));
 sky130_fd_sc_hd__and3_1 _25143_ (.A(_02022_),
    .B(_02065_),
    .C(_02067_),
    .X(_02071_));
 sky130_fd_sc_hd__o211ai_4 _25144_ (.A1(_01914_),
    .A2(_01920_),
    .B1(_02065_),
    .C1(_02067_),
    .Y(_02072_));
 sky130_fd_sc_hd__a31oi_4 _25145_ (.A1(_02022_),
    .A2(_02065_),
    .A3(_02067_),
    .B1(_02020_),
    .Y(_02073_));
 sky130_fd_sc_hd__o211a_2 _25146_ (.A1(_02066_),
    .A2(_02069_),
    .B1(_02068_),
    .C1(_02019_),
    .X(_02074_));
 sky130_fd_sc_hd__nand2_2 _25147_ (.A(_02073_),
    .B(_02068_),
    .Y(_02075_));
 sky130_fd_sc_hd__a2bb2oi_2 _25148_ (.A1_N(_02014_),
    .A2_N(_02018_),
    .B1(_02068_),
    .B2(_02072_),
    .Y(_02076_));
 sky130_fd_sc_hd__a2bb2o_1 _25149_ (.A1_N(_02014_),
    .A2_N(_02018_),
    .B1(_02068_),
    .B2(_02072_),
    .X(_02077_));
 sky130_fd_sc_hd__a221oi_4 _25150_ (.A1(_01821_),
    .A2(_01825_),
    .B1(_02073_),
    .B2(_02068_),
    .C1(_02076_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand3_2 _25151_ (.A(_02077_),
    .B(_01980_),
    .C(_02075_),
    .Y(_02079_));
 sky130_fd_sc_hd__a2bb2oi_2 _25152_ (.A1_N(_01820_),
    .A2_N(_01979_),
    .B1(_02075_),
    .B2(_02077_),
    .Y(_02080_));
 sky130_fd_sc_hd__o22ai_4 _25153_ (.A1(_01820_),
    .A2(_01979_),
    .B1(_02074_),
    .B2(_02076_),
    .Y(_02082_));
 sky130_fd_sc_hd__o22ai_4 _25154_ (.A1(_01927_),
    .A2(_01930_),
    .B1(_02078_),
    .B2(_02080_),
    .Y(_02083_));
 sky130_fd_sc_hd__o311a_1 _25155_ (.A1(_01879_),
    .A2(_01880_),
    .A3(_01925_),
    .B1(_01929_),
    .C1(_02082_),
    .X(_02084_));
 sky130_fd_sc_hd__nand3b_2 _25156_ (.A_N(_01932_),
    .B(_02079_),
    .C(_02082_),
    .Y(_02085_));
 sky130_fd_sc_hd__a22o_1 _25157_ (.A1(_01926_),
    .A2(_01931_),
    .B1(_02079_),
    .B2(_02082_),
    .X(_02086_));
 sky130_fd_sc_hd__o211ai_1 _25158_ (.A1(_01927_),
    .A2(_01930_),
    .B1(_02079_),
    .C1(_02082_),
    .Y(_02087_));
 sky130_fd_sc_hd__a32oi_4 _25159_ (.A1(_01770_),
    .A2(_01771_),
    .A3(_01773_),
    .B1(_01777_),
    .B2(_01829_),
    .Y(_02088_));
 sky130_fd_sc_hd__a2bb2oi_2 _25160_ (.A1_N(_01756_),
    .A2_N(_01751_),
    .B1(_12099_),
    .B2(_01757_),
    .Y(_02089_));
 sky130_fd_sc_hd__o2bb2ai_1 _25161_ (.A1_N(_12099_),
    .A2_N(_01757_),
    .B1(_01756_),
    .B2(_01751_),
    .Y(_02090_));
 sky130_fd_sc_hd__o21a_1 _25162_ (.A1(net140),
    .A2(net136),
    .B1(_01748_),
    .X(_02091_));
 sky130_fd_sc_hd__a32o_1 _25163_ (.A1(_01745_),
    .A2(_01733_),
    .A3(_01744_),
    .B1(_10544_),
    .B2(net139),
    .X(_02093_));
 sky130_fd_sc_hd__a32oi_4 _25164_ (.A1(_01734_),
    .A2(_01746_),
    .A3(_01747_),
    .B1(_01748_),
    .B2(_10546_),
    .Y(_02094_));
 sky130_fd_sc_hd__nor2_1 _25165_ (.A(net144),
    .B(_01740_),
    .Y(_02095_));
 sky130_fd_sc_hd__o22ai_1 _25166_ (.A1(_01735_),
    .A2(_01738_),
    .B1(net144),
    .B2(_01740_),
    .Y(_02096_));
 sky130_fd_sc_hd__or3_2 _25167_ (.A(net57),
    .B(_04266_),
    .C(_04113_),
    .X(_02097_));
 sky130_fd_sc_hd__nand3_4 _25168_ (.A(net209),
    .B(_05074_),
    .C(_08657_),
    .Y(_02098_));
 sky130_fd_sc_hd__o21ai_1 _25169_ (.A1(_04113_),
    .A2(_08660_),
    .B1(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__o311a_1 _25170_ (.A1(_04113_),
    .A2(net57),
    .A3(_04266_),
    .B1(_02098_),
    .C1(net149),
    .X(_02100_));
 sky130_fd_sc_hd__nand3_2 _25171_ (.A(net149),
    .B(_02097_),
    .C(_02098_),
    .Y(_02101_));
 sky130_fd_sc_hd__a21oi_4 _25172_ (.A1(_02097_),
    .A2(_02098_),
    .B1(net149),
    .Y(_02102_));
 sky130_fd_sc_hd__nand2_1 _25173_ (.A(_02099_),
    .B(net157),
    .Y(_02104_));
 sky130_fd_sc_hd__o22a_4 _25174_ (.A1(net237),
    .A2(_09297_),
    .B1(net157),
    .B2(_02099_),
    .X(_02105_));
 sky130_fd_sc_hd__a21oi_2 _25175_ (.A1(_02101_),
    .A2(_02104_),
    .B1(net144),
    .Y(_02106_));
 sky130_fd_sc_hd__o21ai_1 _25176_ (.A1(_02100_),
    .A2(_02102_),
    .B1(net145),
    .Y(_02107_));
 sky130_fd_sc_hd__o21ai_2 _25177_ (.A1(_01740_),
    .A2(_01743_),
    .B1(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__nor3_2 _25178_ (.A(_02096_),
    .B(_02105_),
    .C(_02106_),
    .Y(_02109_));
 sky130_fd_sc_hd__o22a_1 _25179_ (.A1(_01739_),
    .A2(_02095_),
    .B1(_02105_),
    .B2(_02106_),
    .X(_02110_));
 sky130_fd_sc_hd__o22ai_4 _25180_ (.A1(_01739_),
    .A2(_02095_),
    .B1(_02105_),
    .B2(_02106_),
    .Y(_02111_));
 sky130_fd_sc_hd__o22ai_2 _25181_ (.A1(net140),
    .A2(net136),
    .B1(_02109_),
    .B2(_02110_),
    .Y(_02112_));
 sky130_fd_sc_hd__o211ai_2 _25182_ (.A1(_02105_),
    .A2(_02108_),
    .B1(_02111_),
    .C1(_10545_),
    .Y(_02113_));
 sky130_fd_sc_hd__o221ai_4 _25183_ (.A1(net140),
    .A2(net136),
    .B1(_02105_),
    .B2(_02108_),
    .C1(_02111_),
    .Y(_02115_));
 sky130_fd_sc_hd__o21ai_1 _25184_ (.A1(_02109_),
    .A2(_02110_),
    .B1(net133),
    .Y(_02116_));
 sky130_fd_sc_hd__a22oi_1 _25185_ (.A1(_01750_),
    .A2(_02093_),
    .B1(_02112_),
    .B2(_02113_),
    .Y(_02117_));
 sky130_fd_sc_hd__o211ai_4 _25186_ (.A1(_01749_),
    .A2(_02091_),
    .B1(_02115_),
    .C1(_02116_),
    .Y(_02118_));
 sky130_fd_sc_hd__nand3_4 _25187_ (.A(_02112_),
    .B(_02113_),
    .C(_02094_),
    .Y(_02119_));
 sky130_fd_sc_hd__inv_2 _25188_ (.A(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__o2bb2ai_2 _25189_ (.A1_N(_02118_),
    .A2_N(_02119_),
    .B1(net141),
    .B2(_11742_),
    .Y(_02121_));
 sky130_fd_sc_hd__o2111ai_4 _25190_ (.A1(_11737_),
    .A2(_11740_),
    .B1(_02119_),
    .C1(net143),
    .D1(_02118_),
    .Y(_02122_));
 sky130_fd_sc_hd__a21o_1 _25191_ (.A1(_02118_),
    .A2(_02119_),
    .B1(_12099_),
    .X(_02123_));
 sky130_fd_sc_hd__o21ai_2 _25192_ (.A1(net141),
    .A2(_11742_),
    .B1(_02118_),
    .Y(_02124_));
 sky130_fd_sc_hd__nand3_4 _25193_ (.A(_02089_),
    .B(_02121_),
    .C(_02122_),
    .Y(_02126_));
 sky130_fd_sc_hd__inv_2 _25194_ (.A(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__a21oi_1 _25195_ (.A1(_02121_),
    .A2(_02122_),
    .B1(_02089_),
    .Y(_02128_));
 sky130_fd_sc_hd__o211ai_4 _25196_ (.A1(_02124_),
    .A2(_02120_),
    .B1(_02090_),
    .C1(_02123_),
    .Y(_02129_));
 sky130_fd_sc_hd__a22o_1 _25197_ (.A1(_00364_),
    .A2(_00367_),
    .B1(_02126_),
    .B2(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__o2111ai_4 _25198_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_02126_),
    .D1(_02129_),
    .Y(_02131_));
 sky130_fd_sc_hd__o211ai_2 _25199_ (.A1(net130),
    .A2(_00366_),
    .B1(_02126_),
    .C1(_02129_),
    .Y(_02132_));
 sky130_fd_sc_hd__a21o_1 _25200_ (.A1(_02126_),
    .A2(_02129_),
    .B1(_00737_),
    .X(_02133_));
 sky130_fd_sc_hd__o21ai_2 _25201_ (.A1(_00737_),
    .A2(_01762_),
    .B1(_01767_),
    .Y(_02134_));
 sky130_fd_sc_hd__o2111ai_4 _25202_ (.A1(_00737_),
    .A2(_01762_),
    .B1(_01767_),
    .C1(_02132_),
    .D1(_02133_),
    .Y(_02135_));
 sky130_fd_sc_hd__and3_1 _25203_ (.A(_02130_),
    .B(_02134_),
    .C(_02131_),
    .X(_02137_));
 sky130_fd_sc_hd__nand3_4 _25204_ (.A(_02130_),
    .B(_02134_),
    .C(_02131_),
    .Y(_02138_));
 sky130_fd_sc_hd__o22a_1 _25205_ (.A1(_04245_),
    .A2(_05465_),
    .B1(_07772_),
    .B2(_05463_),
    .X(_02139_));
 sky130_fd_sc_hd__a32o_1 _25206_ (.A1(_07771_),
    .A2(_05462_),
    .A3(net166),
    .B1(_05464_),
    .B2(net22),
    .X(_02140_));
 sky130_fd_sc_hd__a32oi_4 _25207_ (.A1(net164),
    .A2(_08208_),
    .A3(_05225_),
    .B1(_05228_),
    .B2(net24),
    .Y(_02141_));
 sky130_fd_sc_hd__a32o_1 _25208_ (.A1(net164),
    .A2(_08208_),
    .A3(_05225_),
    .B1(_05228_),
    .B2(net24),
    .X(_02142_));
 sky130_fd_sc_hd__a21oi_1 _25209_ (.A1(_08665_),
    .A2(_08668_),
    .B1(_04986_),
    .Y(_02143_));
 sky130_fd_sc_hd__o21ai_1 _25210_ (.A1(_08664_),
    .A2(_08666_),
    .B1(net242),
    .Y(_02144_));
 sky130_fd_sc_hd__and3_1 _25211_ (.A(_04124_),
    .B(net25),
    .C(net43),
    .X(_02145_));
 sky130_fd_sc_hd__or3_4 _25212_ (.A(net45),
    .B(net319),
    .C(_04102_),
    .X(_02146_));
 sky130_fd_sc_hd__a21oi_1 _25213_ (.A1(_02144_),
    .A2(_02146_),
    .B1(_02141_),
    .Y(_02148_));
 sky130_fd_sc_hd__o21ai_1 _25214_ (.A1(_02143_),
    .A2(_02145_),
    .B1(_02142_),
    .Y(_02149_));
 sky130_fd_sc_hd__o311a_1 _25215_ (.A1(_04102_),
    .A2(net45),
    .A3(net319),
    .B1(_02141_),
    .C1(_02144_),
    .X(_02150_));
 sky130_fd_sc_hd__o211ai_1 _25216_ (.A1(net319),
    .A2(_04989_),
    .B1(_02141_),
    .C1(_02144_),
    .Y(_02151_));
 sky130_fd_sc_hd__o21ai_1 _25217_ (.A1(_02143_),
    .A2(_02145_),
    .B1(_02141_),
    .Y(_02152_));
 sky130_fd_sc_hd__o221ai_2 _25218_ (.A1(net319),
    .A2(_04989_),
    .B1(_04986_),
    .B2(_08669_),
    .C1(_02142_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand3_1 _25219_ (.A(_02140_),
    .B(_02149_),
    .C(_02151_),
    .Y(_02154_));
 sky130_fd_sc_hd__nand3_2 _25220_ (.A(_02152_),
    .B(_02153_),
    .C(_02139_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _25221_ (.A(_02154_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__o22a_2 _25222_ (.A1(net319),
    .A2(_04898_),
    .B1(_08665_),
    .B2(_04896_),
    .X(_02157_));
 sky130_fd_sc_hd__o2111a_4 _25223_ (.A1(_04481_),
    .A2(_08665_),
    .B1(_01493_),
    .C1(_01497_),
    .D1(_02157_),
    .X(_02159_));
 sky130_fd_sc_hd__nand2_4 _25224_ (.A(_01801_),
    .B(_02157_),
    .Y(_02160_));
 sky130_fd_sc_hd__a31o_1 _25225_ (.A1(net25),
    .A2(_04895_),
    .A3(_08207_),
    .B1(_02159_),
    .X(_02161_));
 sky130_fd_sc_hd__nand2_4 _25226_ (.A(_02156_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__o2111ai_4 _25227_ (.A1(_04896_),
    .A2(_08668_),
    .B1(_02154_),
    .C1(_02155_),
    .D1(_02160_),
    .Y(_02163_));
 sky130_fd_sc_hd__a21o_1 _25228_ (.A1(_02162_),
    .A2(_02163_),
    .B1(_01332_),
    .X(_02164_));
 sky130_fd_sc_hd__and3_1 _25229_ (.A(_01332_),
    .B(_02162_),
    .C(_02163_),
    .X(_02165_));
 sky130_fd_sc_hd__o211ai_2 _25230_ (.A1(_00796_),
    .A2(_01324_),
    .B1(_02162_),
    .C1(_02163_),
    .Y(_02166_));
 sky130_fd_sc_hd__and3_1 _25231_ (.A(_02164_),
    .B(_02166_),
    .C(net130),
    .X(_02167_));
 sky130_fd_sc_hd__o2111ai_1 _25232_ (.A1(_13066_),
    .A2(_00357_),
    .B1(_02166_),
    .C1(_11740_),
    .D1(_02164_),
    .Y(_02168_));
 sky130_fd_sc_hd__o2bb2ai_1 _25233_ (.A1_N(_02164_),
    .A2_N(_02166_),
    .B1(_11741_),
    .B2(_00360_),
    .Y(_02170_));
 sky130_fd_sc_hd__nand2_1 _25234_ (.A(_02168_),
    .B(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__and4_2 _25235_ (.A(_01332_),
    .B(_01813_),
    .C(_01815_),
    .D(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__o311a_2 _25236_ (.A1(_01331_),
    .A2(_01812_),
    .A3(_01814_),
    .B1(_02168_),
    .C1(_02170_),
    .X(_02173_));
 sky130_fd_sc_hd__o31a_1 _25237_ (.A1(_01331_),
    .A2(_01812_),
    .A3(_01814_),
    .B1(_02171_),
    .X(_02174_));
 sky130_fd_sc_hd__nor2_1 _25238_ (.A(_01816_),
    .B(_02171_),
    .Y(_02175_));
 sky130_fd_sc_hd__o211ai_4 _25239_ (.A1(_02172_),
    .A2(_02173_),
    .B1(_02135_),
    .C1(_02138_),
    .Y(_02176_));
 sky130_fd_sc_hd__o2bb2ai_1 _25240_ (.A1_N(_02135_),
    .A2_N(_02138_),
    .B1(_02174_),
    .B2(_02175_),
    .Y(_02177_));
 sky130_fd_sc_hd__o211ai_2 _25241_ (.A1(_02174_),
    .A2(_02175_),
    .B1(_02135_),
    .C1(_02138_),
    .Y(_02178_));
 sky130_fd_sc_hd__o2bb2ai_2 _25242_ (.A1_N(_02135_),
    .A2_N(_02138_),
    .B1(_02172_),
    .B2(_02173_),
    .Y(_02179_));
 sky130_fd_sc_hd__and3_1 _25243_ (.A(_02177_),
    .B(_02088_),
    .C(_02176_),
    .X(_02181_));
 sky130_fd_sc_hd__nand3_1 _25244_ (.A(_02177_),
    .B(_02088_),
    .C(_02176_),
    .Y(_02182_));
 sky130_fd_sc_hd__o2111a_1 _25245_ (.A1(_01829_),
    .A2(_01774_),
    .B1(_01777_),
    .C1(_02178_),
    .D1(_02179_),
    .X(_02183_));
 sky130_fd_sc_hd__o2111ai_4 _25246_ (.A1(_01829_),
    .A2(_01774_),
    .B1(_01777_),
    .C1(_02178_),
    .D1(_02179_),
    .Y(_02184_));
 sky130_fd_sc_hd__nand3_1 _25247_ (.A(_02083_),
    .B(_02085_),
    .C(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand4_2 _25248_ (.A(_02083_),
    .B(_02085_),
    .C(_02182_),
    .D(_02184_),
    .Y(_02186_));
 sky130_fd_sc_hd__a22o_1 _25249_ (.A1(_02083_),
    .A2(_02085_),
    .B1(_02182_),
    .B2(_02184_),
    .X(_02187_));
 sky130_fd_sc_hd__o211a_1 _25250_ (.A1(_02181_),
    .A2(_02185_),
    .B1(_02187_),
    .C1(_01978_),
    .X(_02188_));
 sky130_fd_sc_hd__o211ai_2 _25251_ (.A1(_02181_),
    .A2(_02185_),
    .B1(_02187_),
    .C1(_01978_),
    .Y(_02189_));
 sky130_fd_sc_hd__a21oi_2 _25252_ (.A1(_02186_),
    .A2(_02187_),
    .B1(_01978_),
    .Y(_02190_));
 sky130_fd_sc_hd__a21o_1 _25253_ (.A1(_02186_),
    .A2(_02187_),
    .B1(_01978_),
    .X(_02192_));
 sky130_fd_sc_hd__nand3_2 _25254_ (.A(_02192_),
    .B(_01976_),
    .C(_02189_),
    .Y(_02193_));
 sky130_fd_sc_hd__o22ai_4 _25255_ (.A1(_01936_),
    .A2(_01975_),
    .B1(_02188_),
    .B2(_02190_),
    .Y(_02194_));
 sky130_fd_sc_hd__and3_1 _25256_ (.A(_01974_),
    .B(_02193_),
    .C(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__nand3_1 _25257_ (.A(_01974_),
    .B(_02193_),
    .C(_02194_),
    .Y(_02196_));
 sky130_fd_sc_hd__a21oi_2 _25258_ (.A1(_02193_),
    .A2(_02194_),
    .B1(_01974_),
    .Y(_02197_));
 sky130_fd_sc_hd__a31o_1 _25259_ (.A1(_01974_),
    .A2(_02193_),
    .A3(_02194_),
    .B1(_01877_),
    .X(_02198_));
 sky130_fd_sc_hd__o21ai_1 _25260_ (.A1(_01878_),
    .A2(_02197_),
    .B1(_02196_),
    .Y(_02199_));
 sky130_fd_sc_hd__nand3b_1 _25261_ (.A_N(_02197_),
    .B(_01877_),
    .C(_02196_),
    .Y(_02200_));
 sky130_fd_sc_hd__o22ai_1 _25262_ (.A1(_01874_),
    .A2(_01876_),
    .B1(_02195_),
    .B2(_02197_),
    .Y(_02201_));
 sky130_fd_sc_hd__o21ai_1 _25263_ (.A1(_02195_),
    .A2(_02197_),
    .B1(_01878_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand3_1 _25264_ (.A(_02203_),
    .B(_01972_),
    .C(_02200_),
    .Y(_02204_));
 sky130_fd_sc_hd__o211a_1 _25265_ (.A1(_02198_),
    .A2(_02197_),
    .B1(_01973_),
    .C1(_02201_),
    .X(_02205_));
 sky130_fd_sc_hd__o211ai_1 _25266_ (.A1(_02198_),
    .A2(_02197_),
    .B1(_01973_),
    .C1(_02201_),
    .Y(_02206_));
 sky130_fd_sc_hd__nand2_1 _25267_ (.A(_02204_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__o21a_1 _25268_ (.A1(_01725_),
    .A2(_01968_),
    .B1(_01969_),
    .X(_02208_));
 sky130_fd_sc_hd__xor2_1 _25269_ (.A(_02207_),
    .B(_02208_),
    .X(net111));
 sky130_fd_sc_hd__a32oi_2 _25270_ (.A1(_02088_),
    .A2(_02176_),
    .A3(_02177_),
    .B1(_02085_),
    .B2(_02083_),
    .Y(_02209_));
 sky130_fd_sc_hd__a31oi_1 _25271_ (.A1(_02086_),
    .A2(_02087_),
    .A3(_02182_),
    .B1(_02183_),
    .Y(_02210_));
 sky130_fd_sc_hd__o21ai_1 _25272_ (.A1(_02174_),
    .A2(_02175_),
    .B1(_02138_),
    .Y(_02211_));
 sky130_fd_sc_hd__o21a_1 _25273_ (.A1(_02172_),
    .A2(_02173_),
    .B1(_02135_),
    .X(_02213_));
 sky130_fd_sc_hd__nand2_1 _25274_ (.A(_02135_),
    .B(_02211_),
    .Y(_02214_));
 sky130_fd_sc_hd__o21a_1 _25275_ (.A1(net130),
    .A2(_00366_),
    .B1(_02129_),
    .X(_02215_));
 sky130_fd_sc_hd__a31o_1 _25276_ (.A1(_00364_),
    .A2(_00367_),
    .A3(_02126_),
    .B1(_02128_),
    .X(_02216_));
 sky130_fd_sc_hd__a21oi_4 _25277_ (.A1(net144),
    .A2(_02101_),
    .B1(_02102_),
    .Y(_02217_));
 sky130_fd_sc_hd__a32o_1 _25278_ (.A1(_08876_),
    .A2(_02099_),
    .A3(net319),
    .B1(_02101_),
    .B2(net144),
    .X(_02218_));
 sky130_fd_sc_hd__or3_2 _25279_ (.A(net57),
    .B(_04266_),
    .C(_04135_),
    .X(_02219_));
 sky130_fd_sc_hd__nand3_4 _25280_ (.A(_05290_),
    .B(_05292_),
    .C(_08657_),
    .Y(_02220_));
 sky130_fd_sc_hd__a21oi_4 _25281_ (.A1(_02219_),
    .A2(_02220_),
    .B1(net149),
    .Y(_02221_));
 sky130_fd_sc_hd__a21o_1 _25282_ (.A1(_02219_),
    .A2(_02220_),
    .B1(net149),
    .X(_02222_));
 sky130_fd_sc_hd__o311a_4 _25283_ (.A1(_04135_),
    .A2(net57),
    .A3(_04266_),
    .B1(_02220_),
    .C1(net149),
    .X(_02224_));
 sky130_fd_sc_hd__o211ai_4 _25284_ (.A1(_04135_),
    .A2(_08660_),
    .B1(net149),
    .C1(_02220_),
    .Y(_02225_));
 sky130_fd_sc_hd__o21ai_4 _25285_ (.A1(_02221_),
    .A2(_02224_),
    .B1(net145),
    .Y(_02226_));
 sky130_fd_sc_hd__a31o_1 _25286_ (.A1(net149),
    .A2(_02219_),
    .A3(_02220_),
    .B1(net145),
    .X(_02227_));
 sky130_fd_sc_hd__o22ai_4 _25287_ (.A1(net237),
    .A2(_09297_),
    .B1(_02221_),
    .B2(_02224_),
    .Y(_02228_));
 sky130_fd_sc_hd__nand3_4 _25288_ (.A(_02222_),
    .B(_02225_),
    .C(net145),
    .Y(_02229_));
 sky130_fd_sc_hd__o21ai_1 _25289_ (.A1(net145),
    .A2(_02224_),
    .B1(_02226_),
    .Y(_02230_));
 sky130_fd_sc_hd__a21oi_2 _25290_ (.A1(_02228_),
    .A2(_02229_),
    .B1(_02217_),
    .Y(_02231_));
 sky130_fd_sc_hd__o221ai_4 _25291_ (.A1(_02102_),
    .A2(_02105_),
    .B1(_02224_),
    .B2(net145),
    .C1(_02226_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21oi_2 _25292_ (.A1(_02226_),
    .A2(_02227_),
    .B1(_02218_),
    .Y(_02233_));
 sky130_fd_sc_hd__o2111ai_2 _25293_ (.A1(net145),
    .A2(_02100_),
    .B1(_02104_),
    .C1(_02228_),
    .D1(_02229_),
    .Y(_02235_));
 sky130_fd_sc_hd__o22ai_1 _25294_ (.A1(net140),
    .A2(net136),
    .B1(_02231_),
    .B2(_02233_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand4_1 _25295_ (.A(net139),
    .B(_10544_),
    .C(_02232_),
    .D(_02235_),
    .Y(_02237_));
 sky130_fd_sc_hd__a211o_1 _25296_ (.A1(_02228_),
    .A2(_02229_),
    .B1(_02217_),
    .C1(_10546_),
    .X(_02238_));
 sky130_fd_sc_hd__o2111ai_4 _25297_ (.A1(net140),
    .A2(net136),
    .B1(_02217_),
    .C1(_02228_),
    .D1(_02229_),
    .Y(_02239_));
 sky130_fd_sc_hd__a31oi_2 _25298_ (.A1(_02218_),
    .A2(_02226_),
    .A3(_02227_),
    .B1(_10545_),
    .Y(_02240_));
 sky130_fd_sc_hd__a311oi_4 _25299_ (.A1(_02228_),
    .A2(_02229_),
    .A3(_02217_),
    .B1(net136),
    .C1(net140),
    .Y(_02241_));
 sky130_fd_sc_hd__a31o_1 _25300_ (.A1(_02228_),
    .A2(_02229_),
    .A3(_02217_),
    .B1(_10546_),
    .X(_02242_));
 sky130_fd_sc_hd__a21oi_1 _25301_ (.A1(_02235_),
    .A2(_10545_),
    .B1(_02231_),
    .Y(_02243_));
 sky130_fd_sc_hd__o211ai_4 _25302_ (.A1(_02217_),
    .A2(_02230_),
    .B1(_02239_),
    .C1(_02242_),
    .Y(_02244_));
 sky130_fd_sc_hd__o2bb2ai_1 _25303_ (.A1_N(_10545_),
    .A2_N(_02111_),
    .B1(_02108_),
    .B2(_02105_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21oi_4 _25304_ (.A1(_02111_),
    .A2(_10545_),
    .B1(_02109_),
    .Y(_02247_));
 sky130_fd_sc_hd__o211ai_4 _25305_ (.A1(_10546_),
    .A2(_02232_),
    .B1(_02244_),
    .C1(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__a21oi_2 _25306_ (.A1(_02238_),
    .A2(_02244_),
    .B1(_02247_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand3_2 _25307_ (.A(_02236_),
    .B(_02237_),
    .C(_02246_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21oi_1 _25308_ (.A1(_02248_),
    .A2(_02250_),
    .B1(_12099_),
    .Y(_02251_));
 sky130_fd_sc_hd__a21o_1 _25309_ (.A1(_02248_),
    .A2(_02250_),
    .B1(_12099_),
    .X(_02252_));
 sky130_fd_sc_hd__a31oi_4 _25310_ (.A1(_02238_),
    .A2(_02244_),
    .A3(_02247_),
    .B1(net132),
    .Y(_02253_));
 sky130_fd_sc_hd__o311a_1 _25311_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_02248_),
    .C1(_02250_),
    .X(_02254_));
 sky130_fd_sc_hd__nand2_1 _25312_ (.A(_02253_),
    .B(_02250_),
    .Y(_02255_));
 sky130_fd_sc_hd__o21ai_1 _25313_ (.A1(net132),
    .A2(_02117_),
    .B1(_02119_),
    .Y(_02257_));
 sky130_fd_sc_hd__a221oi_2 _25314_ (.A1(_02253_),
    .A2(_02250_),
    .B1(_02124_),
    .B2(_02119_),
    .C1(_02251_),
    .Y(_02258_));
 sky130_fd_sc_hd__nand3_1 _25315_ (.A(_02252_),
    .B(_02255_),
    .C(_02257_),
    .Y(_02259_));
 sky130_fd_sc_hd__a21oi_1 _25316_ (.A1(_02252_),
    .A2(_02255_),
    .B1(_02257_),
    .Y(_02260_));
 sky130_fd_sc_hd__o21bai_2 _25317_ (.A1(_02251_),
    .A2(_02254_),
    .B1_N(_02257_),
    .Y(_02261_));
 sky130_fd_sc_hd__o2111a_2 _25318_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_02259_),
    .D1(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__o2111ai_2 _25319_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_02259_),
    .D1(_02261_),
    .Y(_02263_));
 sky130_fd_sc_hd__o22a_1 _25320_ (.A1(net130),
    .A2(_00366_),
    .B1(_02258_),
    .B2(_02260_),
    .X(_02264_));
 sky130_fd_sc_hd__o22ai_2 _25321_ (.A1(net130),
    .A2(_00366_),
    .B1(_02258_),
    .B2(_02260_),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2_2 _25322_ (.A(_02216_),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__nand3_2 _25323_ (.A(_02216_),
    .B(_02263_),
    .C(_02265_),
    .Y(_02268_));
 sky130_fd_sc_hd__a2bb2oi_1 _25324_ (.A1_N(_02127_),
    .A2_N(_02215_),
    .B1(_02263_),
    .B2(_02265_),
    .Y(_02269_));
 sky130_fd_sc_hd__o22ai_4 _25325_ (.A1(_02127_),
    .A2(_02215_),
    .B1(_02262_),
    .B2(_02264_),
    .Y(_02270_));
 sky130_fd_sc_hd__o32a_1 _25326_ (.A1(_05463_),
    .A2(_08203_),
    .A3(_08207_),
    .B1(_05465_),
    .B2(_04256_),
    .X(_02271_));
 sky130_fd_sc_hd__a32o_1 _25327_ (.A1(net164),
    .A2(_08208_),
    .A3(_05462_),
    .B1(_05464_),
    .B2(net24),
    .X(_02272_));
 sky130_fd_sc_hd__o211ai_2 _25328_ (.A1(net170),
    .A2(net268),
    .B1(net319),
    .C1(net242),
    .Y(_02273_));
 sky130_fd_sc_hd__a31oi_4 _25329_ (.A1(net319),
    .A2(_08208_),
    .A3(net242),
    .B1(_02145_),
    .Y(_02274_));
 sky130_fd_sc_hd__a21oi_1 _25330_ (.A1(net153),
    .A2(_08668_),
    .B1(_05226_),
    .Y(_02275_));
 sky130_fd_sc_hd__o21ai_2 _25331_ (.A1(_08664_),
    .A2(_08666_),
    .B1(_05225_),
    .Y(_02276_));
 sky130_fd_sc_hd__nor2_1 _25332_ (.A(net319),
    .B(_05229_),
    .Y(_02277_));
 sky130_fd_sc_hd__or3_4 _25333_ (.A(net46),
    .B(net319),
    .C(_04124_),
    .X(_02279_));
 sky130_fd_sc_hd__a22oi_2 _25334_ (.A1(_02146_),
    .A2(_02273_),
    .B1(_02276_),
    .B2(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__o21bai_4 _25335_ (.A1(_02275_),
    .A2(_02277_),
    .B1_N(_02274_),
    .Y(_02281_));
 sky130_fd_sc_hd__o311a_1 _25336_ (.A1(_04124_),
    .A2(net46),
    .A3(net319),
    .B1(_02274_),
    .C1(_02276_),
    .X(_02282_));
 sky130_fd_sc_hd__o2111ai_4 _25337_ (.A1(_04986_),
    .A2(net153),
    .B1(_02146_),
    .C1(_02276_),
    .D1(_02279_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand3_2 _25338_ (.A(_02272_),
    .B(_02281_),
    .C(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__o21ai_1 _25339_ (.A1(_02280_),
    .A2(_02282_),
    .B1(_02271_),
    .Y(_02285_));
 sky130_fd_sc_hd__o21ai_1 _25340_ (.A1(_02280_),
    .A2(_02282_),
    .B1(_02272_),
    .Y(_02286_));
 sky130_fd_sc_hd__nand3_1 _25341_ (.A(_02281_),
    .B(_02283_),
    .C(_02271_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand3_4 _25342_ (.A(_02160_),
    .B(_02284_),
    .C(_02285_),
    .Y(_02288_));
 sky130_fd_sc_hd__inv_2 _25343_ (.A(_02288_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand4_2 _25344_ (.A(_02286_),
    .B(_02287_),
    .C(_01801_),
    .D(_02157_),
    .Y(_02291_));
 sky130_fd_sc_hd__a21oi_2 _25345_ (.A1(_02288_),
    .A2(_02291_),
    .B1(_01332_),
    .Y(_02292_));
 sky130_fd_sc_hd__and3_2 _25346_ (.A(_01332_),
    .B(_02288_),
    .C(_02291_),
    .X(_02293_));
 sky130_fd_sc_hd__a2bb2o_2 _25347_ (.A1_N(_02292_),
    .A2_N(_02293_),
    .B1(_11740_),
    .B2(_00361_),
    .X(_02294_));
 sky130_fd_sc_hd__a2111oi_4 _25348_ (.A1(_13065_),
    .A2(_00358_),
    .B1(_11741_),
    .C1(_02292_),
    .D1(_02293_),
    .Y(_02295_));
 sky130_fd_sc_hd__a2111o_2 _25349_ (.A1(_13065_),
    .A2(_00358_),
    .B1(_11741_),
    .C1(_02292_),
    .D1(_02293_),
    .X(_02296_));
 sky130_fd_sc_hd__nand2_1 _25350_ (.A(_02294_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__and3_1 _25351_ (.A(_02296_),
    .B(_02165_),
    .C(_02294_),
    .X(_02298_));
 sky130_fd_sc_hd__a21oi_2 _25352_ (.A1(_02294_),
    .A2(_02296_),
    .B1(_02165_),
    .Y(_02299_));
 sky130_fd_sc_hd__and4_1 _25353_ (.A(_01332_),
    .B(_02162_),
    .C(_02163_),
    .D(_02297_),
    .X(_02301_));
 sky130_fd_sc_hd__a21o_1 _25354_ (.A1(_02294_),
    .A2(_02296_),
    .B1(_02166_),
    .X(_02302_));
 sky130_fd_sc_hd__and3_1 _25355_ (.A(_02166_),
    .B(_02294_),
    .C(_02296_),
    .X(_02303_));
 sky130_fd_sc_hd__a31o_1 _25356_ (.A1(_01332_),
    .A2(_02162_),
    .A3(_02163_),
    .B1(_02297_),
    .X(_02304_));
 sky130_fd_sc_hd__nor2_1 _25357_ (.A(_02298_),
    .B(_02299_),
    .Y(_02305_));
 sky130_fd_sc_hd__o221ai_4 _25358_ (.A1(_02298_),
    .A2(_02299_),
    .B1(_02262_),
    .B2(_02266_),
    .C1(_02270_),
    .Y(_02306_));
 sky130_fd_sc_hd__o2bb2ai_1 _25359_ (.A1_N(_02268_),
    .A2_N(_02270_),
    .B1(_02301_),
    .B2(_02303_),
    .Y(_02307_));
 sky130_fd_sc_hd__o2bb2ai_1 _25360_ (.A1_N(_02268_),
    .A2_N(_02270_),
    .B1(_02298_),
    .B2(_02299_),
    .Y(_02308_));
 sky130_fd_sc_hd__o221ai_2 _25361_ (.A1(_02301_),
    .A2(_02303_),
    .B1(_02262_),
    .B2(_02266_),
    .C1(_02270_),
    .Y(_02309_));
 sky130_fd_sc_hd__nand3_2 _25362_ (.A(_02214_),
    .B(_02306_),
    .C(_02307_),
    .Y(_02310_));
 sky130_fd_sc_hd__a22oi_2 _25363_ (.A1(_02138_),
    .A2(_02176_),
    .B1(_02306_),
    .B2(_02307_),
    .Y(_02312_));
 sky130_fd_sc_hd__o211ai_2 _25364_ (.A1(_02137_),
    .A2(_02213_),
    .B1(_02308_),
    .C1(_02309_),
    .Y(_02313_));
 sky130_fd_sc_hd__a31o_1 _25365_ (.A1(_02022_),
    .A2(_02065_),
    .A3(_02067_),
    .B1(_02074_),
    .X(_02314_));
 sky130_fd_sc_hd__a41o_1 _25366_ (.A1(_01332_),
    .A2(_01813_),
    .A3(_01815_),
    .A4(_02170_),
    .B1(_02167_),
    .X(_02315_));
 sky130_fd_sc_hd__a31o_1 _25367_ (.A1(_02032_),
    .A2(_02049_),
    .A3(_02051_),
    .B1(_02055_),
    .X(_02316_));
 sky130_fd_sc_hd__o32a_2 _25368_ (.A1(_04896_),
    .A2(_08668_),
    .A3(_01801_),
    .B1(_02159_),
    .B2(_02156_),
    .X(_02317_));
 sky130_fd_sc_hd__a21oi_1 _25369_ (.A1(_02140_),
    .A2(_02151_),
    .B1(_02148_),
    .Y(_02318_));
 sky130_fd_sc_hd__o21ai_1 _25370_ (.A1(_02139_),
    .A2(_02150_),
    .B1(_02149_),
    .Y(_02319_));
 sky130_fd_sc_hd__or3b_1 _25371_ (.A(net49),
    .B(_04223_),
    .C_N(net48),
    .X(_02320_));
 sky130_fd_sc_hd__o211ai_4 _25372_ (.A1(net176),
    .A2(_07501_),
    .B1(net274),
    .C1(_07499_),
    .Y(_02321_));
 sky130_fd_sc_hd__nor2_1 _25373_ (.A(_04245_),
    .B(_05766_),
    .Y(_02323_));
 sky130_fd_sc_hd__or3b_1 _25374_ (.A(net48),
    .B(_04245_),
    .C_N(net47),
    .X(_02324_));
 sky130_fd_sc_hd__a211oi_2 _25375_ (.A1(net204),
    .A2(_07766_),
    .B1(_05763_),
    .C1(_07770_),
    .Y(_02325_));
 sky130_fd_sc_hd__o211ai_2 _25376_ (.A1(net170),
    .A2(_07765_),
    .B1(_05762_),
    .C1(_07771_),
    .Y(_02326_));
 sky130_fd_sc_hd__o2bb2a_1 _25377_ (.A1_N(_02320_),
    .A2_N(_02321_),
    .B1(_02323_),
    .B2(_02325_),
    .X(_02327_));
 sky130_fd_sc_hd__o2bb2ai_2 _25378_ (.A1_N(_02320_),
    .A2_N(_02321_),
    .B1(_02323_),
    .B2(_02325_),
    .Y(_02328_));
 sky130_fd_sc_hd__o2111ai_4 _25379_ (.A1(_04223_),
    .A2(_06030_),
    .B1(_02321_),
    .C1(_02324_),
    .D1(_02326_),
    .Y(_02329_));
 sky130_fd_sc_hd__o311a_1 _25380_ (.A1(net244),
    .A2(net241),
    .A3(_07074_),
    .B1(net273),
    .C1(_07072_),
    .X(_02330_));
 sky130_fd_sc_hd__and3_1 _25381_ (.A(_04190_),
    .B(net20),
    .C(net49),
    .X(_02331_));
 sky130_fd_sc_hd__a31o_1 _25382_ (.A1(_07072_),
    .A2(net170),
    .A3(net273),
    .B1(_02331_),
    .X(_02332_));
 sky130_fd_sc_hd__o211a_1 _25383_ (.A1(_02330_),
    .A2(_02331_),
    .B1(_02328_),
    .C1(_02329_),
    .X(_02334_));
 sky130_fd_sc_hd__o211ai_2 _25384_ (.A1(_02330_),
    .A2(_02331_),
    .B1(_02328_),
    .C1(_02329_),
    .Y(_02335_));
 sky130_fd_sc_hd__a21oi_1 _25385_ (.A1(_02328_),
    .A2(_02329_),
    .B1(_02332_),
    .Y(_02336_));
 sky130_fd_sc_hd__a211o_1 _25386_ (.A1(_02328_),
    .A2(_02329_),
    .B1(_02330_),
    .C1(_02331_),
    .X(_02337_));
 sky130_fd_sc_hd__and3_1 _25387_ (.A(_02319_),
    .B(_02335_),
    .C(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__nand3_1 _25388_ (.A(_02319_),
    .B(_02335_),
    .C(_02337_),
    .Y(_02339_));
 sky130_fd_sc_hd__o21ai_2 _25389_ (.A1(_02334_),
    .A2(_02336_),
    .B1(_02318_),
    .Y(_02340_));
 sky130_fd_sc_hd__o21ai_2 _25390_ (.A1(_02035_),
    .A2(_02046_),
    .B1(_02044_),
    .Y(_02341_));
 sky130_fd_sc_hd__a21oi_2 _25391_ (.A1(_02339_),
    .A2(_02340_),
    .B1(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__a21o_1 _25392_ (.A1(_02339_),
    .A2(_02340_),
    .B1(_02341_),
    .X(_02343_));
 sky130_fd_sc_hd__and3_2 _25393_ (.A(_02339_),
    .B(_02340_),
    .C(_02341_),
    .X(_02345_));
 sky130_fd_sc_hd__nand3_1 _25394_ (.A(_02339_),
    .B(_02340_),
    .C(_02341_),
    .Y(_02346_));
 sky130_fd_sc_hd__a21boi_1 _25395_ (.A1(_02343_),
    .A2(_02346_),
    .B1_N(_02317_),
    .Y(_02347_));
 sky130_fd_sc_hd__o21ai_4 _25396_ (.A1(_02342_),
    .A2(_02345_),
    .B1(_02317_),
    .Y(_02348_));
 sky130_fd_sc_hd__nor3_1 _25397_ (.A(_02317_),
    .B(_02342_),
    .C(_02345_),
    .Y(_02349_));
 sky130_fd_sc_hd__nand3b_2 _25398_ (.A_N(_02317_),
    .B(_02343_),
    .C(_02346_),
    .Y(_02350_));
 sky130_fd_sc_hd__o21bai_2 _25399_ (.A1(_02347_),
    .A2(_02349_),
    .B1_N(_02316_),
    .Y(_02351_));
 sky130_fd_sc_hd__nand3_1 _25400_ (.A(_02316_),
    .B(_02348_),
    .C(_02350_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand4_2 _25401_ (.A(_02053_),
    .B(_02056_),
    .C(_02348_),
    .D(_02350_),
    .Y(_02353_));
 sky130_fd_sc_hd__o2bb2ai_1 _25402_ (.A1_N(_02053_),
    .A2_N(_02056_),
    .B1(_02347_),
    .B2(_02349_),
    .Y(_02354_));
 sky130_fd_sc_hd__and3_1 _25403_ (.A(_02351_),
    .B(_02352_),
    .C(_02063_),
    .X(_02356_));
 sky130_fd_sc_hd__nand3_4 _25404_ (.A(_02351_),
    .B(_02352_),
    .C(_02063_),
    .Y(_02357_));
 sky130_fd_sc_hd__o2111ai_4 _25405_ (.A1(_02061_),
    .A2(_02025_),
    .B1(_02060_),
    .C1(_02353_),
    .D1(_02354_),
    .Y(_02358_));
 sky130_fd_sc_hd__inv_2 _25406_ (.A(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__or4_1 _25407_ (.A(net54),
    .B(_04266_),
    .C(_05548_),
    .D(net207),
    .X(_02360_));
 sky130_fd_sc_hd__or3b_2 _25408_ (.A(_04146_),
    .B(net56),
    .C_N(net54),
    .X(_02361_));
 sky130_fd_sc_hd__o31a_1 _25409_ (.A1(net54),
    .A2(_04266_),
    .A3(_05554_),
    .B1(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__a32o_1 _25410_ (.A1(net178),
    .A2(_05553_),
    .A3(net238),
    .B1(_08006_),
    .B2(net15),
    .X(_02363_));
 sky130_fd_sc_hd__a21boi_2 _25411_ (.A1(_01986_),
    .A2(_02002_),
    .B1_N(_02003_),
    .Y(_02364_));
 sky130_fd_sc_hd__a32o_1 _25412_ (.A1(net176),
    .A2(_05933_),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net16),
    .X(_02365_));
 sky130_fd_sc_hd__o21ai_1 _25413_ (.A1(_01988_),
    .A2(_01996_),
    .B1(_01995_),
    .Y(_02367_));
 sky130_fd_sc_hd__a32o_1 _25414_ (.A1(net202),
    .A2(net173),
    .A3(net239),
    .B1(_07308_),
    .B2(net17),
    .X(_02368_));
 sky130_fd_sc_hd__or3_1 _25415_ (.A(net51),
    .B(_04201_),
    .C(_04190_),
    .X(_02369_));
 sky130_fd_sc_hd__o211ai_4 _25416_ (.A1(net176),
    .A2(_06759_),
    .B1(net240),
    .C1(net191),
    .Y(_02370_));
 sky130_fd_sc_hd__nor2_1 _25417_ (.A(_04179_),
    .B(_07226_),
    .Y(_02371_));
 sky130_fd_sc_hd__o311a_1 _25418_ (.A1(net244),
    .A2(net241),
    .A3(_06451_),
    .B1(net269),
    .C1(net197),
    .X(_02372_));
 sky130_fd_sc_hd__a31oi_1 _25419_ (.A1(net197),
    .A2(_06452_),
    .A3(net269),
    .B1(_02371_),
    .Y(_02373_));
 sky130_fd_sc_hd__o2bb2ai_4 _25420_ (.A1_N(_02369_),
    .A2_N(_02370_),
    .B1(_02371_),
    .B2(_02372_),
    .Y(_02374_));
 sky130_fd_sc_hd__o211ai_2 _25421_ (.A1(_04201_),
    .A2(_06866_),
    .B1(_02370_),
    .C1(_02373_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand3_1 _25422_ (.A(_02368_),
    .B(_02374_),
    .C(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _25423_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_02368_),
    .X(_02378_));
 sky130_fd_sc_hd__a21bo_1 _25424_ (.A1(_02374_),
    .A2(_02375_),
    .B1_N(_02368_),
    .X(_02379_));
 sky130_fd_sc_hd__nand3b_1 _25425_ (.A_N(_02368_),
    .B(_02374_),
    .C(_02375_),
    .Y(_02380_));
 sky130_fd_sc_hd__nand3_1 _25426_ (.A(_02367_),
    .B(_02376_),
    .C(_02378_),
    .Y(_02381_));
 sky130_fd_sc_hd__nand4_2 _25427_ (.A(_01995_),
    .B(_01998_),
    .C(_02379_),
    .D(_02380_),
    .Y(_02382_));
 sky130_fd_sc_hd__nand3b_2 _25428_ (.A_N(_02365_),
    .B(_02381_),
    .C(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__a21bo_1 _25429_ (.A1(_02381_),
    .A2(_02382_),
    .B1_N(_02365_),
    .X(_02384_));
 sky130_fd_sc_hd__a21oi_4 _25430_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_02364_),
    .Y(_02385_));
 sky130_fd_sc_hd__and3_2 _25431_ (.A(_02384_),
    .B(_02364_),
    .C(_02383_),
    .X(_02386_));
 sky130_fd_sc_hd__nor2_1 _25432_ (.A(_02385_),
    .B(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__o221a_1 _25433_ (.A1(_04146_),
    .A2(_08007_),
    .B1(_02385_),
    .B2(_02386_),
    .C1(_02360_),
    .X(_02389_));
 sky130_fd_sc_hd__o21ai_1 _25434_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_02362_),
    .Y(_02390_));
 sky130_fd_sc_hd__a211oi_2 _25435_ (.A1(_02360_),
    .A2(_02361_),
    .B1(_02385_),
    .C1(_02386_),
    .Y(_02391_));
 sky130_fd_sc_hd__or3_1 _25436_ (.A(_02362_),
    .B(_02385_),
    .C(_02386_),
    .X(_02392_));
 sky130_fd_sc_hd__o2bb2a_1 _25437_ (.A1_N(_02360_),
    .A2_N(_02361_),
    .B1(_02385_),
    .B2(_02386_),
    .X(_02393_));
 sky130_fd_sc_hd__o21ai_1 _25438_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_02363_),
    .Y(_02394_));
 sky130_fd_sc_hd__o311a_1 _25439_ (.A1(net54),
    .A2(_04266_),
    .A3(_05554_),
    .B1(_02361_),
    .C1(_02387_),
    .X(_02395_));
 sky130_fd_sc_hd__or3_1 _25440_ (.A(_02363_),
    .B(_02385_),
    .C(_02386_),
    .X(_02396_));
 sky130_fd_sc_hd__nand4_4 _25441_ (.A(_02357_),
    .B(_02358_),
    .C(_02390_),
    .D(_02392_),
    .Y(_02397_));
 sky130_fd_sc_hd__inv_2 _25442_ (.A(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__o2bb2ai_1 _25443_ (.A1_N(_02357_),
    .A2_N(_02358_),
    .B1(_02389_),
    .B2(_02391_),
    .Y(_02400_));
 sky130_fd_sc_hd__o211ai_2 _25444_ (.A1(_02389_),
    .A2(_02391_),
    .B1(_02357_),
    .C1(_02358_),
    .Y(_02401_));
 sky130_fd_sc_hd__o2bb2ai_1 _25445_ (.A1_N(_02357_),
    .A2_N(_02358_),
    .B1(_02393_),
    .B2(_02395_),
    .Y(_02402_));
 sky130_fd_sc_hd__nand3_2 _25446_ (.A(_02400_),
    .B(_02315_),
    .C(_02397_),
    .Y(_02403_));
 sky130_fd_sc_hd__nand3b_4 _25447_ (.A_N(_02315_),
    .B(_02401_),
    .C(_02402_),
    .Y(_02404_));
 sky130_fd_sc_hd__inv_2 _25448_ (.A(_02404_),
    .Y(_02405_));
 sky130_fd_sc_hd__a22oi_1 _25449_ (.A1(_02072_),
    .A2(_02075_),
    .B1(_02403_),
    .B2(_02404_),
    .Y(_02406_));
 sky130_fd_sc_hd__and4_1 _25450_ (.A(_02072_),
    .B(_02075_),
    .C(_02403_),
    .D(_02404_),
    .X(_02407_));
 sky130_fd_sc_hd__o211a_1 _25451_ (.A1(_02071_),
    .A2(_02074_),
    .B1(_02403_),
    .C1(_02404_),
    .X(_02408_));
 sky130_fd_sc_hd__o211ai_2 _25452_ (.A1(_02071_),
    .A2(_02074_),
    .B1(_02403_),
    .C1(_02404_),
    .Y(_02409_));
 sky130_fd_sc_hd__a21oi_1 _25453_ (.A1(_02403_),
    .A2(_02404_),
    .B1(_02314_),
    .Y(_02411_));
 sky130_fd_sc_hd__a21o_1 _25454_ (.A1(_02403_),
    .A2(_02404_),
    .B1(_02314_),
    .X(_02412_));
 sky130_fd_sc_hd__nand4_1 _25455_ (.A(_02310_),
    .B(_02313_),
    .C(_02409_),
    .D(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__o2bb2ai_1 _25456_ (.A1_N(_02310_),
    .A2_N(_02313_),
    .B1(_02408_),
    .B2(_02411_),
    .Y(_02414_));
 sky130_fd_sc_hd__o211ai_1 _25457_ (.A1(_02408_),
    .A2(_02411_),
    .B1(_02310_),
    .C1(_02313_),
    .Y(_02415_));
 sky130_fd_sc_hd__o2bb2ai_1 _25458_ (.A1_N(_02310_),
    .A2_N(_02313_),
    .B1(_02406_),
    .B2(_02407_),
    .Y(_02416_));
 sky130_fd_sc_hd__o211ai_2 _25459_ (.A1(_02183_),
    .A2(_02209_),
    .B1(_02415_),
    .C1(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__and3_1 _25460_ (.A(_02414_),
    .B(_02210_),
    .C(_02413_),
    .X(_02418_));
 sky130_fd_sc_hd__nand3_1 _25461_ (.A(_02414_),
    .B(_02210_),
    .C(_02413_),
    .Y(_02419_));
 sky130_fd_sc_hd__and3_1 _25462_ (.A(_01926_),
    .B(_01931_),
    .C(_02079_),
    .X(_02420_));
 sky130_fd_sc_hd__o2bb2ai_2 _25463_ (.A1_N(_02417_),
    .A2_N(_02419_),
    .B1(_02420_),
    .B2(_02080_),
    .Y(_02422_));
 sky130_fd_sc_hd__o21ai_2 _25464_ (.A1(_02078_),
    .A2(_02084_),
    .B1(_02417_),
    .Y(_02423_));
 sky130_fd_sc_hd__o21ai_1 _25465_ (.A1(_02418_),
    .A2(_02423_),
    .B1(_02422_),
    .Y(_02424_));
 sky130_fd_sc_hd__a31o_1 _25466_ (.A1(_01978_),
    .A2(_02186_),
    .A3(_02187_),
    .B1(_01976_),
    .X(_02425_));
 sky130_fd_sc_hd__o2111ai_4 _25467_ (.A1(_02418_),
    .A2(_02423_),
    .B1(_02425_),
    .C1(_02422_),
    .D1(_02192_),
    .Y(_02426_));
 sky130_fd_sc_hd__o211ai_2 _25468_ (.A1(_02190_),
    .A2(_01977_),
    .B1(_02189_),
    .C1(_02424_),
    .Y(_02427_));
 sky130_fd_sc_hd__a31o_1 _25469_ (.A1(_02006_),
    .A2(_02008_),
    .A3(_02009_),
    .B1(_02018_),
    .X(_02428_));
 sky130_fd_sc_hd__a21oi_1 _25470_ (.A1(_02426_),
    .A2(_02427_),
    .B1(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__a221o_1 _25471_ (.A1(_01983_),
    .A2(_02012_),
    .B1(_02426_),
    .B2(_02427_),
    .C1(_02013_),
    .X(_02430_));
 sky130_fd_sc_hd__and3_1 _25472_ (.A(_02426_),
    .B(_02427_),
    .C(_02428_),
    .X(_02431_));
 sky130_fd_sc_hd__o221a_1 _25473_ (.A1(_01878_),
    .A2(_02197_),
    .B1(_02429_),
    .B2(_02431_),
    .C1(_02196_),
    .X(_02433_));
 sky130_fd_sc_hd__nand3b_1 _25474_ (.A_N(_02431_),
    .B(_02199_),
    .C(_02430_),
    .Y(_02434_));
 sky130_fd_sc_hd__and2b_1 _25475_ (.A_N(_02433_),
    .B(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__nand4_1 _25476_ (.A(_01967_),
    .B(_01969_),
    .C(_02204_),
    .D(_02206_),
    .Y(_02436_));
 sky130_fd_sc_hd__o221a_1 _25477_ (.A1(_02205_),
    .A2(_01969_),
    .B1(_01724_),
    .B2(_02436_),
    .C1(_02204_),
    .X(_02437_));
 sky130_fd_sc_hd__nor2_1 _25478_ (.A(_01723_),
    .B(_02436_),
    .Y(_02438_));
 sky130_fd_sc_hd__o221ai_2 _25479_ (.A1(_01479_),
    .A2(_01482_),
    .B1(_01481_),
    .B2(_12401_),
    .C1(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__nand2_1 _25480_ (.A(_02439_),
    .B(_02437_),
    .Y(_02440_));
 sky130_fd_sc_hd__xor2_1 _25481_ (.A(_02435_),
    .B(_02440_),
    .X(net112));
 sky130_fd_sc_hd__a21boi_1 _25482_ (.A1(_02427_),
    .A2(_02428_),
    .B1_N(_02426_),
    .Y(_02441_));
 sky130_fd_sc_hd__a31oi_2 _25483_ (.A1(_02310_),
    .A2(_02409_),
    .A3(_02412_),
    .B1(_02312_),
    .Y(_02443_));
 sky130_fd_sc_hd__a31o_1 _25484_ (.A1(_02310_),
    .A2(_02409_),
    .A3(_02412_),
    .B1(_02312_),
    .X(_02444_));
 sky130_fd_sc_hd__and3_1 _25485_ (.A(_02357_),
    .B(_02394_),
    .C(_02396_),
    .X(_02445_));
 sky130_fd_sc_hd__a21o_1 _25486_ (.A1(_02340_),
    .A2(_02341_),
    .B1(_02338_),
    .X(_02446_));
 sky130_fd_sc_hd__a22oi_2 _25487_ (.A1(net21),
    .A2(_06326_),
    .B1(_07504_),
    .B2(net273),
    .Y(_02447_));
 sky130_fd_sc_hd__a32oi_2 _25488_ (.A1(_07771_),
    .A2(net274),
    .A3(net166),
    .B1(_06029_),
    .B2(net22),
    .Y(_02448_));
 sky130_fd_sc_hd__a32o_1 _25489_ (.A1(_07771_),
    .A2(net274),
    .A3(net166),
    .B1(_06029_),
    .B2(net22),
    .X(_02449_));
 sky130_fd_sc_hd__nor2_2 _25490_ (.A(_04256_),
    .B(_05766_),
    .Y(_02450_));
 sky130_fd_sc_hd__o311a_1 _25491_ (.A1(_05931_),
    .A2(_07074_),
    .A3(net268),
    .B1(_05762_),
    .C1(net164),
    .X(_02451_));
 sky130_fd_sc_hd__a31oi_2 _25492_ (.A1(net164),
    .A2(_08208_),
    .A3(_05762_),
    .B1(_02450_),
    .Y(_02452_));
 sky130_fd_sc_hd__o21ai_4 _25493_ (.A1(_02450_),
    .A2(_02451_),
    .B1(_02449_),
    .Y(_02454_));
 sky130_fd_sc_hd__nand2_1 _25494_ (.A(_02448_),
    .B(_02452_),
    .Y(_02455_));
 sky130_fd_sc_hd__o21ai_1 _25495_ (.A1(_02450_),
    .A2(_02451_),
    .B1(_02448_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _25496_ (.A(_02449_),
    .B(_02452_),
    .Y(_02457_));
 sky130_fd_sc_hd__nand3b_4 _25497_ (.A_N(_02447_),
    .B(_02454_),
    .C(_02455_),
    .Y(_02458_));
 sky130_fd_sc_hd__nand3_2 _25498_ (.A(_02456_),
    .B(_02457_),
    .C(_02447_),
    .Y(_02459_));
 sky130_fd_sc_hd__nand2_2 _25499_ (.A(_02458_),
    .B(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__a21oi_1 _25500_ (.A1(_02272_),
    .A2(_02283_),
    .B1(_02280_),
    .Y(_02461_));
 sky130_fd_sc_hd__o21ai_1 _25501_ (.A1(_02271_),
    .A2(_02282_),
    .B1(_02281_),
    .Y(_02462_));
 sky130_fd_sc_hd__a21oi_4 _25502_ (.A1(_02458_),
    .A2(_02459_),
    .B1(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__a21oi_4 _25503_ (.A1(_02281_),
    .A2(_02284_),
    .B1(_02460_),
    .Y(_02465_));
 sky130_fd_sc_hd__a21o_1 _25504_ (.A1(_02281_),
    .A2(_02284_),
    .B1(_02460_),
    .X(_02466_));
 sky130_fd_sc_hd__a21oi_1 _25505_ (.A1(_02329_),
    .A2(_02332_),
    .B1(_02327_),
    .Y(_02467_));
 sky130_fd_sc_hd__nand3b_1 _25506_ (.A_N(_02463_),
    .B(_02466_),
    .C(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__o22ai_1 _25507_ (.A1(_02327_),
    .A2(_02334_),
    .B1(_02463_),
    .B2(_02465_),
    .Y(_02469_));
 sky130_fd_sc_hd__o21ai_1 _25508_ (.A1(_02463_),
    .A2(_02465_),
    .B1(_02467_),
    .Y(_02470_));
 sky130_fd_sc_hd__o2bb2a_2 _25509_ (.A1_N(_02461_),
    .A2_N(_02460_),
    .B1(_02334_),
    .B2(_02327_),
    .X(_02471_));
 sky130_fd_sc_hd__a22o_1 _25510_ (.A1(_02328_),
    .A2(_02335_),
    .B1(_02460_),
    .B2(_02461_),
    .X(_02472_));
 sky130_fd_sc_hd__nand3_2 _25511_ (.A(_02288_),
    .B(_02468_),
    .C(_02469_),
    .Y(_02473_));
 sky130_fd_sc_hd__o211ai_4 _25512_ (.A1(_02465_),
    .A2(_02472_),
    .B1(_02290_),
    .C1(_02470_),
    .Y(_02474_));
 sky130_fd_sc_hd__a21oi_1 _25513_ (.A1(_02473_),
    .A2(_02474_),
    .B1(_02446_),
    .Y(_02476_));
 sky130_fd_sc_hd__a21o_1 _25514_ (.A1(_02473_),
    .A2(_02474_),
    .B1(_02446_),
    .X(_02477_));
 sky130_fd_sc_hd__o211a_1 _25515_ (.A1(_02338_),
    .A2(_02345_),
    .B1(_02473_),
    .C1(_02474_),
    .X(_02478_));
 sky130_fd_sc_hd__o211ai_2 _25516_ (.A1(_02338_),
    .A2(_02345_),
    .B1(_02473_),
    .C1(_02474_),
    .Y(_02479_));
 sky130_fd_sc_hd__o211ai_2 _25517_ (.A1(_02047_),
    .A2(_02052_),
    .B1(_02056_),
    .C1(_02350_),
    .Y(_02480_));
 sky130_fd_sc_hd__a21oi_1 _25518_ (.A1(_02316_),
    .A2(_02348_),
    .B1(_02349_),
    .Y(_02481_));
 sky130_fd_sc_hd__nand4_4 _25519_ (.A(_02348_),
    .B(_02477_),
    .C(_02479_),
    .D(_02480_),
    .Y(_02482_));
 sky130_fd_sc_hd__o21ai_2 _25520_ (.A1(_02476_),
    .A2(_02478_),
    .B1(_02481_),
    .Y(_02483_));
 sky130_fd_sc_hd__o2bb2a_1 _25521_ (.A1_N(_05934_),
    .A2_N(net238),
    .B1(_08007_),
    .B2(_04157_),
    .X(_02484_));
 sky130_fd_sc_hd__a32o_1 _25522_ (.A1(net202),
    .A2(_06221_),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net17),
    .X(_02485_));
 sky130_fd_sc_hd__nand2_1 _25523_ (.A(_02374_),
    .B(_02376_),
    .Y(_02487_));
 sky130_fd_sc_hd__a32o_1 _25524_ (.A1(_06449_),
    .A2(_06452_),
    .A3(net239),
    .B1(_07308_),
    .B2(net18),
    .X(_02488_));
 sky130_fd_sc_hd__or3_1 _25525_ (.A(net51),
    .B(_04212_),
    .C(_04190_),
    .X(_02489_));
 sky130_fd_sc_hd__o221ai_4 _25526_ (.A1(net176),
    .A2(_07074_),
    .B1(_04212_),
    .B2(net190),
    .C1(net240),
    .Y(_02490_));
 sky130_fd_sc_hd__o31a_1 _25527_ (.A1(_04190_),
    .A2(net51),
    .A3(_04212_),
    .B1(_02490_),
    .X(_02491_));
 sky130_fd_sc_hd__nor2_1 _25528_ (.A(_04201_),
    .B(_07226_),
    .Y(_02492_));
 sky130_fd_sc_hd__o311a_1 _25529_ (.A1(net244),
    .A2(net241),
    .A3(_06759_),
    .B1(net269),
    .C1(net192),
    .X(_02493_));
 sky130_fd_sc_hd__a31oi_4 _25530_ (.A1(net192),
    .A2(_06762_),
    .A3(net269),
    .B1(_02492_),
    .Y(_02494_));
 sky130_fd_sc_hd__o2bb2ai_2 _25531_ (.A1_N(_02489_),
    .A2_N(_02490_),
    .B1(_02492_),
    .B2(_02493_),
    .Y(_02495_));
 sky130_fd_sc_hd__o211ai_4 _25532_ (.A1(_04212_),
    .A2(_06866_),
    .B1(_02490_),
    .C1(_02494_),
    .Y(_02496_));
 sky130_fd_sc_hd__nand3_2 _25533_ (.A(_02488_),
    .B(_02495_),
    .C(_02496_),
    .Y(_02498_));
 sky130_fd_sc_hd__a21o_1 _25534_ (.A1(_02495_),
    .A2(_02496_),
    .B1(_02488_),
    .X(_02499_));
 sky130_fd_sc_hd__a21bo_1 _25535_ (.A1(_02495_),
    .A2(_02496_),
    .B1_N(_02488_),
    .X(_02500_));
 sky130_fd_sc_hd__nand3b_1 _25536_ (.A_N(_02488_),
    .B(_02495_),
    .C(_02496_),
    .Y(_02501_));
 sky130_fd_sc_hd__nand3_1 _25537_ (.A(_02487_),
    .B(_02498_),
    .C(_02499_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand4_1 _25538_ (.A(_02374_),
    .B(_02376_),
    .C(_02500_),
    .D(_02501_),
    .Y(_02503_));
 sky130_fd_sc_hd__a21bo_1 _25539_ (.A1(_02502_),
    .A2(_02503_),
    .B1_N(_02485_),
    .X(_02504_));
 sky130_fd_sc_hd__nand3b_1 _25540_ (.A_N(_02485_),
    .B(_02502_),
    .C(_02503_),
    .Y(_02505_));
 sky130_fd_sc_hd__a21boi_1 _25541_ (.A1(_02365_),
    .A2(_02382_),
    .B1_N(_02381_),
    .Y(_02506_));
 sky130_fd_sc_hd__a21o_1 _25542_ (.A1(_02504_),
    .A2(_02505_),
    .B1(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__nand3_1 _25543_ (.A(_02504_),
    .B(_02505_),
    .C(_02506_),
    .Y(_02509_));
 sky130_fd_sc_hd__nand2_1 _25544_ (.A(_02507_),
    .B(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__and2_1 _25545_ (.A(_02510_),
    .B(_02484_),
    .X(_02511_));
 sky130_fd_sc_hd__nor2_1 _25546_ (.A(_02484_),
    .B(_02510_),
    .Y(_02512_));
 sky130_fd_sc_hd__and3_1 _25547_ (.A(_02507_),
    .B(_02509_),
    .C(_02484_),
    .X(_02513_));
 sky130_fd_sc_hd__a21oi_1 _25548_ (.A1(_02507_),
    .A2(_02509_),
    .B1(_02484_),
    .Y(_02514_));
 sky130_fd_sc_hd__o2bb2ai_2 _25549_ (.A1_N(_02482_),
    .A2_N(_02483_),
    .B1(_02511_),
    .B2(_02512_),
    .Y(_02515_));
 sky130_fd_sc_hd__o211ai_4 _25550_ (.A1(_02513_),
    .A2(_02514_),
    .B1(_02482_),
    .C1(_02483_),
    .Y(_02516_));
 sky130_fd_sc_hd__and4_1 _25551_ (.A(_01332_),
    .B(_02162_),
    .C(_02163_),
    .D(_02294_),
    .X(_02517_));
 sky130_fd_sc_hd__a41o_1 _25552_ (.A1(_01332_),
    .A2(_02162_),
    .A3(_02163_),
    .A4(_02294_),
    .B1(_02295_),
    .X(_02518_));
 sky130_fd_sc_hd__o211a_1 _25553_ (.A1(_02295_),
    .A2(_02517_),
    .B1(_02516_),
    .C1(_02515_),
    .X(_02520_));
 sky130_fd_sc_hd__o211ai_4 _25554_ (.A1(_02295_),
    .A2(_02517_),
    .B1(_02516_),
    .C1(_02515_),
    .Y(_02521_));
 sky130_fd_sc_hd__a21oi_2 _25555_ (.A1(_02515_),
    .A2(_02516_),
    .B1(_02518_),
    .Y(_02522_));
 sky130_fd_sc_hd__a21o_1 _25556_ (.A1(_02515_),
    .A2(_02516_),
    .B1(_02518_),
    .X(_02523_));
 sky130_fd_sc_hd__o211ai_4 _25557_ (.A1(_02359_),
    .A2(_02445_),
    .B1(_02521_),
    .C1(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__o22ai_4 _25558_ (.A1(_02356_),
    .A2(_02398_),
    .B1(_02520_),
    .B2(_02522_),
    .Y(_02525_));
 sky130_fd_sc_hd__o211a_1 _25559_ (.A1(_02356_),
    .A2(_02398_),
    .B1(_02521_),
    .C1(_02523_),
    .X(_02526_));
 sky130_fd_sc_hd__a211o_1 _25560_ (.A1(_02357_),
    .A2(_02397_),
    .B1(_02520_),
    .C1(_02522_),
    .X(_02527_));
 sky130_fd_sc_hd__o22a_1 _25561_ (.A1(_02359_),
    .A2(_02445_),
    .B1(_02520_),
    .B2(_02522_),
    .X(_02528_));
 sky130_fd_sc_hd__a2bb2o_1 _25562_ (.A1_N(_02359_),
    .A2_N(_02445_),
    .B1(_02521_),
    .B2(_02523_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _25563_ (.A(_02524_),
    .B(_02525_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_2 _25564_ (.A(net319),
    .B(_05465_),
    .Y(_02532_));
 sky130_fd_sc_hd__a21oi_1 _25565_ (.A1(net153),
    .A2(net158),
    .B1(_05463_),
    .Y(_02533_));
 sky130_fd_sc_hd__a21oi_2 _25566_ (.A1(_08670_),
    .A2(_05462_),
    .B1(_02532_),
    .Y(_02534_));
 sky130_fd_sc_hd__o211ai_4 _25567_ (.A1(net170),
    .A2(net268),
    .B1(net319),
    .C1(_05225_),
    .Y(_02535_));
 sky130_fd_sc_hd__and4_4 _25568_ (.A(_02146_),
    .B(_02273_),
    .C(_02279_),
    .D(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__o2111ai_4 _25569_ (.A1(_04986_),
    .A2(net153),
    .B1(_02146_),
    .C1(_02279_),
    .D1(_02535_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2_1 _25570_ (.A(_02534_),
    .B(_02536_),
    .Y(_02538_));
 sky130_fd_sc_hd__o21a_2 _25571_ (.A1(_02532_),
    .A2(_02533_),
    .B1(_02537_),
    .X(_02539_));
 sky130_fd_sc_hd__o21ai_2 _25572_ (.A1(_02532_),
    .A2(_02533_),
    .B1(_02537_),
    .Y(_02540_));
 sky130_fd_sc_hd__a21o_2 _25573_ (.A1(_02538_),
    .A2(_02540_),
    .B1(_02160_),
    .X(_02542_));
 sky130_fd_sc_hd__and3_1 _25574_ (.A(_02160_),
    .B(_02538_),
    .C(_02540_),
    .X(_02543_));
 sky130_fd_sc_hd__nand3_4 _25575_ (.A(_02160_),
    .B(_02538_),
    .C(_02540_),
    .Y(_02544_));
 sky130_fd_sc_hd__o211ai_4 _25576_ (.A1(_00796_),
    .A2(_01324_),
    .B1(_02542_),
    .C1(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__o2bb2ai_2 _25577_ (.A1_N(_02542_),
    .A2_N(_02544_),
    .B1(_00796_),
    .B2(_01324_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand3_1 _25578_ (.A(_02542_),
    .B(_02544_),
    .C(_01331_),
    .Y(_02547_));
 sky130_fd_sc_hd__a221o_1 _25579_ (.A1(_13065_),
    .A2(_00358_),
    .B1(_02546_),
    .B2(_02547_),
    .C1(_11741_),
    .X(_02548_));
 sky130_fd_sc_hd__inv_2 _25580_ (.A(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__o211ai_2 _25581_ (.A1(_00360_),
    .A2(_11741_),
    .B1(_02547_),
    .C1(_02546_),
    .Y(_02550_));
 sky130_fd_sc_hd__a2bb2o_1 _25582_ (.A1_N(_00360_),
    .A2_N(_11741_),
    .B1(_02547_),
    .B2(_02546_),
    .X(_02551_));
 sky130_fd_sc_hd__nand4_1 _25583_ (.A(_00361_),
    .B(_02546_),
    .C(_02547_),
    .D(_11740_),
    .Y(_02553_));
 sky130_fd_sc_hd__nand2_1 _25584_ (.A(_02551_),
    .B(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__and3_1 _25585_ (.A(_02548_),
    .B(_02550_),
    .C(_02293_),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _25586_ (.A(_02293_),
    .B(_02554_),
    .Y(_02556_));
 sky130_fd_sc_hd__a31o_1 _25587_ (.A1(_01332_),
    .A2(_02288_),
    .A3(_02291_),
    .B1(_02554_),
    .X(_02557_));
 sky130_fd_sc_hd__nand2_1 _25588_ (.A(_02556_),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__a21oi_1 _25589_ (.A1(_02261_),
    .A2(_00736_),
    .B1(_02258_),
    .Y(_02559_));
 sky130_fd_sc_hd__o21ai_1 _25590_ (.A1(net129),
    .A2(_02260_),
    .B1(_02259_),
    .Y(_02560_));
 sky130_fd_sc_hd__a21oi_2 _25591_ (.A1(_12099_),
    .A2(_02248_),
    .B1(_02249_),
    .Y(_02561_));
 sky130_fd_sc_hd__or3_2 _25592_ (.A(net57),
    .B(_04266_),
    .C(_04146_),
    .X(_02562_));
 sky130_fd_sc_hd__nand3_2 _25593_ (.A(net178),
    .B(_05553_),
    .C(_08657_),
    .Y(_02564_));
 sky130_fd_sc_hd__o21ai_1 _25594_ (.A1(_04146_),
    .A2(_08660_),
    .B1(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__a21oi_1 _25595_ (.A1(_02562_),
    .A2(_02564_),
    .B1(net149),
    .Y(_02566_));
 sky130_fd_sc_hd__a21o_1 _25596_ (.A1(_02562_),
    .A2(_02564_),
    .B1(net149),
    .X(_02567_));
 sky130_fd_sc_hd__o311a_4 _25597_ (.A1(_08658_),
    .A2(net207),
    .A3(_05548_),
    .B1(_02562_),
    .C1(net149),
    .X(_02568_));
 sky130_fd_sc_hd__a31o_1 _25598_ (.A1(net149),
    .A2(_02562_),
    .A3(_02564_),
    .B1(net145),
    .X(_02569_));
 sky130_fd_sc_hd__o21ai_2 _25599_ (.A1(_02566_),
    .A2(_02568_),
    .B1(net145),
    .Y(_02570_));
 sky130_fd_sc_hd__o21ai_2 _25600_ (.A1(_02566_),
    .A2(_02568_),
    .B1(net144),
    .Y(_02571_));
 sky130_fd_sc_hd__nand3b_2 _25601_ (.A_N(_02568_),
    .B(net145),
    .C(_02567_),
    .Y(_02572_));
 sky130_fd_sc_hd__o21ai_4 _25602_ (.A1(net145),
    .A2(_02224_),
    .B1(_02222_),
    .Y(_02573_));
 sky130_fd_sc_hd__a21oi_2 _25603_ (.A1(net144),
    .A2(_02225_),
    .B1(_02221_),
    .Y(_02575_));
 sky130_fd_sc_hd__o211a_2 _25604_ (.A1(net145),
    .A2(_02568_),
    .B1(_02573_),
    .C1(_02570_),
    .X(_02576_));
 sky130_fd_sc_hd__o211ai_4 _25605_ (.A1(net145),
    .A2(_02568_),
    .B1(_02573_),
    .C1(_02570_),
    .Y(_02577_));
 sky130_fd_sc_hd__and3_1 _25606_ (.A(_02571_),
    .B(_02572_),
    .C(_02575_),
    .X(_02578_));
 sky130_fd_sc_hd__nand3_2 _25607_ (.A(_02571_),
    .B(_02572_),
    .C(_02575_),
    .Y(_02579_));
 sky130_fd_sc_hd__a22o_1 _25608_ (.A1(net139),
    .A2(_10544_),
    .B1(_02577_),
    .B2(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__a31oi_2 _25609_ (.A1(_02571_),
    .A2(_02572_),
    .A3(_02575_),
    .B1(_10546_),
    .Y(_02581_));
 sky130_fd_sc_hd__a31o_1 _25610_ (.A1(_02571_),
    .A2(_02572_),
    .A3(_02575_),
    .B1(_10546_),
    .X(_02582_));
 sky130_fd_sc_hd__o211ai_4 _25611_ (.A1(net140),
    .A2(net136),
    .B1(_02577_),
    .C1(_02579_),
    .Y(_02583_));
 sky130_fd_sc_hd__a21o_1 _25612_ (.A1(_02577_),
    .A2(_02579_),
    .B1(_10546_),
    .X(_02584_));
 sky130_fd_sc_hd__o211ai_4 _25613_ (.A1(_02233_),
    .A2(_02240_),
    .B1(_02583_),
    .C1(_02584_),
    .Y(_02586_));
 sky130_fd_sc_hd__o221a_1 _25614_ (.A1(_02231_),
    .A2(_02241_),
    .B1(_02576_),
    .B2(_02582_),
    .C1(_02580_),
    .X(_02587_));
 sky130_fd_sc_hd__o221ai_4 _25615_ (.A1(_02231_),
    .A2(_02241_),
    .B1(_02576_),
    .B2(_02582_),
    .C1(_02580_),
    .Y(_02588_));
 sky130_fd_sc_hd__o2bb2ai_2 _25616_ (.A1_N(_02586_),
    .A2_N(_02588_),
    .B1(net141),
    .B2(_11742_),
    .Y(_02589_));
 sky130_fd_sc_hd__o2111ai_4 _25617_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net143),
    .C1(_02586_),
    .D1(_02588_),
    .Y(_02590_));
 sky130_fd_sc_hd__a21o_1 _25618_ (.A1(_02586_),
    .A2(_02588_),
    .B1(_12099_),
    .X(_02591_));
 sky130_fd_sc_hd__a31o_1 _25619_ (.A1(_02243_),
    .A2(_02583_),
    .A3(_02584_),
    .B1(net132),
    .X(_02592_));
 sky130_fd_sc_hd__a21oi_4 _25620_ (.A1(_02589_),
    .A2(_02590_),
    .B1(_02561_),
    .Y(_02593_));
 sky130_fd_sc_hd__o221ai_4 _25621_ (.A1(_02249_),
    .A2(_02253_),
    .B1(_02587_),
    .B2(_02592_),
    .C1(_02591_),
    .Y(_02594_));
 sky130_fd_sc_hd__nand3_2 _25622_ (.A(_02561_),
    .B(_02589_),
    .C(_02590_),
    .Y(_02595_));
 sky130_fd_sc_hd__o211a_1 _25623_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_02595_),
    .X(_02597_));
 sky130_fd_sc_hd__a31o_1 _25624_ (.A1(_02561_),
    .A2(_02589_),
    .A3(_02590_),
    .B1(net129),
    .X(_02598_));
 sky130_fd_sc_hd__a22o_1 _25625_ (.A1(_00364_),
    .A2(_00367_),
    .B1(_02594_),
    .B2(_02595_),
    .X(_02599_));
 sky130_fd_sc_hd__o211ai_2 _25626_ (.A1(_00363_),
    .A2(_00366_),
    .B1(_02594_),
    .C1(_02595_),
    .Y(_02600_));
 sky130_fd_sc_hd__a21o_1 _25627_ (.A1(_02594_),
    .A2(_02595_),
    .B1(net129),
    .X(_02601_));
 sky130_fd_sc_hd__o211a_1 _25628_ (.A1(_02598_),
    .A2(_02593_),
    .B1(_02560_),
    .C1(_02599_),
    .X(_02602_));
 sky130_fd_sc_hd__o211ai_2 _25629_ (.A1(_02598_),
    .A2(_02593_),
    .B1(_02560_),
    .C1(_02599_),
    .Y(_02603_));
 sky130_fd_sc_hd__nand3_2 _25630_ (.A(_02601_),
    .B(_02559_),
    .C(_02600_),
    .Y(_02604_));
 sky130_fd_sc_hd__a31o_1 _25631_ (.A1(_02601_),
    .A2(_02559_),
    .A3(_02600_),
    .B1(_02558_),
    .X(_02605_));
 sky130_fd_sc_hd__a22o_1 _25632_ (.A1(_02556_),
    .A2(_02557_),
    .B1(_02603_),
    .B2(_02604_),
    .X(_02606_));
 sky130_fd_sc_hd__nand3_1 _25633_ (.A(_02558_),
    .B(_02603_),
    .C(_02604_),
    .Y(_02608_));
 sky130_fd_sc_hd__a21o_1 _25634_ (.A1(_02603_),
    .A2(_02604_),
    .B1(_02558_),
    .X(_02609_));
 sky130_fd_sc_hd__o21a_1 _25635_ (.A1(_02602_),
    .A2(_02605_),
    .B1(_02606_),
    .X(_02610_));
 sky130_fd_sc_hd__a31oi_4 _25636_ (.A1(_02268_),
    .A2(_02302_),
    .A3(_02304_),
    .B1(_02269_),
    .Y(_02611_));
 sky130_fd_sc_hd__a2bb2oi_2 _25637_ (.A1_N(_02262_),
    .A2_N(_02266_),
    .B1(_02305_),
    .B2(_02270_),
    .Y(_02612_));
 sky130_fd_sc_hd__nand3_4 _25638_ (.A(_02608_),
    .B(_02609_),
    .C(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__o211ai_4 _25639_ (.A1(_02602_),
    .A2(_02605_),
    .B1(_02611_),
    .C1(_02606_),
    .Y(_02614_));
 sky130_fd_sc_hd__nand3_4 _25640_ (.A(_02524_),
    .B(_02525_),
    .C(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__o21a_1 _25641_ (.A1(_02610_),
    .A2(_02611_),
    .B1(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__nand2_1 _25642_ (.A(_02613_),
    .B(_02614_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand4_1 _25643_ (.A(_02524_),
    .B(_02525_),
    .C(_02613_),
    .D(_02614_),
    .Y(_02619_));
 sky130_fd_sc_hd__nand2_1 _25644_ (.A(_02531_),
    .B(_02617_),
    .Y(_02620_));
 sky130_fd_sc_hd__o21ai_1 _25645_ (.A1(_02526_),
    .A2(_02528_),
    .B1(_02617_),
    .Y(_02621_));
 sky130_fd_sc_hd__nand4_1 _25646_ (.A(_02527_),
    .B(_02529_),
    .C(_02613_),
    .D(_02614_),
    .Y(_02622_));
 sky130_fd_sc_hd__nand3_1 _25647_ (.A(_02620_),
    .B(_02443_),
    .C(_02619_),
    .Y(_02623_));
 sky130_fd_sc_hd__a21oi_1 _25648_ (.A1(_02619_),
    .A2(_02620_),
    .B1(_02443_),
    .Y(_02624_));
 sky130_fd_sc_hd__nand3_1 _25649_ (.A(_02444_),
    .B(_02621_),
    .C(_02622_),
    .Y(_02625_));
 sky130_fd_sc_hd__and3_1 _25650_ (.A(_02072_),
    .B(_02075_),
    .C(_02403_),
    .X(_02626_));
 sky130_fd_sc_hd__a31o_1 _25651_ (.A1(_02315_),
    .A2(_02397_),
    .A3(_02400_),
    .B1(_02408_),
    .X(_02627_));
 sky130_fd_sc_hd__o2bb2ai_1 _25652_ (.A1_N(_02623_),
    .A2_N(_02625_),
    .B1(_02626_),
    .B2(_02405_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand3_1 _25653_ (.A(_02623_),
    .B(_02625_),
    .C(_02627_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2_1 _25654_ (.A(_02419_),
    .B(_02423_),
    .Y(_02631_));
 sky130_fd_sc_hd__nand3_2 _25655_ (.A(_02628_),
    .B(_02631_),
    .C(_02630_),
    .Y(_02632_));
 sky130_fd_sc_hd__a21o_1 _25656_ (.A1(_02628_),
    .A2(_02630_),
    .B1(_02631_),
    .X(_02633_));
 sky130_fd_sc_hd__o21ai_1 _25657_ (.A1(_02385_),
    .A2(_02391_),
    .B1(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__a221oi_2 _25658_ (.A1(_02387_),
    .A2(_02363_),
    .B1(_02633_),
    .B2(_02632_),
    .C1(_02385_),
    .Y(_02635_));
 sky130_fd_sc_hd__o211a_1 _25659_ (.A1(_02385_),
    .A2(_02391_),
    .B1(_02632_),
    .C1(_02633_),
    .X(_02636_));
 sky130_fd_sc_hd__nor3_1 _25660_ (.A(_02636_),
    .B(_02441_),
    .C(_02635_),
    .Y(_02637_));
 sky130_fd_sc_hd__o21a_1 _25661_ (.A1(_02635_),
    .A2(_02636_),
    .B1(_02441_),
    .X(_02638_));
 sky130_fd_sc_hd__nor2_1 _25662_ (.A(_02637_),
    .B(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hd__a31o_1 _25663_ (.A1(_02434_),
    .A2(_02439_),
    .A3(_02437_),
    .B1(_02433_),
    .X(_02641_));
 sky130_fd_sc_hd__xnor2_1 _25664_ (.A(_02639_),
    .B(_02641_),
    .Y(net113));
 sky130_fd_sc_hd__o21ai_1 _25665_ (.A1(_02484_),
    .A2(_02510_),
    .B1(_02507_),
    .Y(_02642_));
 sky130_fd_sc_hd__o21a_1 _25666_ (.A1(_02484_),
    .A2(_02510_),
    .B1(_02507_),
    .X(_02643_));
 sky130_fd_sc_hd__a21o_1 _25667_ (.A1(_02623_),
    .A2(_02627_),
    .B1(_02624_),
    .X(_02644_));
 sky130_fd_sc_hd__a21oi_1 _25668_ (.A1(_02623_),
    .A2(_02627_),
    .B1(_02624_),
    .Y(_02645_));
 sky130_fd_sc_hd__a31oi_2 _25669_ (.A1(_02569_),
    .A2(_02570_),
    .A3(_02573_),
    .B1(_10545_),
    .Y(_02646_));
 sky130_fd_sc_hd__a21oi_1 _25670_ (.A1(_02565_),
    .A2(net157),
    .B1(net144),
    .Y(_02647_));
 sky130_fd_sc_hd__o21ai_1 _25671_ (.A1(net145),
    .A2(_02568_),
    .B1(_02567_),
    .Y(_02648_));
 sky130_fd_sc_hd__o21a_1 _25672_ (.A1(net145),
    .A2(_02568_),
    .B1(_02567_),
    .X(_02649_));
 sky130_fd_sc_hd__o211ai_4 _25673_ (.A1(net233),
    .A2(_05927_),
    .B1(_08657_),
    .C1(_05933_),
    .Y(_02651_));
 sky130_fd_sc_hd__or3_2 _25674_ (.A(net57),
    .B(_04266_),
    .C(_04157_),
    .X(_02652_));
 sky130_fd_sc_hd__o31ai_4 _25675_ (.A1(net204),
    .A2(_08658_),
    .A3(_05932_),
    .B1(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__a21oi_2 _25676_ (.A1(_02651_),
    .A2(_02652_),
    .B1(net149),
    .Y(_02654_));
 sky130_fd_sc_hd__a21o_1 _25677_ (.A1(_02651_),
    .A2(_02652_),
    .B1(net149),
    .X(_02655_));
 sky130_fd_sc_hd__o311a_4 _25678_ (.A1(_04157_),
    .A2(_04266_),
    .A3(net57),
    .B1(net149),
    .C1(_02651_),
    .X(_02656_));
 sky130_fd_sc_hd__o221ai_4 _25679_ (.A1(_05935_),
    .A2(_08658_),
    .B1(_08660_),
    .B2(_04157_),
    .C1(net149),
    .Y(_02657_));
 sky130_fd_sc_hd__nand3_4 _25680_ (.A(_02655_),
    .B(_02657_),
    .C(net145),
    .Y(_02658_));
 sky130_fd_sc_hd__o22ai_4 _25681_ (.A1(net237),
    .A2(_09297_),
    .B1(_02654_),
    .B2(_02656_),
    .Y(_02659_));
 sky130_fd_sc_hd__o21ai_1 _25682_ (.A1(_02654_),
    .A2(_02656_),
    .B1(net145),
    .Y(_02660_));
 sky130_fd_sc_hd__o211ai_4 _25683_ (.A1(net145),
    .A2(_02656_),
    .B1(_02648_),
    .C1(_02660_),
    .Y(_02662_));
 sky130_fd_sc_hd__o211ai_4 _25684_ (.A1(_02568_),
    .A2(_02647_),
    .B1(_02658_),
    .C1(_02659_),
    .Y(_02663_));
 sky130_fd_sc_hd__a21oi_2 _25685_ (.A1(_02662_),
    .A2(_02663_),
    .B1(_10545_),
    .Y(_02664_));
 sky130_fd_sc_hd__a22o_1 _25686_ (.A1(net139),
    .A2(_10544_),
    .B1(_02662_),
    .B2(_02663_),
    .X(_02665_));
 sky130_fd_sc_hd__nand4_2 _25687_ (.A(net139),
    .B(_10544_),
    .C(_02662_),
    .D(_02663_),
    .Y(_02666_));
 sky130_fd_sc_hd__o211ai_2 _25688_ (.A1(net140),
    .A2(net136),
    .B1(_02662_),
    .C1(_02663_),
    .Y(_02667_));
 sky130_fd_sc_hd__a21o_1 _25689_ (.A1(_02662_),
    .A2(_02663_),
    .B1(_10546_),
    .X(_02668_));
 sky130_fd_sc_hd__o21ai_2 _25690_ (.A1(_02576_),
    .A2(_02581_),
    .B1(_02666_),
    .Y(_02669_));
 sky130_fd_sc_hd__o211ai_2 _25691_ (.A1(_02576_),
    .A2(_02581_),
    .B1(_02665_),
    .C1(_02666_),
    .Y(_02670_));
 sky130_fd_sc_hd__o211ai_4 _25692_ (.A1(_02578_),
    .A2(_02646_),
    .B1(_02667_),
    .C1(_02668_),
    .Y(_02671_));
 sky130_fd_sc_hd__a21oi_2 _25693_ (.A1(_02670_),
    .A2(_02671_),
    .B1(_12099_),
    .Y(_02673_));
 sky130_fd_sc_hd__a21o_1 _25694_ (.A1(_02670_),
    .A2(_02671_),
    .B1(_12099_),
    .X(_02674_));
 sky130_fd_sc_hd__o221a_1 _25695_ (.A1(net141),
    .A2(_11742_),
    .B1(_02664_),
    .B2(_02669_),
    .C1(_02671_),
    .X(_02675_));
 sky130_fd_sc_hd__o221ai_4 _25696_ (.A1(net141),
    .A2(_11742_),
    .B1(_02664_),
    .B2(_02669_),
    .C1(_02671_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _25697_ (.A(_02674_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__a32oi_2 _25698_ (.A1(_02243_),
    .A2(_02583_),
    .A3(_02584_),
    .B1(_02588_),
    .B2(net132),
    .Y(_02678_));
 sky130_fd_sc_hd__a32o_2 _25699_ (.A1(_02243_),
    .A2(_02583_),
    .A3(_02584_),
    .B1(_02588_),
    .B2(net132),
    .X(_02679_));
 sky130_fd_sc_hd__a21oi_1 _25700_ (.A1(_02674_),
    .A2(_02676_),
    .B1(_02678_),
    .Y(_02680_));
 sky130_fd_sc_hd__o21ai_2 _25701_ (.A1(_02673_),
    .A2(_02675_),
    .B1(_02679_),
    .Y(_02681_));
 sky130_fd_sc_hd__nor3_4 _25702_ (.A(_02673_),
    .B(_02675_),
    .C(_02679_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand3_1 _25703_ (.A(_02674_),
    .B(_02676_),
    .C(_02678_),
    .Y(_02684_));
 sky130_fd_sc_hd__o22ai_4 _25704_ (.A1(_00363_),
    .A2(_00366_),
    .B1(_02680_),
    .B2(_02682_),
    .Y(_02685_));
 sky130_fd_sc_hd__a21oi_2 _25705_ (.A1(_02677_),
    .A2(_02679_),
    .B1(net129),
    .Y(_02686_));
 sky130_fd_sc_hd__o2111ai_4 _25706_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_02681_),
    .D1(_02684_),
    .Y(_02687_));
 sky130_fd_sc_hd__nand2_1 _25707_ (.A(_02685_),
    .B(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__a31o_1 _25708_ (.A1(_00364_),
    .A2(_00367_),
    .A3(_02595_),
    .B1(_02593_),
    .X(_02689_));
 sky130_fd_sc_hd__a32o_1 _25709_ (.A1(_02561_),
    .A2(_02589_),
    .A3(_02590_),
    .B1(_02594_),
    .B2(net129),
    .X(_02690_));
 sky130_fd_sc_hd__a21oi_2 _25710_ (.A1(_02685_),
    .A2(_02687_),
    .B1(_02689_),
    .Y(_02691_));
 sky130_fd_sc_hd__a21o_1 _25711_ (.A1(_02685_),
    .A2(_02687_),
    .B1(_02689_),
    .X(_02692_));
 sky130_fd_sc_hd__o211a_2 _25712_ (.A1(_02593_),
    .A2(_02597_),
    .B1(_02685_),
    .C1(_02687_),
    .X(_02693_));
 sky130_fd_sc_hd__o211ai_4 _25713_ (.A1(_02593_),
    .A2(_02597_),
    .B1(_02685_),
    .C1(_02687_),
    .Y(_02695_));
 sky130_fd_sc_hd__a31oi_4 _25714_ (.A1(net319),
    .A2(_08208_),
    .A3(_05462_),
    .B1(_02532_),
    .Y(_02696_));
 sky130_fd_sc_hd__o2111a_1 _25715_ (.A1(_05226_),
    .A2(net153),
    .B1(_02279_),
    .C1(_02696_),
    .D1(_02274_),
    .X(_02697_));
 sky130_fd_sc_hd__a311o_1 _25716_ (.A1(net319),
    .A2(_05462_),
    .A3(_08208_),
    .B1(_02532_),
    .C1(_02537_),
    .X(_02698_));
 sky130_fd_sc_hd__a31oi_4 _25717_ (.A1(_02274_),
    .A2(_02279_),
    .A3(_02535_),
    .B1(_02696_),
    .Y(_02699_));
 sky130_fd_sc_hd__a31o_2 _25718_ (.A1(_02274_),
    .A2(_02279_),
    .A3(_02535_),
    .B1(_02696_),
    .X(_02700_));
 sky130_fd_sc_hd__nand2_2 _25719_ (.A(_02698_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__o21ai_2 _25720_ (.A1(_02697_),
    .A2(_02699_),
    .B1(_02159_),
    .Y(_02702_));
 sky130_fd_sc_hd__and3_2 _25721_ (.A(_02160_),
    .B(_02698_),
    .C(_02700_),
    .X(_02703_));
 sky130_fd_sc_hd__a211o_4 _25722_ (.A1(_01801_),
    .A2(_02157_),
    .B1(_02697_),
    .C1(_02699_),
    .X(_02704_));
 sky130_fd_sc_hd__and2_4 _25723_ (.A(_02702_),
    .B(_02704_),
    .X(_02706_));
 sky130_fd_sc_hd__o21ai_1 _25724_ (.A1(_00796_),
    .A2(_01324_),
    .B1(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__a21oi_4 _25725_ (.A1(_02702_),
    .A2(_02704_),
    .B1(_01332_),
    .Y(_02708_));
 sky130_fd_sc_hd__a211o_2 _25726_ (.A1(_02702_),
    .A2(_02704_),
    .B1(_00796_),
    .C1(_01324_),
    .X(_02709_));
 sky130_fd_sc_hd__a21oi_1 _25727_ (.A1(_02707_),
    .A2(_02709_),
    .B1(net131),
    .Y(_02710_));
 sky130_fd_sc_hd__o221a_4 _25728_ (.A1(_13066_),
    .A2(_00357_),
    .B1(_01332_),
    .B2(_02706_),
    .C1(_11740_),
    .X(_02711_));
 sky130_fd_sc_hd__or4_4 _25729_ (.A(_10544_),
    .B(_11735_),
    .C(_00360_),
    .D(_02708_),
    .X(_02712_));
 sky130_fd_sc_hd__a21oi_2 _25730_ (.A1(_02711_),
    .A2(_02707_),
    .B1(_02710_),
    .Y(_02713_));
 sky130_fd_sc_hd__xor2_4 _25731_ (.A(_02545_),
    .B(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__o21bai_1 _25732_ (.A1(_02691_),
    .A2(_02693_),
    .B1_N(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand3_1 _25733_ (.A(_02692_),
    .B(_02695_),
    .C(_02714_),
    .Y(_02717_));
 sky130_fd_sc_hd__o21ai_4 _25734_ (.A1(_02691_),
    .A2(_02693_),
    .B1(_02714_),
    .Y(_02718_));
 sky130_fd_sc_hd__a21oi_2 _25735_ (.A1(_02688_),
    .A2(_02690_),
    .B1(_02714_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand3b_4 _25736_ (.A_N(_02714_),
    .B(_02695_),
    .C(_02692_),
    .Y(_02720_));
 sky130_fd_sc_hd__nand2_2 _25737_ (.A(_02603_),
    .B(_02605_),
    .Y(_02721_));
 sky130_fd_sc_hd__a31oi_2 _25738_ (.A1(_02556_),
    .A2(_02557_),
    .A3(_02604_),
    .B1(_02602_),
    .Y(_02722_));
 sky130_fd_sc_hd__a21oi_4 _25739_ (.A1(_02718_),
    .A2(_02720_),
    .B1(_02721_),
    .Y(_02723_));
 sky130_fd_sc_hd__nand3_2 _25740_ (.A(_02715_),
    .B(_02717_),
    .C(_02722_),
    .Y(_02724_));
 sky130_fd_sc_hd__a21oi_1 _25741_ (.A1(_02715_),
    .A2(_02717_),
    .B1(_02722_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand3_4 _25742_ (.A(_02718_),
    .B(_02721_),
    .C(_02720_),
    .Y(_02726_));
 sky130_fd_sc_hd__nand2_2 _25743_ (.A(_02482_),
    .B(_02516_),
    .Y(_02728_));
 sky130_fd_sc_hd__a21oi_2 _25744_ (.A1(_02293_),
    .A2(_02550_),
    .B1(_02549_),
    .Y(_02729_));
 sky130_fd_sc_hd__a21boi_1 _25745_ (.A1(_02446_),
    .A2(_02473_),
    .B1_N(_02474_),
    .Y(_02730_));
 sky130_fd_sc_hd__nand2_1 _25746_ (.A(_02474_),
    .B(_02479_),
    .Y(_02731_));
 sky130_fd_sc_hd__and3_1 _25747_ (.A(_02328_),
    .B(_02335_),
    .C(_02466_),
    .X(_02732_));
 sky130_fd_sc_hd__o21ai_1 _25748_ (.A1(_02448_),
    .A2(_02452_),
    .B1(_02458_),
    .Y(_02733_));
 sky130_fd_sc_hd__nor2_2 _25749_ (.A(_04256_),
    .B(_06030_),
    .Y(_02734_));
 sky130_fd_sc_hd__o311a_1 _25750_ (.A1(_05931_),
    .A2(_07074_),
    .A3(net268),
    .B1(net274),
    .C1(net164),
    .X(_02735_));
 sky130_fd_sc_hd__a31oi_2 _25751_ (.A1(net164),
    .A2(_08208_),
    .A3(net274),
    .B1(_02734_),
    .Y(_02736_));
 sky130_fd_sc_hd__a21oi_2 _25752_ (.A1(net153),
    .A2(net158),
    .B1(_05763_),
    .Y(_02737_));
 sky130_fd_sc_hd__o21ai_1 _25753_ (.A1(_08664_),
    .A2(_08666_),
    .B1(_05762_),
    .Y(_02739_));
 sky130_fd_sc_hd__nor2_4 _25754_ (.A(net319),
    .B(_05766_),
    .Y(_02740_));
 sky130_fd_sc_hd__or3b_4 _25755_ (.A(net48),
    .B(net319),
    .C_N(net47),
    .X(_02741_));
 sky130_fd_sc_hd__o22a_2 _25756_ (.A1(_02734_),
    .A2(_02735_),
    .B1(_02737_),
    .B2(_02740_),
    .X(_02742_));
 sky130_fd_sc_hd__o22ai_4 _25757_ (.A1(_02734_),
    .A2(_02735_),
    .B1(_02737_),
    .B2(_02740_),
    .Y(_02743_));
 sky130_fd_sc_hd__o211ai_4 _25758_ (.A1(net319),
    .A2(_05766_),
    .B1(_02736_),
    .C1(_02739_),
    .Y(_02744_));
 sky130_fd_sc_hd__a32o_2 _25759_ (.A1(_07771_),
    .A2(net273),
    .A3(net166),
    .B1(_06326_),
    .B2(net22),
    .X(_02745_));
 sky130_fd_sc_hd__a21oi_1 _25760_ (.A1(_02743_),
    .A2(_02744_),
    .B1(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__a21o_2 _25761_ (.A1(_02743_),
    .A2(_02744_),
    .B1(_02745_),
    .X(_02747_));
 sky130_fd_sc_hd__and3_2 _25762_ (.A(_02743_),
    .B(_02744_),
    .C(_02745_),
    .X(_02748_));
 sky130_fd_sc_hd__nand3_4 _25763_ (.A(_02743_),
    .B(_02744_),
    .C(_02745_),
    .Y(_02750_));
 sky130_fd_sc_hd__o22ai_4 _25764_ (.A1(_02534_),
    .A2(_02536_),
    .B1(_02746_),
    .B2(_02748_),
    .Y(_02751_));
 sky130_fd_sc_hd__nand3_1 _25765_ (.A(_02747_),
    .B(_02750_),
    .C(_02539_),
    .Y(_02752_));
 sky130_fd_sc_hd__a21oi_1 _25766_ (.A1(_02751_),
    .A2(_02752_),
    .B1(_02733_),
    .Y(_02753_));
 sky130_fd_sc_hd__a21o_1 _25767_ (.A1(_02751_),
    .A2(_02752_),
    .B1(_02733_),
    .X(_02754_));
 sky130_fd_sc_hd__a32oi_4 _25768_ (.A1(_02747_),
    .A2(_02750_),
    .A3(_02539_),
    .B1(_02458_),
    .B2(_02454_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _25769_ (.A(_02755_),
    .B(_02751_),
    .Y(_02756_));
 sky130_fd_sc_hd__a211oi_2 _25770_ (.A1(_02751_),
    .A2(_02755_),
    .B1(_02544_),
    .C1(_02753_),
    .Y(_02757_));
 sky130_fd_sc_hd__a211o_2 _25771_ (.A1(_02751_),
    .A2(_02755_),
    .B1(_02544_),
    .C1(_02753_),
    .X(_02758_));
 sky130_fd_sc_hd__a21oi_2 _25772_ (.A1(_02754_),
    .A2(_02756_),
    .B1(_02543_),
    .Y(_02759_));
 sky130_fd_sc_hd__a21o_2 _25773_ (.A1(_02754_),
    .A2(_02756_),
    .B1(_02543_),
    .X(_02761_));
 sky130_fd_sc_hd__o22ai_2 _25774_ (.A1(_02465_),
    .A2(_02471_),
    .B1(_02757_),
    .B2(_02759_),
    .Y(_02762_));
 sky130_fd_sc_hd__o211ai_2 _25775_ (.A1(_02463_),
    .A2(_02732_),
    .B1(_02758_),
    .C1(_02761_),
    .Y(_02763_));
 sky130_fd_sc_hd__o22ai_4 _25776_ (.A1(_02463_),
    .A2(_02732_),
    .B1(_02757_),
    .B2(_02759_),
    .Y(_02764_));
 sky130_fd_sc_hd__o21ai_1 _25777_ (.A1(_02465_),
    .A2(_02471_),
    .B1(_02761_),
    .Y(_02765_));
 sky130_fd_sc_hd__o211ai_4 _25778_ (.A1(_02465_),
    .A2(_02471_),
    .B1(_02758_),
    .C1(_02761_),
    .Y(_02766_));
 sky130_fd_sc_hd__and3_1 _25779_ (.A(_02762_),
    .B(_02763_),
    .C(_02730_),
    .X(_02767_));
 sky130_fd_sc_hd__nand3_2 _25780_ (.A(_02762_),
    .B(_02763_),
    .C(_02730_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand3_4 _25781_ (.A(_02731_),
    .B(_02764_),
    .C(_02766_),
    .Y(_02769_));
 sky130_fd_sc_hd__inv_2 _25782_ (.A(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__a32oi_4 _25783_ (.A1(_06219_),
    .A2(_06221_),
    .A3(net238),
    .B1(_08006_),
    .B2(net17),
    .Y(_02772_));
 sky130_fd_sc_hd__a32o_1 _25784_ (.A1(_06219_),
    .A2(_06221_),
    .A3(net238),
    .B1(_08006_),
    .B2(net17),
    .X(_02773_));
 sky130_fd_sc_hd__a32o_1 _25785_ (.A1(_06449_),
    .A2(_06452_),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net18),
    .X(_02774_));
 sky130_fd_sc_hd__a32o_1 _25786_ (.A1(net192),
    .A2(_06762_),
    .A3(net239),
    .B1(_07308_),
    .B2(net19),
    .X(_02775_));
 sky130_fd_sc_hd__or3b_1 _25787_ (.A(net52),
    .B(_04212_),
    .C_N(net51),
    .X(_02776_));
 sky130_fd_sc_hd__o221ai_2 _25788_ (.A1(net176),
    .A2(_07074_),
    .B1(_04212_),
    .B2(net190),
    .C1(net269),
    .Y(_02777_));
 sky130_fd_sc_hd__nor2_1 _25789_ (.A(_04223_),
    .B(_06866_),
    .Y(_02778_));
 sky130_fd_sc_hd__a211oi_1 _25790_ (.A1(net204),
    .A2(_07500_),
    .B1(_06864_),
    .C1(_07498_),
    .Y(_02779_));
 sky130_fd_sc_hd__a31oi_1 _25791_ (.A1(_07499_),
    .A2(_07503_),
    .A3(net240),
    .B1(_02778_),
    .Y(_02780_));
 sky130_fd_sc_hd__o2bb2ai_1 _25792_ (.A1_N(_02776_),
    .A2_N(_02777_),
    .B1(_02778_),
    .B2(_02779_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand3_2 _25793_ (.A(_02780_),
    .B(_02777_),
    .C(_02776_),
    .Y(_02783_));
 sky130_fd_sc_hd__a21oi_2 _25794_ (.A1(_02781_),
    .A2(_02783_),
    .B1(_02775_),
    .Y(_02784_));
 sky130_fd_sc_hd__and3_1 _25795_ (.A(_02775_),
    .B(_02781_),
    .C(_02783_),
    .X(_02785_));
 sky130_fd_sc_hd__a211oi_1 _25796_ (.A1(_02495_),
    .A2(_02498_),
    .B1(_02784_),
    .C1(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__a211o_1 _25797_ (.A1(_02495_),
    .A2(_02498_),
    .B1(_02784_),
    .C1(_02785_),
    .X(_02787_));
 sky130_fd_sc_hd__o221ai_4 _25798_ (.A1(_02491_),
    .A2(_02494_),
    .B1(_02784_),
    .B2(_02785_),
    .C1(_02498_),
    .Y(_02788_));
 sky130_fd_sc_hd__a21o_1 _25799_ (.A1(_02787_),
    .A2(_02788_),
    .B1(_02774_),
    .X(_02789_));
 sky130_fd_sc_hd__nand3_2 _25800_ (.A(_02774_),
    .B(_02787_),
    .C(_02788_),
    .Y(_02790_));
 sky130_fd_sc_hd__and2_1 _25801_ (.A(_02789_),
    .B(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__a32o_1 _25802_ (.A1(_02487_),
    .A2(_02498_),
    .A3(_02499_),
    .B1(_02503_),
    .B2(_02485_),
    .X(_02792_));
 sky130_fd_sc_hd__a21oi_2 _25803_ (.A1(_02789_),
    .A2(_02790_),
    .B1(_02792_),
    .Y(_02794_));
 sky130_fd_sc_hd__and3_2 _25804_ (.A(_02789_),
    .B(_02790_),
    .C(_02792_),
    .X(_02795_));
 sky130_fd_sc_hd__nand2_1 _25805_ (.A(_02791_),
    .B(_02792_),
    .Y(_02796_));
 sky130_fd_sc_hd__nor3_1 _25806_ (.A(_02773_),
    .B(_02794_),
    .C(_02795_),
    .Y(_02797_));
 sky130_fd_sc_hd__o21a_1 _25807_ (.A1(_02794_),
    .A2(_02795_),
    .B1(_02773_),
    .X(_02798_));
 sky130_fd_sc_hd__nor3_1 _25808_ (.A(_02773_),
    .B(_02792_),
    .C(_02791_),
    .Y(_02799_));
 sky130_fd_sc_hd__nor3_4 _25809_ (.A(_02772_),
    .B(_02794_),
    .C(_02795_),
    .Y(_02800_));
 sky130_fd_sc_hd__a31o_1 _25810_ (.A1(_02789_),
    .A2(_02790_),
    .A3(_02792_),
    .B1(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__o21a_1 _25811_ (.A1(_02794_),
    .A2(_02795_),
    .B1(_02772_),
    .X(_02802_));
 sky130_fd_sc_hd__o21a_1 _25812_ (.A1(_02797_),
    .A2(_02798_),
    .B1(_02768_),
    .X(_02803_));
 sky130_fd_sc_hd__o211ai_2 _25813_ (.A1(_02797_),
    .A2(_02798_),
    .B1(_02768_),
    .C1(_02769_),
    .Y(_02805_));
 sky130_fd_sc_hd__o2bb2ai_2 _25814_ (.A1_N(_02768_),
    .A2_N(_02769_),
    .B1(_02800_),
    .B2(_02802_),
    .Y(_02806_));
 sky130_fd_sc_hd__o2bb2ai_1 _25815_ (.A1_N(_02768_),
    .A2_N(_02769_),
    .B1(_02797_),
    .B2(_02798_),
    .Y(_02807_));
 sky130_fd_sc_hd__o211ai_2 _25816_ (.A1(_02800_),
    .A2(_02802_),
    .B1(_02768_),
    .C1(_02769_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _25817_ (.A(_02805_),
    .B(_02806_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand3_4 _25818_ (.A(_02808_),
    .B(_02729_),
    .C(_02807_),
    .Y(_02810_));
 sky130_fd_sc_hd__o211ai_4 _25819_ (.A1(_02549_),
    .A2(_02555_),
    .B1(_02805_),
    .C1(_02806_),
    .Y(_02811_));
 sky130_fd_sc_hd__a21oi_2 _25820_ (.A1(_02810_),
    .A2(_02811_),
    .B1(_02728_),
    .Y(_02812_));
 sky130_fd_sc_hd__a21o_1 _25821_ (.A1(_02810_),
    .A2(_02811_),
    .B1(_02728_),
    .X(_02813_));
 sky130_fd_sc_hd__and3_1 _25822_ (.A(_02728_),
    .B(_02810_),
    .C(_02811_),
    .X(_02814_));
 sky130_fd_sc_hd__nand3_4 _25823_ (.A(_02728_),
    .B(_02810_),
    .C(_02811_),
    .Y(_02816_));
 sky130_fd_sc_hd__a22o_1 _25824_ (.A1(_02482_),
    .A2(_02516_),
    .B1(_02810_),
    .B2(_02811_),
    .X(_02817_));
 sky130_fd_sc_hd__nand4_1 _25825_ (.A(_02482_),
    .B(_02516_),
    .C(_02810_),
    .D(_02811_),
    .Y(_02818_));
 sky130_fd_sc_hd__o22a_1 _25826_ (.A1(_02723_),
    .A2(_02725_),
    .B1(_02812_),
    .B2(_02814_),
    .X(_02819_));
 sky130_fd_sc_hd__o2bb2ai_4 _25827_ (.A1_N(_02724_),
    .A2_N(_02726_),
    .B1(_02812_),
    .B2(_02814_),
    .Y(_02820_));
 sky130_fd_sc_hd__nand3_2 _25828_ (.A(_02726_),
    .B(_02813_),
    .C(_02816_),
    .Y(_02821_));
 sky130_fd_sc_hd__nand4_2 _25829_ (.A(_02724_),
    .B(_02726_),
    .C(_02813_),
    .D(_02816_),
    .Y(_02822_));
 sky130_fd_sc_hd__a22oi_4 _25830_ (.A1(_02613_),
    .A2(_02615_),
    .B1(_02820_),
    .B2(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__a31o_2 _25831_ (.A1(_02357_),
    .A2(_02397_),
    .A3(_02521_),
    .B1(_02522_),
    .X(_02824_));
 sky130_fd_sc_hd__o31a_1 _25832_ (.A1(_02356_),
    .A2(_02398_),
    .A3(_02520_),
    .B1(_02523_),
    .X(_02825_));
 sky130_fd_sc_hd__a211oi_2 _25833_ (.A1(_02820_),
    .A2(_02822_),
    .B1(_02825_),
    .C1(_02616_),
    .Y(_02827_));
 sky130_fd_sc_hd__o211ai_2 _25834_ (.A1(_02723_),
    .A2(_02821_),
    .B1(_02613_),
    .C1(_02615_),
    .Y(_02828_));
 sky130_fd_sc_hd__o2111a_1 _25835_ (.A1(_02723_),
    .A2(_02821_),
    .B1(_02820_),
    .C1(_02613_),
    .D1(_02615_),
    .X(_02829_));
 sky130_fd_sc_hd__o2111ai_4 _25836_ (.A1(_02723_),
    .A2(_02821_),
    .B1(_02820_),
    .C1(_02613_),
    .D1(_02615_),
    .Y(_02830_));
 sky130_fd_sc_hd__o22ai_4 _25837_ (.A1(_02819_),
    .A2(_02828_),
    .B1(_02824_),
    .B2(_02823_),
    .Y(_02831_));
 sky130_fd_sc_hd__nand3b_1 _25838_ (.A_N(_02823_),
    .B(_02825_),
    .C(_02830_),
    .Y(_02832_));
 sky130_fd_sc_hd__o21ai_1 _25839_ (.A1(_02823_),
    .A2(_02829_),
    .B1(_02824_),
    .Y(_02833_));
 sky130_fd_sc_hd__nand3_1 _25840_ (.A(_02644_),
    .B(_02832_),
    .C(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__o221ai_4 _25841_ (.A1(_02830_),
    .A2(_02824_),
    .B1(_02827_),
    .B2(_02831_),
    .C1(_02645_),
    .Y(_02835_));
 sky130_fd_sc_hd__a31o_1 _25842_ (.A1(_02644_),
    .A2(_02832_),
    .A3(_02833_),
    .B1(_02642_),
    .X(_02836_));
 sky130_fd_sc_hd__nand2_1 _25843_ (.A(_02834_),
    .B(_02835_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21oi_1 _25844_ (.A1(_02834_),
    .A2(_02835_),
    .B1(_02642_),
    .Y(_02839_));
 sky130_fd_sc_hd__and3_1 _25845_ (.A(_02834_),
    .B(_02835_),
    .C(_02642_),
    .X(_02840_));
 sky130_fd_sc_hd__o211ai_1 _25846_ (.A1(_02839_),
    .A2(_02840_),
    .B1(_02632_),
    .C1(_02634_),
    .Y(_02841_));
 sky130_fd_sc_hd__a21oi_1 _25847_ (.A1(_02632_),
    .A2(_02634_),
    .B1(_02839_),
    .Y(_02842_));
 sky130_fd_sc_hd__o21ai_1 _25848_ (.A1(_02643_),
    .A2(_02838_),
    .B1(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__nand2_1 _25849_ (.A(_02841_),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__and3b_1 _25850_ (.A_N(_02433_),
    .B(_02639_),
    .C(_02434_),
    .X(_02845_));
 sky130_fd_sc_hd__o21bai_1 _25851_ (.A1(_02434_),
    .A2(_02638_),
    .B1_N(_02637_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21oi_2 _25852_ (.A1(_02440_),
    .A2(_02845_),
    .B1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__xor2_1 _25853_ (.A(_02844_),
    .B(_02847_),
    .X(net114));
 sky130_fd_sc_hd__o21ai_1 _25854_ (.A1(_02729_),
    .A2(_02809_),
    .B1(_02816_),
    .Y(_02849_));
 sky130_fd_sc_hd__a2bb2o_1 _25855_ (.A1_N(_02545_),
    .A2_N(_02710_),
    .B1(_02711_),
    .B2(_02707_),
    .X(_02850_));
 sky130_fd_sc_hd__a311o_1 _25856_ (.A1(_02754_),
    .A2(_02756_),
    .A3(_02543_),
    .B1(_02471_),
    .C1(_02465_),
    .X(_02851_));
 sky130_fd_sc_hd__o31a_1 _25857_ (.A1(_02463_),
    .A2(_02732_),
    .A3(_02759_),
    .B1(_02758_),
    .X(_02852_));
 sky130_fd_sc_hd__a32oi_4 _25858_ (.A1(_02539_),
    .A2(_02747_),
    .A3(_02750_),
    .B1(_02755_),
    .B2(_02751_),
    .Y(_02853_));
 sky130_fd_sc_hd__a32o_1 _25859_ (.A1(_02539_),
    .A2(_02747_),
    .A3(_02750_),
    .B1(_02755_),
    .B2(_02751_),
    .X(_02854_));
 sky130_fd_sc_hd__a21o_1 _25860_ (.A1(_02744_),
    .A2(_02745_),
    .B1(_02742_),
    .X(_02855_));
 sky130_fd_sc_hd__o311a_1 _25861_ (.A1(net22),
    .A2(net24),
    .A3(_07503_),
    .B1(_05762_),
    .C1(net319),
    .X(_02856_));
 sky130_fd_sc_hd__a31oi_4 _25862_ (.A1(net319),
    .A2(net163),
    .A3(_05762_),
    .B1(_02740_),
    .Y(_02857_));
 sky130_fd_sc_hd__nor2_1 _25863_ (.A(net319),
    .B(_06030_),
    .Y(_02859_));
 sky130_fd_sc_hd__or3b_2 _25864_ (.A(net49),
    .B(net319),
    .C_N(net48),
    .X(_02860_));
 sky130_fd_sc_hd__a21oi_2 _25865_ (.A1(net153),
    .A2(net158),
    .B1(_06028_),
    .Y(_02861_));
 sky130_fd_sc_hd__o22a_1 _25866_ (.A1(net319),
    .A2(_06030_),
    .B1(_06028_),
    .B2(_08669_),
    .X(_02862_));
 sky130_fd_sc_hd__o221ai_4 _25867_ (.A1(net319),
    .A2(_06030_),
    .B1(_06028_),
    .B2(_08669_),
    .C1(_02857_),
    .Y(_02863_));
 sky130_fd_sc_hd__o22a_1 _25868_ (.A1(_02740_),
    .A2(_02856_),
    .B1(_02859_),
    .B2(_02861_),
    .X(_02864_));
 sky130_fd_sc_hd__o22ai_4 _25869_ (.A1(_02740_),
    .A2(_02856_),
    .B1(_02859_),
    .B2(_02861_),
    .Y(_02865_));
 sky130_fd_sc_hd__and3_1 _25870_ (.A(_04190_),
    .B(net24),
    .C(net49),
    .X(_02866_));
 sky130_fd_sc_hd__o311a_1 _25871_ (.A1(_05931_),
    .A2(_07074_),
    .A3(net268),
    .B1(net273),
    .C1(net164),
    .X(_02867_));
 sky130_fd_sc_hd__a31o_1 _25872_ (.A1(net164),
    .A2(net163),
    .A3(net273),
    .B1(_02866_),
    .X(_02868_));
 sky130_fd_sc_hd__a21oi_4 _25873_ (.A1(_02863_),
    .A2(_02865_),
    .B1(_02868_),
    .Y(_02870_));
 sky130_fd_sc_hd__o211a_1 _25874_ (.A1(_02866_),
    .A2(_02867_),
    .B1(_02863_),
    .C1(_02865_),
    .X(_02871_));
 sky130_fd_sc_hd__o211ai_4 _25875_ (.A1(_02866_),
    .A2(_02867_),
    .B1(_02863_),
    .C1(_02865_),
    .Y(_02872_));
 sky130_fd_sc_hd__a31o_2 _25876_ (.A1(_02863_),
    .A2(_02865_),
    .A3(_02868_),
    .B1(_02700_),
    .X(_02873_));
 sky130_fd_sc_hd__nor2_1 _25877_ (.A(_02870_),
    .B(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand3b_1 _25878_ (.A_N(_02870_),
    .B(_02872_),
    .C(_02699_),
    .Y(_02875_));
 sky130_fd_sc_hd__o22a_1 _25879_ (.A1(_02536_),
    .A2(_02696_),
    .B1(_02870_),
    .B2(_02871_),
    .X(_02876_));
 sky130_fd_sc_hd__o22ai_4 _25880_ (.A1(_02536_),
    .A2(_02696_),
    .B1(_02870_),
    .B2(_02871_),
    .Y(_02877_));
 sky130_fd_sc_hd__a21o_1 _25881_ (.A1(_02875_),
    .A2(_02877_),
    .B1(_02855_),
    .X(_02878_));
 sky130_fd_sc_hd__o21ai_4 _25882_ (.A1(_02742_),
    .A2(_02748_),
    .B1(_02877_),
    .Y(_02879_));
 sky130_fd_sc_hd__o22ai_2 _25883_ (.A1(_02742_),
    .A2(_02748_),
    .B1(_02874_),
    .B2(_02876_),
    .Y(_02881_));
 sky130_fd_sc_hd__o2111ai_4 _25884_ (.A1(_02873_),
    .A2(_02870_),
    .B1(_02750_),
    .C1(_02743_),
    .D1(_02877_),
    .Y(_02882_));
 sky130_fd_sc_hd__o211ai_4 _25885_ (.A1(_02701_),
    .A2(_02159_),
    .B1(_02882_),
    .C1(_02881_),
    .Y(_02883_));
 sky130_fd_sc_hd__o211ai_4 _25886_ (.A1(_02874_),
    .A2(_02879_),
    .B1(_02703_),
    .C1(_02878_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _25887_ (.A(_02883_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__a21oi_2 _25888_ (.A1(_02883_),
    .A2(_02884_),
    .B1(_02854_),
    .Y(_02886_));
 sky130_fd_sc_hd__a21o_1 _25889_ (.A1(_02883_),
    .A2(_02884_),
    .B1(_02854_),
    .X(_02887_));
 sky130_fd_sc_hd__a31o_1 _25890_ (.A1(_02704_),
    .A2(_02881_),
    .A3(_02882_),
    .B1(_02853_),
    .X(_02888_));
 sky130_fd_sc_hd__and3_1 _25891_ (.A(_02854_),
    .B(_02883_),
    .C(_02884_),
    .X(_02889_));
 sky130_fd_sc_hd__nand3_1 _25892_ (.A(_02854_),
    .B(_02883_),
    .C(_02884_),
    .Y(_02890_));
 sky130_fd_sc_hd__a22oi_2 _25893_ (.A1(_02885_),
    .A2(_02853_),
    .B1(_02765_),
    .B2(_02758_),
    .Y(_02892_));
 sky130_fd_sc_hd__a22oi_4 _25894_ (.A1(_02761_),
    .A2(_02851_),
    .B1(_02887_),
    .B2(_02890_),
    .Y(_02893_));
 sky130_fd_sc_hd__o21ai_1 _25895_ (.A1(_02886_),
    .A2(_02889_),
    .B1(_02852_),
    .Y(_02894_));
 sky130_fd_sc_hd__a32oi_2 _25896_ (.A1(_06449_),
    .A2(_06452_),
    .A3(net238),
    .B1(_08006_),
    .B2(net18),
    .Y(_02895_));
 sky130_fd_sc_hd__a32o_1 _25897_ (.A1(_06449_),
    .A2(_06452_),
    .A3(net238),
    .B1(_08006_),
    .B2(net18),
    .X(_02896_));
 sky130_fd_sc_hd__a32o_1 _25898_ (.A1(net192),
    .A2(_06762_),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net19),
    .X(_02897_));
 sky130_fd_sc_hd__a21boi_2 _25899_ (.A1(_02775_),
    .A2(_02783_),
    .B1_N(_02781_),
    .Y(_02898_));
 sky130_fd_sc_hd__a32o_1 _25900_ (.A1(_07072_),
    .A2(net170),
    .A3(net239),
    .B1(_07308_),
    .B2(net20),
    .X(_02899_));
 sky130_fd_sc_hd__or3b_1 _25901_ (.A(net52),
    .B(_04223_),
    .C_N(net51),
    .X(_02900_));
 sky130_fd_sc_hd__nand3_2 _25902_ (.A(_07499_),
    .B(_07503_),
    .C(net269),
    .Y(_02901_));
 sky130_fd_sc_hd__or3_2 _25903_ (.A(net51),
    .B(_04245_),
    .C(_04190_),
    .X(_02903_));
 sky130_fd_sc_hd__o211ai_2 _25904_ (.A1(net170),
    .A2(_07765_),
    .B1(net240),
    .C1(_07771_),
    .Y(_02904_));
 sky130_fd_sc_hd__a22oi_1 _25905_ (.A1(_02900_),
    .A2(_02901_),
    .B1(_02903_),
    .B2(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__a22o_1 _25906_ (.A1(_02900_),
    .A2(_02901_),
    .B1(_02903_),
    .B2(_02904_),
    .X(_02906_));
 sky130_fd_sc_hd__o2111a_1 _25907_ (.A1(_04223_),
    .A2(_07226_),
    .B1(_02901_),
    .C1(_02903_),
    .D1(_02904_),
    .X(_02907_));
 sky130_fd_sc_hd__o2111ai_2 _25908_ (.A1(_04223_),
    .A2(_07226_),
    .B1(_02901_),
    .C1(_02903_),
    .D1(_02904_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand3_1 _25909_ (.A(_02899_),
    .B(_02906_),
    .C(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__o21ai_1 _25910_ (.A1(_02905_),
    .A2(_02907_),
    .B1(_02899_),
    .Y(_02910_));
 sky130_fd_sc_hd__nand3b_1 _25911_ (.A_N(_02899_),
    .B(_02906_),
    .C(_02908_),
    .Y(_02911_));
 sky130_fd_sc_hd__nand3_1 _25912_ (.A(_02898_),
    .B(_02910_),
    .C(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__a21oi_1 _25913_ (.A1(_02910_),
    .A2(_02911_),
    .B1(_02898_),
    .Y(_02914_));
 sky130_fd_sc_hd__a21o_1 _25914_ (.A1(_02910_),
    .A2(_02911_),
    .B1(_02898_),
    .X(_02915_));
 sky130_fd_sc_hd__a21bo_1 _25915_ (.A1(_02912_),
    .A2(_02915_),
    .B1_N(_02897_),
    .X(_02916_));
 sky130_fd_sc_hd__nand3b_2 _25916_ (.A_N(_02897_),
    .B(_02912_),
    .C(_02915_),
    .Y(_02917_));
 sky130_fd_sc_hd__a21oi_2 _25917_ (.A1(_02774_),
    .A2(_02788_),
    .B1(_02786_),
    .Y(_02918_));
 sky130_fd_sc_hd__and3_1 _25918_ (.A(_02916_),
    .B(_02917_),
    .C(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__nand2_1 _25919_ (.A(_02895_),
    .B(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__a21oi_4 _25920_ (.A1(_02916_),
    .A2(_02917_),
    .B1(_02918_),
    .Y(_02921_));
 sky130_fd_sc_hd__a31oi_2 _25921_ (.A1(_02916_),
    .A2(_02917_),
    .A3(_02918_),
    .B1(_02895_),
    .Y(_02922_));
 sky130_fd_sc_hd__nor2_4 _25922_ (.A(_02921_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__a22oi_4 _25923_ (.A1(_02896_),
    .A2(_02921_),
    .B1(_02923_),
    .B2(_02920_),
    .Y(_02925_));
 sky130_fd_sc_hd__a22o_1 _25924_ (.A1(_02896_),
    .A2(_02921_),
    .B1(_02923_),
    .B2(_02920_),
    .X(_02926_));
 sky130_fd_sc_hd__o21ai_1 _25925_ (.A1(_02892_),
    .A2(_02893_),
    .B1(_02925_),
    .Y(_02927_));
 sky130_fd_sc_hd__o21ai_1 _25926_ (.A1(_02852_),
    .A2(_02886_),
    .B1(_02926_),
    .Y(_02928_));
 sky130_fd_sc_hd__o21ai_1 _25927_ (.A1(_02892_),
    .A2(_02893_),
    .B1(_02926_),
    .Y(_02929_));
 sky130_fd_sc_hd__o211ai_2 _25928_ (.A1(_02852_),
    .A2(_02886_),
    .B1(_02925_),
    .C1(_02894_),
    .Y(_02930_));
 sky130_fd_sc_hd__nand3b_4 _25929_ (.A_N(_02850_),
    .B(_02929_),
    .C(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__inv_2 _25930_ (.A(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__o211ai_4 _25931_ (.A1(_02893_),
    .A2(_02928_),
    .B1(_02927_),
    .C1(_02850_),
    .Y(_02933_));
 sky130_fd_sc_hd__o221a_1 _25932_ (.A1(_02772_),
    .A2(_02796_),
    .B1(_02799_),
    .B2(_02801_),
    .C1(_02769_),
    .X(_02934_));
 sky130_fd_sc_hd__a31o_1 _25933_ (.A1(_02731_),
    .A2(_02764_),
    .A3(_02766_),
    .B1(_02803_),
    .X(_02936_));
 sky130_fd_sc_hd__o211a_1 _25934_ (.A1(_02770_),
    .A2(_02803_),
    .B1(_02931_),
    .C1(_02933_),
    .X(_02937_));
 sky130_fd_sc_hd__o211ai_1 _25935_ (.A1(_02770_),
    .A2(_02803_),
    .B1(_02931_),
    .C1(_02933_),
    .Y(_02938_));
 sky130_fd_sc_hd__a21oi_1 _25936_ (.A1(_02931_),
    .A2(_02933_),
    .B1(_02936_),
    .Y(_02939_));
 sky130_fd_sc_hd__o2bb2ai_1 _25937_ (.A1_N(_02931_),
    .A2_N(_02933_),
    .B1(_02934_),
    .B2(_02767_),
    .Y(_02940_));
 sky130_fd_sc_hd__a2bb2o_1 _25938_ (.A1_N(_02770_),
    .A2_N(_02803_),
    .B1(_02931_),
    .B2(_02933_),
    .X(_02941_));
 sky130_fd_sc_hd__o211ai_1 _25939_ (.A1(_02767_),
    .A2(_02934_),
    .B1(_02933_),
    .C1(_02931_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2_1 _25940_ (.A(_02938_),
    .B(_02940_),
    .Y(_02943_));
 sky130_fd_sc_hd__a31o_4 _25941_ (.A1(_00361_),
    .A2(_10542_),
    .A3(_11736_),
    .B1(_01332_),
    .X(_02944_));
 sky130_fd_sc_hd__o31a_4 _25942_ (.A1(_10544_),
    .A2(_11735_),
    .A3(_00360_),
    .B1(_02708_),
    .X(_02945_));
 sky130_fd_sc_hd__a31o_2 _25943_ (.A1(_00361_),
    .A2(_10542_),
    .A3(_11736_),
    .B1(_02709_),
    .X(_02947_));
 sky130_fd_sc_hd__o21a_2 _25944_ (.A1(_02706_),
    .A2(_02944_),
    .B1(_02712_),
    .X(_02948_));
 sky130_fd_sc_hd__o21ai_4 _25945_ (.A1(_02706_),
    .A2(_02944_),
    .B1(_02712_),
    .Y(_02949_));
 sky130_fd_sc_hd__a21oi_2 _25946_ (.A1(_02681_),
    .A2(_00736_),
    .B1(_02682_),
    .Y(_02950_));
 sky130_fd_sc_hd__a2bb2oi_1 _25947_ (.A1_N(_02669_),
    .A2_N(_02664_),
    .B1(_12099_),
    .B2(_02671_),
    .Y(_02951_));
 sky130_fd_sc_hd__a2bb2o_2 _25948_ (.A1_N(_02664_),
    .A2_N(_02669_),
    .B1(_02671_),
    .B2(_12099_),
    .X(_02952_));
 sky130_fd_sc_hd__a21oi_1 _25949_ (.A1(_02653_),
    .A2(net157),
    .B1(net144),
    .Y(_02953_));
 sky130_fd_sc_hd__a31o_2 _25950_ (.A1(_02653_),
    .A2(_08664_),
    .A3(net33),
    .B1(net144),
    .X(_02954_));
 sky130_fd_sc_hd__nor2_1 _25951_ (.A(_04168_),
    .B(_08660_),
    .Y(_02955_));
 sky130_fd_sc_hd__a31oi_2 _25952_ (.A1(_06219_),
    .A2(_06221_),
    .A3(_08657_),
    .B1(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__a31o_1 _25953_ (.A1(_06219_),
    .A2(_06221_),
    .A3(_08657_),
    .B1(_02955_),
    .X(_02958_));
 sky130_fd_sc_hd__o21ai_4 _25954_ (.A1(_03286_),
    .A2(net152),
    .B1(_02956_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand3_4 _25955_ (.A(_02958_),
    .B(_08664_),
    .C(net33),
    .Y(_02960_));
 sky130_fd_sc_hd__a21oi_4 _25956_ (.A1(_02959_),
    .A2(_02960_),
    .B1(net144),
    .Y(_02961_));
 sky130_fd_sc_hd__a21o_1 _25957_ (.A1(_02959_),
    .A2(_02960_),
    .B1(net144),
    .X(_02962_));
 sky130_fd_sc_hd__o211a_1 _25958_ (.A1(net237),
    .A2(_09297_),
    .B1(_02959_),
    .C1(_02960_),
    .X(_02963_));
 sky130_fd_sc_hd__o211ai_4 _25959_ (.A1(net237),
    .A2(_09297_),
    .B1(_02959_),
    .C1(_02960_),
    .Y(_02964_));
 sky130_fd_sc_hd__o211ai_4 _25960_ (.A1(_02653_),
    .A2(net157),
    .B1(_02964_),
    .C1(_02954_),
    .Y(_02965_));
 sky130_fd_sc_hd__o2111ai_4 _25961_ (.A1(net157),
    .A2(_02653_),
    .B1(_02954_),
    .C1(_02962_),
    .D1(_02964_),
    .Y(_02966_));
 sky130_fd_sc_hd__a22oi_4 _25962_ (.A1(_02657_),
    .A2(_02954_),
    .B1(_02962_),
    .B2(_02964_),
    .Y(_02967_));
 sky130_fd_sc_hd__o22ai_4 _25963_ (.A1(_02656_),
    .A2(_02953_),
    .B1(_02961_),
    .B2(_02963_),
    .Y(_02969_));
 sky130_fd_sc_hd__a21oi_2 _25964_ (.A1(_02966_),
    .A2(_02969_),
    .B1(_10545_),
    .Y(_02970_));
 sky130_fd_sc_hd__a22o_1 _25965_ (.A1(net139),
    .A2(_10544_),
    .B1(_02966_),
    .B2(_02969_),
    .X(_02971_));
 sky130_fd_sc_hd__nand2_1 _25966_ (.A(_02969_),
    .B(_10545_),
    .Y(_02972_));
 sky130_fd_sc_hd__o211ai_2 _25967_ (.A1(_02961_),
    .A2(_02965_),
    .B1(_10545_),
    .C1(_02969_),
    .Y(_02973_));
 sky130_fd_sc_hd__o221ai_4 _25968_ (.A1(net140),
    .A2(_10542_),
    .B1(_02961_),
    .B2(_02965_),
    .C1(_02969_),
    .Y(_02974_));
 sky130_fd_sc_hd__a21o_1 _25969_ (.A1(_02966_),
    .A2(_02969_),
    .B1(_10546_),
    .X(_02975_));
 sky130_fd_sc_hd__a32oi_4 _25970_ (.A1(_02649_),
    .A2(_02658_),
    .A3(_02659_),
    .B1(_02662_),
    .B2(_10546_),
    .Y(_02976_));
 sky130_fd_sc_hd__a32o_1 _25971_ (.A1(_02649_),
    .A2(_02658_),
    .A3(_02659_),
    .B1(_02662_),
    .B2(_10546_),
    .X(_02977_));
 sky130_fd_sc_hd__nand3_4 _25972_ (.A(_02974_),
    .B(_02975_),
    .C(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__nand2_2 _25973_ (.A(_02976_),
    .B(_02973_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand3_1 _25974_ (.A(_02971_),
    .B(_02973_),
    .C(_02976_),
    .Y(_02981_));
 sky130_fd_sc_hd__o221a_1 _25975_ (.A1(net141),
    .A2(_11742_),
    .B1(_02970_),
    .B2(_02980_),
    .C1(_02978_),
    .X(_02982_));
 sky130_fd_sc_hd__o221ai_4 _25976_ (.A1(net141),
    .A2(_11742_),
    .B1(_02970_),
    .B2(_02980_),
    .C1(_02978_),
    .Y(_02983_));
 sky130_fd_sc_hd__a21oi_1 _25977_ (.A1(_02978_),
    .A2(_02981_),
    .B1(_12099_),
    .Y(_02984_));
 sky130_fd_sc_hd__a21o_1 _25978_ (.A1(_02978_),
    .A2(_02981_),
    .B1(_12099_),
    .X(_02985_));
 sky130_fd_sc_hd__nor3_2 _25979_ (.A(_02951_),
    .B(_02982_),
    .C(_02984_),
    .Y(_02986_));
 sky130_fd_sc_hd__nand3_4 _25980_ (.A(_02952_),
    .B(_02983_),
    .C(_02985_),
    .Y(_02987_));
 sky130_fd_sc_hd__a21oi_4 _25981_ (.A1(_02983_),
    .A2(_02985_),
    .B1(_02952_),
    .Y(_02988_));
 sky130_fd_sc_hd__o21ai_2 _25982_ (.A1(_02982_),
    .A2(_02984_),
    .B1(_02951_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand2_1 _25983_ (.A(_02989_),
    .B(_00736_),
    .Y(_02991_));
 sky130_fd_sc_hd__o2111ai_4 _25984_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_02987_),
    .D1(_02989_),
    .Y(_02992_));
 sky130_fd_sc_hd__o22ai_4 _25985_ (.A1(net131),
    .A2(_00366_),
    .B1(_02986_),
    .B2(_02988_),
    .Y(_02993_));
 sky130_fd_sc_hd__o211ai_2 _25986_ (.A1(net131),
    .A2(_00366_),
    .B1(_02987_),
    .C1(_02989_),
    .Y(_02994_));
 sky130_fd_sc_hd__o21ai_2 _25987_ (.A1(_02986_),
    .A2(_02988_),
    .B1(_00736_),
    .Y(_02995_));
 sky130_fd_sc_hd__o211a_1 _25988_ (.A1(_02682_),
    .A2(_02686_),
    .B1(_02992_),
    .C1(_02993_),
    .X(_02996_));
 sky130_fd_sc_hd__o211ai_4 _25989_ (.A1(_02682_),
    .A2(_02686_),
    .B1(_02992_),
    .C1(_02993_),
    .Y(_02997_));
 sky130_fd_sc_hd__a21boi_4 _25990_ (.A1(_02992_),
    .A2(_02993_),
    .B1_N(_02950_),
    .Y(_02998_));
 sky130_fd_sc_hd__a31oi_1 _25991_ (.A1(_02995_),
    .A2(_02950_),
    .A3(_02994_),
    .B1(_02949_),
    .Y(_02999_));
 sky130_fd_sc_hd__nand2_2 _25992_ (.A(_02999_),
    .B(_02997_),
    .Y(_03000_));
 sky130_fd_sc_hd__o22ai_4 _25993_ (.A1(_02711_),
    .A2(_02945_),
    .B1(_02996_),
    .B2(_02998_),
    .Y(_03002_));
 sky130_fd_sc_hd__o21ai_2 _25994_ (.A1(_02714_),
    .A2(_02691_),
    .B1(_02695_),
    .Y(_03003_));
 sky130_fd_sc_hd__o211a_1 _25995_ (.A1(_02693_),
    .A2(_02719_),
    .B1(_03000_),
    .C1(_03002_),
    .X(_03004_));
 sky130_fd_sc_hd__o211ai_4 _25996_ (.A1(_02693_),
    .A2(_02719_),
    .B1(_03000_),
    .C1(_03002_),
    .Y(_03005_));
 sky130_fd_sc_hd__a21oi_4 _25997_ (.A1(_03000_),
    .A2(_03002_),
    .B1(_03003_),
    .Y(_03006_));
 sky130_fd_sc_hd__a21o_1 _25998_ (.A1(_03000_),
    .A2(_03002_),
    .B1(_03003_),
    .X(_03007_));
 sky130_fd_sc_hd__o2bb2ai_1 _25999_ (.A1_N(_02941_),
    .A2_N(_02942_),
    .B1(_03004_),
    .B2(_03006_),
    .Y(_03008_));
 sky130_fd_sc_hd__o211ai_2 _26000_ (.A1(_02937_),
    .A2(_02939_),
    .B1(_03005_),
    .C1(_03007_),
    .Y(_03009_));
 sky130_fd_sc_hd__o22ai_2 _26001_ (.A1(_02937_),
    .A2(_02939_),
    .B1(_03004_),
    .B2(_03006_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand3_1 _26002_ (.A(_02938_),
    .B(_02940_),
    .C(_03005_),
    .Y(_03011_));
 sky130_fd_sc_hd__a31oi_2 _26003_ (.A1(_02726_),
    .A2(_02817_),
    .A3(_02818_),
    .B1(_02723_),
    .Y(_03013_));
 sky130_fd_sc_hd__a31oi_2 _26004_ (.A1(_02724_),
    .A2(_02813_),
    .A3(_02816_),
    .B1(_02725_),
    .Y(_03014_));
 sky130_fd_sc_hd__o211ai_4 _26005_ (.A1(_03006_),
    .A2(_03011_),
    .B1(_03013_),
    .C1(_03010_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand3_4 _26006_ (.A(_03008_),
    .B(_03009_),
    .C(_03014_),
    .Y(_03016_));
 sky130_fd_sc_hd__nand3_1 _26007_ (.A(_03016_),
    .B(_02849_),
    .C(_03015_),
    .Y(_03017_));
 sky130_fd_sc_hd__a21o_1 _26008_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_02849_),
    .X(_03018_));
 sky130_fd_sc_hd__a22o_1 _26009_ (.A1(_02811_),
    .A2(_02816_),
    .B1(_03015_),
    .B2(_03016_),
    .X(_03019_));
 sky130_fd_sc_hd__nand4_1 _26010_ (.A(_02811_),
    .B(_02816_),
    .C(_03015_),
    .D(_03016_),
    .Y(_03020_));
 sky130_fd_sc_hd__nand3b_2 _26011_ (.A_N(_02831_),
    .B(_03019_),
    .C(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__nand3_4 _26012_ (.A(_03018_),
    .B(_02831_),
    .C(_03017_),
    .Y(_03022_));
 sky130_fd_sc_hd__a21oi_1 _26013_ (.A1(_03021_),
    .A2(_03022_),
    .B1(_02801_),
    .Y(_03024_));
 sky130_fd_sc_hd__a21o_1 _26014_ (.A1(_03021_),
    .A2(_03022_),
    .B1(_02801_),
    .X(_03025_));
 sky130_fd_sc_hd__and3_1 _26015_ (.A(_03021_),
    .B(_03022_),
    .C(_02801_),
    .X(_03026_));
 sky130_fd_sc_hd__o211ai_4 _26016_ (.A1(_02795_),
    .A2(_02800_),
    .B1(_03021_),
    .C1(_03022_),
    .Y(_03027_));
 sky130_fd_sc_hd__o2bb2a_1 _26017_ (.A1_N(_02835_),
    .A2_N(_02836_),
    .B1(_03024_),
    .B2(_03026_),
    .X(_03028_));
 sky130_fd_sc_hd__o2bb2ai_1 _26018_ (.A1_N(_02835_),
    .A2_N(_02836_),
    .B1(_03024_),
    .B2(_03026_),
    .Y(_03029_));
 sky130_fd_sc_hd__nand4_1 _26019_ (.A(_02835_),
    .B(_02836_),
    .C(_03025_),
    .D(_03027_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand2_1 _26020_ (.A(_03029_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__o21ai_1 _26021_ (.A1(_02844_),
    .A2(_02847_),
    .B1(_02843_),
    .Y(_03032_));
 sky130_fd_sc_hd__xnor2_1 _26022_ (.A(_03031_),
    .B(_03032_),
    .Y(net115));
 sky130_fd_sc_hd__nand2_1 _26023_ (.A(_03022_),
    .B(_03027_),
    .Y(_03034_));
 sky130_fd_sc_hd__o211ai_2 _26024_ (.A1(_02729_),
    .A2(_02809_),
    .B1(_02816_),
    .C1(_03015_),
    .Y(_03035_));
 sky130_fd_sc_hd__a21bo_1 _26025_ (.A1(_02849_),
    .A2(_03016_),
    .B1_N(_03015_),
    .X(_03036_));
 sky130_fd_sc_hd__a31oi_1 _26026_ (.A1(_02941_),
    .A2(_02942_),
    .A3(_03005_),
    .B1(_03006_),
    .Y(_03037_));
 sky130_fd_sc_hd__and3_2 _26027_ (.A(_04190_),
    .B(net25),
    .C(net49),
    .X(_03038_));
 sky130_fd_sc_hd__or3b_1 _26028_ (.A(net50),
    .B(net319),
    .C_N(net49),
    .X(_03039_));
 sky130_fd_sc_hd__a21oi_2 _26029_ (.A1(net153),
    .A2(net158),
    .B1(_06325_),
    .Y(_03040_));
 sky130_fd_sc_hd__o211ai_4 _26030_ (.A1(_07076_),
    .A2(net268),
    .B1(net319),
    .C1(net274),
    .Y(_03041_));
 sky130_fd_sc_hd__o2111a_1 _26031_ (.A1(_05763_),
    .A2(net153),
    .B1(_02741_),
    .C1(_02860_),
    .D1(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__o2111ai_4 _26032_ (.A1(_05763_),
    .A2(net153),
    .B1(_02741_),
    .C1(_02860_),
    .D1(_03041_),
    .Y(_03043_));
 sky130_fd_sc_hd__o211ai_2 _26033_ (.A1(_06325_),
    .A2(_08669_),
    .B1(_03039_),
    .C1(_03042_),
    .Y(_03045_));
 sky130_fd_sc_hd__o21ai_2 _26034_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_03043_),
    .Y(_03046_));
 sky130_fd_sc_hd__nand3_1 _26035_ (.A(_03045_),
    .B(_03046_),
    .C(_02699_),
    .Y(_03047_));
 sky130_fd_sc_hd__a2bb2o_1 _26036_ (.A1_N(_02536_),
    .A2_N(_02696_),
    .B1(_03045_),
    .B2(_03046_),
    .X(_03048_));
 sky130_fd_sc_hd__a21o_1 _26037_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_02700_),
    .X(_03049_));
 sky130_fd_sc_hd__o211ai_2 _26038_ (.A1(_02536_),
    .A2(_02696_),
    .B1(_03045_),
    .C1(_03046_),
    .Y(_03050_));
 sky130_fd_sc_hd__a22o_1 _26039_ (.A1(_02865_),
    .A2(_02872_),
    .B1(_03049_),
    .B2(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__o2111ai_1 _26040_ (.A1(_02857_),
    .A2(_02862_),
    .B1(_02872_),
    .C1(_03049_),
    .D1(_03050_),
    .Y(_03052_));
 sky130_fd_sc_hd__o2111ai_4 _26041_ (.A1(_02857_),
    .A2(_02862_),
    .B1(_02872_),
    .C1(_03047_),
    .D1(_03048_),
    .Y(_03053_));
 sky130_fd_sc_hd__o211ai_2 _26042_ (.A1(_02864_),
    .A2(_02871_),
    .B1(_03049_),
    .C1(_03050_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand3_2 _26043_ (.A(_03051_),
    .B(_03052_),
    .C(_02703_),
    .Y(_03056_));
 sky130_fd_sc_hd__o211ai_4 _26044_ (.A1(_02701_),
    .A2(_02159_),
    .B1(_03054_),
    .C1(_03053_),
    .Y(_03057_));
 sky130_fd_sc_hd__and2_1 _26045_ (.A(_03056_),
    .B(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__a2bb2o_1 _26046_ (.A1_N(_02873_),
    .A2_N(_02870_),
    .B1(_02855_),
    .B2(_02877_),
    .X(_03059_));
 sky130_fd_sc_hd__a22o_1 _26047_ (.A1(_02875_),
    .A2(_02879_),
    .B1(_03056_),
    .B2(_03057_),
    .X(_03060_));
 sky130_fd_sc_hd__o2111ai_4 _26048_ (.A1(_02870_),
    .A2(_02873_),
    .B1(_02879_),
    .C1(_03056_),
    .D1(_03057_),
    .Y(_03061_));
 sky130_fd_sc_hd__a32o_1 _26049_ (.A1(_02704_),
    .A2(_03053_),
    .A3(_03054_),
    .B1(_02875_),
    .B2(_02879_),
    .X(_03062_));
 sky130_fd_sc_hd__o2bb2ai_2 _26050_ (.A1_N(_02884_),
    .A2_N(_02888_),
    .B1(_03058_),
    .B2(_03059_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand4_4 _26051_ (.A(_02884_),
    .B(_02888_),
    .C(_03060_),
    .D(_03061_),
    .Y(_03064_));
 sky130_fd_sc_hd__o2bb2a_1 _26052_ (.A1_N(_06763_),
    .A2_N(net238),
    .B1(_08007_),
    .B2(_04201_),
    .X(_03065_));
 sky130_fd_sc_hd__and3b_1 _26053_ (.A_N(net54),
    .B(net53),
    .C(net20),
    .X(_03067_));
 sky130_fd_sc_hd__o311a_1 _26054_ (.A1(net244),
    .A2(net241),
    .A3(_07074_),
    .B1(_07642_),
    .C1(_07072_),
    .X(_03068_));
 sky130_fd_sc_hd__a21oi_1 _26055_ (.A1(_07077_),
    .A2(_07642_),
    .B1(_03067_),
    .Y(_03069_));
 sky130_fd_sc_hd__a21o_1 _26056_ (.A1(_02899_),
    .A2(_02908_),
    .B1(_02905_),
    .X(_03070_));
 sky130_fd_sc_hd__o2bb2a_1 _26057_ (.A1_N(net21),
    .A2_N(_07308_),
    .B1(_07506_),
    .B2(_07306_),
    .X(_03071_));
 sky130_fd_sc_hd__a32o_1 _26058_ (.A1(_07499_),
    .A2(_07503_),
    .A3(net239),
    .B1(_07308_),
    .B2(net21),
    .X(_03072_));
 sky130_fd_sc_hd__or3b_2 _26059_ (.A(net52),
    .B(_04245_),
    .C_N(net51),
    .X(_03073_));
 sky130_fd_sc_hd__o211ai_4 _26060_ (.A1(net170),
    .A2(_07765_),
    .B1(net269),
    .C1(_07771_),
    .Y(_03074_));
 sky130_fd_sc_hd__or3_2 _26061_ (.A(net51),
    .B(_04256_),
    .C(_04190_),
    .X(_03075_));
 sky130_fd_sc_hd__o211ai_4 _26062_ (.A1(net170),
    .A2(net268),
    .B1(net240),
    .C1(_08204_),
    .Y(_03076_));
 sky130_fd_sc_hd__a22oi_4 _26063_ (.A1(_03073_),
    .A2(_03074_),
    .B1(_03075_),
    .B2(_03076_),
    .Y(_03078_));
 sky130_fd_sc_hd__a22o_1 _26064_ (.A1(_03073_),
    .A2(_03074_),
    .B1(_03075_),
    .B2(_03076_),
    .X(_03079_));
 sky130_fd_sc_hd__o2111a_1 _26065_ (.A1(_04245_),
    .A2(_07226_),
    .B1(_03074_),
    .C1(_03075_),
    .D1(_03076_),
    .X(_03080_));
 sky130_fd_sc_hd__o2111ai_2 _26066_ (.A1(_04245_),
    .A2(_07226_),
    .B1(_03074_),
    .C1(_03075_),
    .D1(_03076_),
    .Y(_03081_));
 sky130_fd_sc_hd__o21ai_2 _26067_ (.A1(_03078_),
    .A2(_03080_),
    .B1(_03071_),
    .Y(_03082_));
 sky130_fd_sc_hd__nor3_1 _26068_ (.A(_03071_),
    .B(_03078_),
    .C(_03080_),
    .Y(_03083_));
 sky130_fd_sc_hd__nand3_2 _26069_ (.A(_03072_),
    .B(_03079_),
    .C(_03081_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand3_2 _26070_ (.A(_03070_),
    .B(_03082_),
    .C(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__a21o_1 _26071_ (.A1(_03082_),
    .A2(_03084_),
    .B1(_03070_),
    .X(_03086_));
 sky130_fd_sc_hd__a22o_1 _26072_ (.A1(_02906_),
    .A2(_02909_),
    .B1(_03082_),
    .B2(_03084_),
    .X(_03087_));
 sky130_fd_sc_hd__nand4_1 _26073_ (.A(_02906_),
    .B(_02909_),
    .C(_03082_),
    .D(_03084_),
    .Y(_03089_));
 sky130_fd_sc_hd__o211ai_4 _26074_ (.A1(_03067_),
    .A2(_03068_),
    .B1(_03085_),
    .C1(_03086_),
    .Y(_03090_));
 sky130_fd_sc_hd__nand3_2 _26075_ (.A(_03087_),
    .B(_03089_),
    .C(_03069_),
    .Y(_03091_));
 sky130_fd_sc_hd__a21oi_1 _26076_ (.A1(_02897_),
    .A2(_02912_),
    .B1(_02914_),
    .Y(_03092_));
 sky130_fd_sc_hd__nand3b_4 _26077_ (.A_N(_03092_),
    .B(_03091_),
    .C(_03090_),
    .Y(_03093_));
 sky130_fd_sc_hd__a21bo_1 _26078_ (.A1(_03090_),
    .A2(_03091_),
    .B1_N(_03092_),
    .X(_03094_));
 sky130_fd_sc_hd__nand3b_2 _26079_ (.A_N(_03065_),
    .B(_03093_),
    .C(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a21bo_1 _26080_ (.A1(_03093_),
    .A2(_03094_),
    .B1_N(_03065_),
    .X(_03096_));
 sky130_fd_sc_hd__nand2_1 _26081_ (.A(_03095_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__a21o_1 _26082_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__nand3_1 _26083_ (.A(_03063_),
    .B(_03064_),
    .C(_03097_),
    .Y(_03100_));
 sky130_fd_sc_hd__a22o_1 _26084_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_03095_),
    .B2(_03096_),
    .X(_03101_));
 sky130_fd_sc_hd__nand4_1 _26085_ (.A(_03063_),
    .B(_03064_),
    .C(_03095_),
    .D(_03096_),
    .Y(_03102_));
 sky130_fd_sc_hd__o211ai_2 _26086_ (.A1(_02708_),
    .A2(_00364_),
    .B1(_03100_),
    .C1(_03098_),
    .Y(_03103_));
 sky130_fd_sc_hd__o2111ai_4 _26087_ (.A1(_01332_),
    .A2(_02706_),
    .B1(_03102_),
    .C1(net131),
    .D1(_03101_),
    .Y(_03104_));
 sky130_fd_sc_hd__a32o_1 _26088_ (.A1(_02761_),
    .A2(_02851_),
    .A3(_02887_),
    .B1(_02894_),
    .B2(_02926_),
    .X(_03105_));
 sky130_fd_sc_hd__o22a_1 _26089_ (.A1(_02886_),
    .A2(_02852_),
    .B1(_02925_),
    .B2(_02893_),
    .X(_03106_));
 sky130_fd_sc_hd__a21o_1 _26090_ (.A1(_03103_),
    .A2(_03104_),
    .B1(_03105_),
    .X(_03107_));
 sky130_fd_sc_hd__nand3_1 _26091_ (.A(_03103_),
    .B(_03104_),
    .C(_03105_),
    .Y(_03108_));
 sky130_fd_sc_hd__a21o_1 _26092_ (.A1(_03103_),
    .A2(_03104_),
    .B1(_03106_),
    .X(_03109_));
 sky130_fd_sc_hd__nand3_1 _26093_ (.A(_03103_),
    .B(_03104_),
    .C(_03106_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _26094_ (.A(_03107_),
    .B(_03108_),
    .Y(_03112_));
 sky130_fd_sc_hd__a21boi_2 _26095_ (.A1(_12099_),
    .A2(_02978_),
    .B1_N(_02981_),
    .Y(_03113_));
 sky130_fd_sc_hd__o2bb2ai_2 _26096_ (.A1_N(_12099_),
    .A2_N(_02978_),
    .B1(_02980_),
    .B2(_02970_),
    .Y(_03114_));
 sky130_fd_sc_hd__o22a_1 _26097_ (.A1(net140),
    .A2(_10542_),
    .B1(_02961_),
    .B2(_02965_),
    .X(_03115_));
 sky130_fd_sc_hd__o22ai_4 _26098_ (.A1(_02961_),
    .A2(_02965_),
    .B1(_10546_),
    .B2(_02967_),
    .Y(_03116_));
 sky130_fd_sc_hd__a21boi_4 _26099_ (.A1(net144),
    .A2(_02959_),
    .B1_N(_02960_),
    .Y(_03117_));
 sky130_fd_sc_hd__o21ai_1 _26100_ (.A1(net149),
    .A2(_02956_),
    .B1(_02964_),
    .Y(_03118_));
 sky130_fd_sc_hd__or3_1 _26101_ (.A(net57),
    .B(_04266_),
    .C(_04179_),
    .X(_03119_));
 sky130_fd_sc_hd__nand3_4 _26102_ (.A(_06449_),
    .B(_06452_),
    .C(_08657_),
    .Y(_03120_));
 sky130_fd_sc_hd__a21oi_2 _26103_ (.A1(_03119_),
    .A2(_03120_),
    .B1(net149),
    .Y(_03122_));
 sky130_fd_sc_hd__a21o_1 _26104_ (.A1(_03119_),
    .A2(_03120_),
    .B1(net149),
    .X(_03123_));
 sky130_fd_sc_hd__o311a_2 _26105_ (.A1(_04179_),
    .A2(net57),
    .A3(_04266_),
    .B1(_03120_),
    .C1(net149),
    .X(_03124_));
 sky130_fd_sc_hd__o211ai_4 _26106_ (.A1(_04179_),
    .A2(_08660_),
    .B1(net149),
    .C1(_03120_),
    .Y(_03125_));
 sky130_fd_sc_hd__o211ai_2 _26107_ (.A1(net237),
    .A2(_09297_),
    .B1(_03123_),
    .C1(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__o21ai_1 _26108_ (.A1(_03122_),
    .A2(_03124_),
    .B1(net145),
    .Y(_03127_));
 sky130_fd_sc_hd__o22ai_4 _26109_ (.A1(net237),
    .A2(_09297_),
    .B1(_03122_),
    .B2(_03124_),
    .Y(_03128_));
 sky130_fd_sc_hd__nand3_4 _26110_ (.A(_03123_),
    .B(_03125_),
    .C(_09299_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand3_4 _26111_ (.A(_03117_),
    .B(_03128_),
    .C(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__inv_2 _26112_ (.A(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__a21oi_1 _26113_ (.A1(_03128_),
    .A2(_03129_),
    .B1(_03117_),
    .Y(_03133_));
 sky130_fd_sc_hd__nand3_4 _26114_ (.A(_03118_),
    .B(_03126_),
    .C(_03127_),
    .Y(_03134_));
 sky130_fd_sc_hd__a2bb2oi_1 _26115_ (.A1_N(net140),
    .A2_N(net136),
    .B1(_03130_),
    .B2(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__a22o_1 _26116_ (.A1(net139),
    .A2(_10544_),
    .B1(_03130_),
    .B2(_03134_),
    .X(_03136_));
 sky130_fd_sc_hd__a31oi_4 _26117_ (.A1(_03117_),
    .A2(_03128_),
    .A3(_03129_),
    .B1(_10546_),
    .Y(_03137_));
 sky130_fd_sc_hd__nand2_1 _26118_ (.A(_03137_),
    .B(_03134_),
    .Y(_03138_));
 sky130_fd_sc_hd__o211a_1 _26119_ (.A1(net140),
    .A2(net136),
    .B1(_03130_),
    .C1(_03134_),
    .X(_03139_));
 sky130_fd_sc_hd__o211ai_2 _26120_ (.A1(net140),
    .A2(net136),
    .B1(_03130_),
    .C1(_03134_),
    .Y(_03140_));
 sky130_fd_sc_hd__a21oi_1 _26121_ (.A1(_03130_),
    .A2(_03134_),
    .B1(_10546_),
    .Y(_03141_));
 sky130_fd_sc_hd__a21o_1 _26122_ (.A1(_03130_),
    .A2(_03134_),
    .B1(_10546_),
    .X(_03142_));
 sky130_fd_sc_hd__a221oi_4 _26123_ (.A1(_03137_),
    .A2(_03134_),
    .B1(_02972_),
    .B2(_02966_),
    .C1(_03135_),
    .Y(_03144_));
 sky130_fd_sc_hd__o21ai_2 _26124_ (.A1(_03139_),
    .A2(_03141_),
    .B1(_03116_),
    .Y(_03145_));
 sky130_fd_sc_hd__a21oi_2 _26125_ (.A1(_03136_),
    .A2(_03138_),
    .B1(_03116_),
    .Y(_03146_));
 sky130_fd_sc_hd__o211ai_4 _26126_ (.A1(_02967_),
    .A2(_03115_),
    .B1(_03140_),
    .C1(_03142_),
    .Y(_03147_));
 sky130_fd_sc_hd__o21ai_1 _26127_ (.A1(_03144_),
    .A2(_03146_),
    .B1(_12098_),
    .Y(_03148_));
 sky130_fd_sc_hd__o21ai_2 _26128_ (.A1(net141),
    .A2(_11742_),
    .B1(_03147_),
    .Y(_03149_));
 sky130_fd_sc_hd__o22ai_4 _26129_ (.A1(net141),
    .A2(_11742_),
    .B1(_03144_),
    .B2(_03146_),
    .Y(_03150_));
 sky130_fd_sc_hd__o2111ai_4 _26130_ (.A1(_11737_),
    .A2(_11740_),
    .B1(_03147_),
    .C1(net143),
    .D1(_03145_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand3_2 _26131_ (.A(_03113_),
    .B(_03150_),
    .C(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__o211ai_4 _26132_ (.A1(_03149_),
    .A2(_03144_),
    .B1(_03114_),
    .C1(_03148_),
    .Y(_03153_));
 sky130_fd_sc_hd__o211a_1 _26133_ (.A1(net131),
    .A2(_00366_),
    .B1(_03152_),
    .C1(_03153_),
    .X(_03155_));
 sky130_fd_sc_hd__o211ai_2 _26134_ (.A1(net131),
    .A2(_00366_),
    .B1(_03152_),
    .C1(_03153_),
    .Y(_03156_));
 sky130_fd_sc_hd__a21oi_1 _26135_ (.A1(_03152_),
    .A2(_03153_),
    .B1(net129),
    .Y(_03157_));
 sky130_fd_sc_hd__a21o_1 _26136_ (.A1(_03152_),
    .A2(_03153_),
    .B1(net129),
    .X(_03158_));
 sky130_fd_sc_hd__o2bb2ai_4 _26137_ (.A1_N(_02987_),
    .A2_N(_02991_),
    .B1(_03155_),
    .B2(_03157_),
    .Y(_03159_));
 sky130_fd_sc_hd__o2111ai_4 _26138_ (.A1(_02988_),
    .A2(net129),
    .B1(_02987_),
    .C1(_03156_),
    .D1(_03158_),
    .Y(_03160_));
 sky130_fd_sc_hd__a22o_1 _26139_ (.A1(_02712_),
    .A2(_02947_),
    .B1(_03159_),
    .B2(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__o2111ai_4 _26140_ (.A1(_02944_),
    .A2(_02706_),
    .B1(_02712_),
    .C1(_03159_),
    .D1(_03160_),
    .Y(_03162_));
 sky130_fd_sc_hd__o211ai_2 _26141_ (.A1(_02711_),
    .A2(_02945_),
    .B1(_03159_),
    .C1(_03160_),
    .Y(_03163_));
 sky130_fd_sc_hd__a21o_1 _26142_ (.A1(_03159_),
    .A2(_03160_),
    .B1(_02949_),
    .X(_03164_));
 sky130_fd_sc_hd__a32oi_4 _26143_ (.A1(_02950_),
    .A2(_02994_),
    .A3(_02995_),
    .B1(_02997_),
    .B2(_02949_),
    .Y(_03166_));
 sky130_fd_sc_hd__o2111a_1 _26144_ (.A1(_02998_),
    .A2(_02949_),
    .B1(_02997_),
    .C1(_03163_),
    .D1(_03164_),
    .X(_03167_));
 sky130_fd_sc_hd__o2111ai_4 _26145_ (.A1(_02998_),
    .A2(_02949_),
    .B1(_02997_),
    .C1(_03163_),
    .D1(_03164_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand3_4 _26146_ (.A(_03161_),
    .B(_03162_),
    .C(_03166_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand4_2 _26147_ (.A(_03109_),
    .B(_03111_),
    .C(_03168_),
    .D(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__a22o_1 _26148_ (.A1(_03109_),
    .A2(_03111_),
    .B1(_03168_),
    .B2(_03169_),
    .X(_03171_));
 sky130_fd_sc_hd__nand4_1 _26149_ (.A(_03107_),
    .B(_03108_),
    .C(_03168_),
    .D(_03169_),
    .Y(_03172_));
 sky130_fd_sc_hd__a22o_1 _26150_ (.A1(_03107_),
    .A2(_03108_),
    .B1(_03168_),
    .B2(_03169_),
    .X(_03173_));
 sky130_fd_sc_hd__o2111ai_4 _26151_ (.A1(_03006_),
    .A2(_02943_),
    .B1(_03005_),
    .C1(_03170_),
    .D1(_03171_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand3_1 _26152_ (.A(_03037_),
    .B(_03172_),
    .C(_03173_),
    .Y(_03175_));
 sky130_fd_sc_hd__o311a_1 _26153_ (.A1(_02767_),
    .A2(_02800_),
    .A3(_02802_),
    .B1(_02933_),
    .C1(_02769_),
    .X(_03178_));
 sky130_fd_sc_hd__nor2_1 _26154_ (.A(_02932_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__o2bb2ai_1 _26155_ (.A1_N(_03174_),
    .A2_N(_03175_),
    .B1(_03178_),
    .B2(_02932_),
    .Y(_03180_));
 sky130_fd_sc_hd__nand3_1 _26156_ (.A(_03174_),
    .B(_03175_),
    .C(_03179_),
    .Y(_03181_));
 sky130_fd_sc_hd__a22oi_2 _26157_ (.A1(_03016_),
    .A2(_03035_),
    .B1(_03180_),
    .B2(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__nand2_1 _26158_ (.A(_03182_),
    .B(_02923_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand4_1 _26159_ (.A(_03016_),
    .B(_03035_),
    .C(_03180_),
    .D(_03181_),
    .Y(_03184_));
 sky130_fd_sc_hd__o21ai_1 _26160_ (.A1(_02923_),
    .A2(_03182_),
    .B1(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__o21a_1 _26161_ (.A1(_02923_),
    .A2(_03182_),
    .B1(_03184_),
    .X(_03186_));
 sky130_fd_sc_hd__nand2_1 _26162_ (.A(_03183_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__and4b_1 _26163_ (.A_N(_02923_),
    .B(_03036_),
    .C(_03180_),
    .D(_03181_),
    .X(_03189_));
 sky130_fd_sc_hd__or2_1 _26164_ (.A(_02923_),
    .B(_03184_),
    .X(_03190_));
 sky130_fd_sc_hd__a211oi_1 _26165_ (.A1(_03183_),
    .A2(_03186_),
    .B1(_03189_),
    .C1(_03034_),
    .Y(_03191_));
 sky130_fd_sc_hd__a22oi_4 _26166_ (.A1(_03022_),
    .A2(_03027_),
    .B1(_03187_),
    .B2(_03190_),
    .Y(_03192_));
 sky130_fd_sc_hd__nor2_1 _26167_ (.A(_03191_),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__and4_1 _26168_ (.A(_02841_),
    .B(_02843_),
    .C(_03029_),
    .D(_03030_),
    .X(_03194_));
 sky130_fd_sc_hd__nand3_1 _26169_ (.A(_02435_),
    .B(_02639_),
    .C(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__and4_1 _26170_ (.A(_02435_),
    .B(_02438_),
    .C(_02639_),
    .D(_03194_),
    .X(_03196_));
 sky130_fd_sc_hd__o221ai_4 _26171_ (.A1(_01479_),
    .A2(_01482_),
    .B1(_01481_),
    .B2(_12401_),
    .C1(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__o21ai_1 _26172_ (.A1(_02843_),
    .A2(_03028_),
    .B1(_03030_),
    .Y(_03198_));
 sky130_fd_sc_hd__a21oi_1 _26173_ (.A1(_02846_),
    .A2(_03194_),
    .B1(_03198_),
    .Y(_03200_));
 sky130_fd_sc_hd__o21a_2 _26174_ (.A1(_02437_),
    .A2(_03195_),
    .B1(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__nand2_1 _26175_ (.A(_03197_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__xor2_1 _26176_ (.A(_03193_),
    .B(_03202_),
    .X(net116));
 sky130_fd_sc_hd__nand2_1 _26177_ (.A(_03093_),
    .B(_03095_),
    .Y(_03203_));
 sky130_fd_sc_hd__a21boi_2 _26178_ (.A1(_03174_),
    .A2(_03179_),
    .B1_N(_03175_),
    .Y(_03204_));
 sky130_fd_sc_hd__o21ai_1 _26179_ (.A1(_03167_),
    .A2(_03112_),
    .B1(_03169_),
    .Y(_03205_));
 sky130_fd_sc_hd__a32o_1 _26180_ (.A1(_07072_),
    .A2(net170),
    .A3(net238),
    .B1(_08006_),
    .B2(net20),
    .X(_03206_));
 sky130_fd_sc_hd__nand2_1 _26181_ (.A(_03085_),
    .B(_03090_),
    .Y(_03207_));
 sky130_fd_sc_hd__a22oi_1 _26182_ (.A1(_07504_),
    .A2(_07642_),
    .B1(_07643_),
    .B2(net21),
    .Y(_03208_));
 sky130_fd_sc_hd__a32o_1 _26183_ (.A1(_07499_),
    .A2(_07503_),
    .A3(_07642_),
    .B1(_07643_),
    .B2(net21),
    .X(_03210_));
 sky130_fd_sc_hd__a21oi_1 _26184_ (.A1(_03072_),
    .A2(_03081_),
    .B1(_03078_),
    .Y(_03211_));
 sky130_fd_sc_hd__a32o_1 _26185_ (.A1(_07771_),
    .A2(net239),
    .A3(net166),
    .B1(_07308_),
    .B2(net22),
    .X(_03212_));
 sky130_fd_sc_hd__a32oi_4 _26186_ (.A1(_08204_),
    .A2(net163),
    .A3(net269),
    .B1(_07225_),
    .B2(net24),
    .Y(_03213_));
 sky130_fd_sc_hd__o21ai_1 _26187_ (.A1(net160),
    .A2(_08666_),
    .B1(net240),
    .Y(_03214_));
 sky130_fd_sc_hd__nor2_2 _26188_ (.A(net319),
    .B(_06866_),
    .Y(_03215_));
 sky130_fd_sc_hd__or3_1 _26189_ (.A(net51),
    .B(net319),
    .C(_04190_),
    .X(_03216_));
 sky130_fd_sc_hd__a21oi_1 _26190_ (.A1(_03214_),
    .A2(_03216_),
    .B1(_03213_),
    .Y(_03217_));
 sky130_fd_sc_hd__a21o_1 _26191_ (.A1(_03214_),
    .A2(_03216_),
    .B1(_03213_),
    .X(_03218_));
 sky130_fd_sc_hd__o221a_1 _26192_ (.A1(net319),
    .A2(_06866_),
    .B1(_06864_),
    .B2(_08669_),
    .C1(_03213_),
    .X(_03219_));
 sky130_fd_sc_hd__o221ai_4 _26193_ (.A1(net319),
    .A2(_06866_),
    .B1(_06864_),
    .B2(_08669_),
    .C1(_03213_),
    .Y(_03221_));
 sky130_fd_sc_hd__nand3_2 _26194_ (.A(_03212_),
    .B(_03218_),
    .C(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__o21bai_1 _26195_ (.A1(_03217_),
    .A2(_03219_),
    .B1_N(_03212_),
    .Y(_03223_));
 sky130_fd_sc_hd__o21ai_1 _26196_ (.A1(_03217_),
    .A2(_03219_),
    .B1(_03212_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand3b_1 _26197_ (.A_N(_03212_),
    .B(_03218_),
    .C(_03221_),
    .Y(_03225_));
 sky130_fd_sc_hd__o211ai_2 _26198_ (.A1(_03078_),
    .A2(_03083_),
    .B1(_03222_),
    .C1(_03223_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand3_1 _26199_ (.A(_03224_),
    .B(_03225_),
    .C(_03211_),
    .Y(_03227_));
 sky130_fd_sc_hd__nand3_1 _26200_ (.A(_03223_),
    .B(_03211_),
    .C(_03222_),
    .Y(_03228_));
 sky130_fd_sc_hd__o211ai_1 _26201_ (.A1(_03078_),
    .A2(_03083_),
    .B1(_03224_),
    .C1(_03225_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand3_1 _26202_ (.A(_03210_),
    .B(_03226_),
    .C(_03227_),
    .Y(_03230_));
 sky130_fd_sc_hd__nand3_1 _26203_ (.A(_03229_),
    .B(_03208_),
    .C(_03228_),
    .Y(_03232_));
 sky130_fd_sc_hd__nand3_1 _26204_ (.A(_03226_),
    .B(_03227_),
    .C(_03208_),
    .Y(_03233_));
 sky130_fd_sc_hd__nand3_1 _26205_ (.A(_03210_),
    .B(_03228_),
    .C(_03229_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand3_2 _26206_ (.A(_03207_),
    .B(_03230_),
    .C(_03232_),
    .Y(_03235_));
 sky130_fd_sc_hd__nand4_2 _26207_ (.A(_03085_),
    .B(_03090_),
    .C(_03233_),
    .D(_03234_),
    .Y(_03236_));
 sky130_fd_sc_hd__a21o_1 _26208_ (.A1(_03235_),
    .A2(_03236_),
    .B1(_03206_),
    .X(_03237_));
 sky130_fd_sc_hd__nand3_2 _26209_ (.A(_03206_),
    .B(_03235_),
    .C(_03236_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand2_1 _26210_ (.A(_03237_),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__nand2_1 _26211_ (.A(_03047_),
    .B(_03051_),
    .Y(_03240_));
 sky130_fd_sc_hd__a21oi_1 _26212_ (.A1(net273),
    .A2(net160),
    .B1(_03038_),
    .Y(_03241_));
 sky130_fd_sc_hd__a31o_1 _26213_ (.A1(net319),
    .A2(net163),
    .A3(net273),
    .B1(_03038_),
    .X(_03243_));
 sky130_fd_sc_hd__o2111ai_1 _26214_ (.A1(_06028_),
    .A2(net153),
    .B1(_02857_),
    .C1(_02860_),
    .D1(_03241_),
    .Y(_03244_));
 sky130_fd_sc_hd__a31o_1 _26215_ (.A1(_02857_),
    .A2(_02860_),
    .A3(_03041_),
    .B1(_03241_),
    .X(_03245_));
 sky130_fd_sc_hd__a31o_1 _26216_ (.A1(_02857_),
    .A2(_02860_),
    .A3(_03041_),
    .B1(_03243_),
    .X(_03246_));
 sky130_fd_sc_hd__nand2_1 _26217_ (.A(_03042_),
    .B(_03243_),
    .Y(_03247_));
 sky130_fd_sc_hd__o211ai_4 _26218_ (.A1(_02536_),
    .A2(_02696_),
    .B1(_03246_),
    .C1(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__nand3_2 _26219_ (.A(_03245_),
    .B(_02699_),
    .C(_03244_),
    .Y(_03249_));
 sky130_fd_sc_hd__nand2_2 _26220_ (.A(_03248_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__a21boi_1 _26221_ (.A1(_03248_),
    .A2(_03249_),
    .B1_N(_03046_),
    .Y(_03251_));
 sky130_fd_sc_hd__o2111a_1 _26222_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_03043_),
    .C1(_03248_),
    .D1(_03249_),
    .X(_03252_));
 sky130_fd_sc_hd__o2111ai_2 _26223_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_03043_),
    .C1(_03248_),
    .D1(_03249_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand3b_2 _26224_ (.A_N(_03251_),
    .B(_03254_),
    .C(_02703_),
    .Y(_03255_));
 sky130_fd_sc_hd__o22ai_2 _26225_ (.A1(_02159_),
    .A2(_02701_),
    .B1(_03251_),
    .B2(_03252_),
    .Y(_03256_));
 sky130_fd_sc_hd__and2_1 _26226_ (.A(_03255_),
    .B(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__o2bb2ai_2 _26227_ (.A1_N(_03056_),
    .A2_N(_03062_),
    .B1(_03240_),
    .B2(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__a21o_1 _26228_ (.A1(_03250_),
    .A2(_02857_),
    .B1(_02704_),
    .X(_03259_));
 sky130_fd_sc_hd__o2111ai_4 _26229_ (.A1(_05763_),
    .A2(net153),
    .B1(_02704_),
    .C1(_02741_),
    .D1(_03250_),
    .Y(_03260_));
 sky130_fd_sc_hd__o21ai_1 _26230_ (.A1(_03046_),
    .A2(_03250_),
    .B1(_03249_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand3_1 _26231_ (.A(_03259_),
    .B(_03260_),
    .C(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__inv_2 _26232_ (.A(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__and4_2 _26233_ (.A(_02857_),
    .B(_03250_),
    .C(_02700_),
    .D(_02704_),
    .X(_03265_));
 sky130_fd_sc_hd__or4_1 _26234_ (.A(_02740_),
    .B(_03248_),
    .C(_02856_),
    .D(_02703_),
    .X(_03266_));
 sky130_fd_sc_hd__o21ai_1 _26235_ (.A1(_02699_),
    .A2(_03260_),
    .B1(_03262_),
    .Y(_03267_));
 sky130_fd_sc_hd__a31o_1 _26236_ (.A1(_03240_),
    .A2(_03255_),
    .A3(_03256_),
    .B1(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__a31oi_2 _26237_ (.A1(_03240_),
    .A2(_03255_),
    .A3(_03256_),
    .B1(_03267_),
    .Y(_03269_));
 sky130_fd_sc_hd__a22o_1 _26238_ (.A1(_03237_),
    .A2(_03238_),
    .B1(_03258_),
    .B2(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__nand4_2 _26239_ (.A(_03237_),
    .B(_03238_),
    .C(_03258_),
    .D(_03269_),
    .Y(_03271_));
 sky130_fd_sc_hd__o2bb2ai_2 _26240_ (.A1_N(_03270_),
    .A2_N(_03271_),
    .B1(_00364_),
    .B2(_02708_),
    .Y(_03272_));
 sky130_fd_sc_hd__nand4_4 _26241_ (.A(_03270_),
    .B(net131),
    .C(_02709_),
    .D(_03271_),
    .Y(_03273_));
 sky130_fd_sc_hd__inv_2 _26242_ (.A(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_1 _26243_ (.A(_03063_),
    .B(_03097_),
    .Y(_03276_));
 sky130_fd_sc_hd__a22o_1 _26244_ (.A1(_03272_),
    .A2(_03273_),
    .B1(_03276_),
    .B2(_03064_),
    .X(_03277_));
 sky130_fd_sc_hd__nand3_2 _26245_ (.A(_03064_),
    .B(_03272_),
    .C(_03276_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand4_1 _26246_ (.A(_03064_),
    .B(_03272_),
    .C(_03273_),
    .D(_03276_),
    .Y(_03279_));
 sky130_fd_sc_hd__o21ai_2 _26247_ (.A1(_03274_),
    .A2(_03278_),
    .B1(_03277_),
    .Y(_03280_));
 sky130_fd_sc_hd__a311oi_2 _26248_ (.A1(_03136_),
    .A2(_03138_),
    .A3(_03116_),
    .B1(_11742_),
    .C1(net141),
    .Y(_03281_));
 sky130_fd_sc_hd__o32a_1 _26249_ (.A1(_03116_),
    .A2(_03139_),
    .A3(_03141_),
    .B1(_12099_),
    .B2(_03144_),
    .X(_03282_));
 sky130_fd_sc_hd__a21o_1 _26250_ (.A1(_03130_),
    .A2(_10545_),
    .B1(_03133_),
    .X(_03283_));
 sky130_fd_sc_hd__a32o_1 _26251_ (.A1(_03117_),
    .A2(_03128_),
    .A3(_03129_),
    .B1(_03134_),
    .B2(_10546_),
    .X(_03284_));
 sky130_fd_sc_hd__a21oi_2 _26252_ (.A1(net144),
    .A2(_03125_),
    .B1(_03122_),
    .Y(_03285_));
 sky130_fd_sc_hd__o21ai_2 _26253_ (.A1(_09299_),
    .A2(_03124_),
    .B1(_03123_),
    .Y(_03288_));
 sky130_fd_sc_hd__or3_1 _26254_ (.A(net57),
    .B(_04266_),
    .C(_04201_),
    .X(_03289_));
 sky130_fd_sc_hd__nand3_2 _26255_ (.A(net192),
    .B(_06762_),
    .C(_08657_),
    .Y(_03290_));
 sky130_fd_sc_hd__o311a_2 _26256_ (.A1(_08658_),
    .A2(net190),
    .A3(_06756_),
    .B1(_03289_),
    .C1(net149),
    .X(_03291_));
 sky130_fd_sc_hd__o221ai_4 _26257_ (.A1(_04201_),
    .A2(_08660_),
    .B1(net152),
    .B2(_03286_),
    .C1(_03290_),
    .Y(_03292_));
 sky130_fd_sc_hd__a21oi_1 _26258_ (.A1(_03289_),
    .A2(_03290_),
    .B1(net149),
    .Y(_03293_));
 sky130_fd_sc_hd__a21o_2 _26259_ (.A1(_03289_),
    .A2(_03290_),
    .B1(net149),
    .X(_03294_));
 sky130_fd_sc_hd__o211ai_4 _26260_ (.A1(net237),
    .A2(_09297_),
    .B1(_03292_),
    .C1(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__o21ai_2 _26261_ (.A1(_03291_),
    .A2(_03293_),
    .B1(_09299_),
    .Y(_03296_));
 sky130_fd_sc_hd__o21ai_2 _26262_ (.A1(_03291_),
    .A2(_03293_),
    .B1(net144),
    .Y(_03297_));
 sky130_fd_sc_hd__o2111ai_4 _26263_ (.A1(_04495_),
    .A2(net152),
    .B1(_08882_),
    .C1(_03292_),
    .D1(_03294_),
    .Y(_03299_));
 sky130_fd_sc_hd__nand3_4 _26264_ (.A(_03297_),
    .B(_03299_),
    .C(_03285_),
    .Y(_03300_));
 sky130_fd_sc_hd__inv_2 _26265_ (.A(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand3_4 _26266_ (.A(_03288_),
    .B(_03295_),
    .C(_03296_),
    .Y(_03302_));
 sky130_fd_sc_hd__a22o_1 _26267_ (.A1(net139),
    .A2(_10544_),
    .B1(_03300_),
    .B2(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__nand4_2 _26268_ (.A(net139),
    .B(_10544_),
    .C(_03300_),
    .D(_03302_),
    .Y(_03304_));
 sky130_fd_sc_hd__o211ai_4 _26269_ (.A1(net140),
    .A2(_10542_),
    .B1(_03300_),
    .C1(_03302_),
    .Y(_03305_));
 sky130_fd_sc_hd__a21o_2 _26270_ (.A1(_03300_),
    .A2(_03302_),
    .B1(_10546_),
    .X(_03306_));
 sky130_fd_sc_hd__a2bb2oi_2 _26271_ (.A1_N(_03133_),
    .A2_N(_03137_),
    .B1(_03305_),
    .B2(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand3_4 _26272_ (.A(_03303_),
    .B(_03304_),
    .C(_03283_),
    .Y(_03308_));
 sky130_fd_sc_hd__a21oi_2 _26273_ (.A1(_03303_),
    .A2(_03304_),
    .B1(_03283_),
    .Y(_03310_));
 sky130_fd_sc_hd__o2111ai_4 _26274_ (.A1(_10546_),
    .A2(_03131_),
    .B1(_03134_),
    .C1(_03305_),
    .D1(_03306_),
    .Y(_03311_));
 sky130_fd_sc_hd__o2bb2ai_2 _26275_ (.A1_N(_03308_),
    .A2_N(_03311_),
    .B1(net141),
    .B2(_11742_),
    .Y(_03312_));
 sky130_fd_sc_hd__o2111ai_4 _26276_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net143),
    .C1(_03308_),
    .D1(_03311_),
    .Y(_03313_));
 sky130_fd_sc_hd__a31oi_4 _26277_ (.A1(_03284_),
    .A2(_03305_),
    .A3(_03306_),
    .B1(_12098_),
    .Y(_03314_));
 sky130_fd_sc_hd__nand2_1 _26278_ (.A(_03314_),
    .B(_03308_),
    .Y(_03315_));
 sky130_fd_sc_hd__o21ai_1 _26279_ (.A1(_03307_),
    .A2(_03310_),
    .B1(_12098_),
    .Y(_03316_));
 sky130_fd_sc_hd__a22oi_2 _26280_ (.A1(_03145_),
    .A2(_03149_),
    .B1(_03312_),
    .B2(_03313_),
    .Y(_03317_));
 sky130_fd_sc_hd__nand3_1 _26281_ (.A(_03316_),
    .B(_03282_),
    .C(_03315_),
    .Y(_03318_));
 sky130_fd_sc_hd__o211a_1 _26282_ (.A1(_03146_),
    .A2(_03281_),
    .B1(_03312_),
    .C1(_03313_),
    .X(_03319_));
 sky130_fd_sc_hd__o211ai_2 _26283_ (.A1(_03146_),
    .A2(_03281_),
    .B1(_03312_),
    .C1(_03313_),
    .Y(_03321_));
 sky130_fd_sc_hd__o21ai_2 _26284_ (.A1(_03317_),
    .A2(_03319_),
    .B1(net129),
    .Y(_03322_));
 sky130_fd_sc_hd__a31o_1 _26285_ (.A1(_03315_),
    .A2(_03316_),
    .A3(_03282_),
    .B1(net129),
    .X(_03323_));
 sky130_fd_sc_hd__o2111ai_1 _26286_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_03318_),
    .D1(_03321_),
    .Y(_03324_));
 sky130_fd_sc_hd__a32oi_4 _26287_ (.A1(_03113_),
    .A2(_03150_),
    .A3(_03151_),
    .B1(_03153_),
    .B2(net129),
    .Y(_03325_));
 sky130_fd_sc_hd__a21oi_1 _26288_ (.A1(_03322_),
    .A2(_03324_),
    .B1(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__a21o_1 _26289_ (.A1(_03322_),
    .A2(_03324_),
    .B1(_03325_),
    .X(_03327_));
 sky130_fd_sc_hd__o211a_1 _26290_ (.A1(_03319_),
    .A2(_03323_),
    .B1(_03325_),
    .C1(_03322_),
    .X(_03328_));
 sky130_fd_sc_hd__o211ai_2 _26291_ (.A1(_03319_),
    .A2(_03323_),
    .B1(_03325_),
    .C1(_03322_),
    .Y(_03329_));
 sky130_fd_sc_hd__a22o_1 _26292_ (.A1(_02712_),
    .A2(_02947_),
    .B1(_03327_),
    .B2(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__o2111ai_1 _26293_ (.A1(_02944_),
    .A2(_02706_),
    .B1(_02712_),
    .C1(_03327_),
    .D1(_03329_),
    .Y(_03332_));
 sky130_fd_sc_hd__o211ai_1 _26294_ (.A1(_02711_),
    .A2(_02945_),
    .B1(_03327_),
    .C1(_03329_),
    .Y(_03333_));
 sky130_fd_sc_hd__o21ai_1 _26295_ (.A1(_03326_),
    .A2(_03328_),
    .B1(_02948_),
    .Y(_03334_));
 sky130_fd_sc_hd__a21boi_1 _26296_ (.A1(_02948_),
    .A2(_03160_),
    .B1_N(_03159_),
    .Y(_03335_));
 sky130_fd_sc_hd__and3_1 _26297_ (.A(_03333_),
    .B(_03334_),
    .C(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__nand3_2 _26298_ (.A(_03333_),
    .B(_03334_),
    .C(_03335_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand3b_2 _26299_ (.A_N(_03335_),
    .B(_03332_),
    .C(_03330_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand3_1 _26300_ (.A(_03280_),
    .B(_03337_),
    .C(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__a21o_1 _26301_ (.A1(_03337_),
    .A2(_03338_),
    .B1(_03280_),
    .X(_03340_));
 sky130_fd_sc_hd__o2111ai_1 _26302_ (.A1(_03278_),
    .A2(_03274_),
    .B1(_03277_),
    .C1(_03337_),
    .D1(_03338_),
    .Y(_03341_));
 sky130_fd_sc_hd__a22o_1 _26303_ (.A1(_03277_),
    .A2(_03279_),
    .B1(_03337_),
    .B2(_03338_),
    .X(_03343_));
 sky130_fd_sc_hd__nand3_1 _26304_ (.A(_03343_),
    .B(_03205_),
    .C(_03341_),
    .Y(_03344_));
 sky130_fd_sc_hd__o2111ai_2 _26305_ (.A1(_03112_),
    .A2(_03167_),
    .B1(_03169_),
    .C1(_03339_),
    .D1(_03340_),
    .Y(_03345_));
 sky130_fd_sc_hd__a32o_1 _26306_ (.A1(_02712_),
    .A2(_03098_),
    .A3(_03100_),
    .B1(_03104_),
    .B2(_03106_),
    .X(_03346_));
 sky130_fd_sc_hd__nand3_1 _26307_ (.A(_03344_),
    .B(_03345_),
    .C(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__a21o_1 _26308_ (.A1(_03344_),
    .A2(_03345_),
    .B1(_03346_),
    .X(_03348_));
 sky130_fd_sc_hd__a21o_1 _26309_ (.A1(_03347_),
    .A2(_03348_),
    .B1(_03204_),
    .X(_03349_));
 sky130_fd_sc_hd__nand3_1 _26310_ (.A(_03204_),
    .B(_03347_),
    .C(_03348_),
    .Y(_03350_));
 sky130_fd_sc_hd__a32o_1 _26311_ (.A1(_03204_),
    .A2(_03347_),
    .A3(_03348_),
    .B1(_03095_),
    .B2(_03093_),
    .X(_03351_));
 sky130_fd_sc_hd__nand3_1 _26312_ (.A(_03203_),
    .B(_03349_),
    .C(_03350_),
    .Y(_03352_));
 sky130_fd_sc_hd__a21o_1 _26313_ (.A1(_03349_),
    .A2(_03350_),
    .B1(_03203_),
    .X(_03354_));
 sky130_fd_sc_hd__nand3_1 _26314_ (.A(_03354_),
    .B(_03185_),
    .C(_03352_),
    .Y(_03355_));
 sky130_fd_sc_hd__a21o_1 _26315_ (.A1(_03352_),
    .A2(_03354_),
    .B1(_03185_),
    .X(_03356_));
 sky130_fd_sc_hd__nand2_1 _26316_ (.A(_03355_),
    .B(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__o21ba_1 _26317_ (.A1(_03192_),
    .A2(_03202_),
    .B1_N(_03191_),
    .X(_03358_));
 sky130_fd_sc_hd__xnor2_1 _26318_ (.A(_03357_),
    .B(_03358_),
    .Y(net117));
 sky130_fd_sc_hd__nand2_1 _26319_ (.A(_03349_),
    .B(_03351_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand2_1 _26320_ (.A(_03235_),
    .B(_03238_),
    .Y(_03360_));
 sky130_fd_sc_hd__nand2_1 _26321_ (.A(_03344_),
    .B(_03346_),
    .Y(_03361_));
 sky130_fd_sc_hd__nand2_1 _26322_ (.A(_03345_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__o21ai_1 _26323_ (.A1(_03280_),
    .A2(_03336_),
    .B1(_03338_),
    .Y(_03364_));
 sky130_fd_sc_hd__and3_1 _26324_ (.A(_07499_),
    .B(_07503_),
    .C(net238),
    .X(_03365_));
 sky130_fd_sc_hd__and3_1 _26325_ (.A(_04266_),
    .B(net54),
    .C(net21),
    .X(_03366_));
 sky130_fd_sc_hd__a31o_1 _26326_ (.A1(_07499_),
    .A2(_07503_),
    .A3(net238),
    .B1(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__and3b_1 _26327_ (.A_N(net54),
    .B(net22),
    .C(net53),
    .X(_03368_));
 sky130_fd_sc_hd__o311a_1 _26328_ (.A1(net233),
    .A2(_05927_),
    .A3(_07767_),
    .B1(_07771_),
    .C1(_07642_),
    .X(_03369_));
 sky130_fd_sc_hd__a31o_1 _26329_ (.A1(_07771_),
    .A2(_07642_),
    .A3(net166),
    .B1(_03368_),
    .X(_03370_));
 sky130_fd_sc_hd__a21o_1 _26330_ (.A1(_03212_),
    .A2(_03221_),
    .B1(_03217_),
    .X(_03371_));
 sky130_fd_sc_hd__a32o_2 _26331_ (.A1(_08204_),
    .A2(net163),
    .A3(net239),
    .B1(_07308_),
    .B2(net24),
    .X(_03372_));
 sky130_fd_sc_hd__o311a_1 _26332_ (.A1(net22),
    .A2(net24),
    .A3(_07503_),
    .B1(net240),
    .C1(net319),
    .X(_03373_));
 sky130_fd_sc_hd__a21oi_4 _26333_ (.A1(_06863_),
    .A2(net160),
    .B1(_03215_),
    .Y(_03375_));
 sky130_fd_sc_hd__nor2_2 _26334_ (.A(net319),
    .B(_07226_),
    .Y(_03376_));
 sky130_fd_sc_hd__a21oi_2 _26335_ (.A1(net153),
    .A2(net158),
    .B1(_07224_),
    .Y(_03377_));
 sky130_fd_sc_hd__o221ai_4 _26336_ (.A1(net319),
    .A2(_07226_),
    .B1(_07224_),
    .B2(_08669_),
    .C1(_03375_),
    .Y(_03378_));
 sky130_fd_sc_hd__o22a_1 _26337_ (.A1(_03215_),
    .A2(_03373_),
    .B1(_03376_),
    .B2(_03377_),
    .X(_03379_));
 sky130_fd_sc_hd__o22ai_4 _26338_ (.A1(_03215_),
    .A2(_03373_),
    .B1(_03376_),
    .B2(_03377_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand3_2 _26339_ (.A(_03372_),
    .B(_03378_),
    .C(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__a21o_1 _26340_ (.A1(_03378_),
    .A2(_03380_),
    .B1(_03372_),
    .X(_03382_));
 sky130_fd_sc_hd__a21bo_1 _26341_ (.A1(_03378_),
    .A2(_03380_),
    .B1_N(_03372_),
    .X(_03383_));
 sky130_fd_sc_hd__nand3b_1 _26342_ (.A_N(_03372_),
    .B(_03378_),
    .C(_03380_),
    .Y(_03384_));
 sky130_fd_sc_hd__nand3_2 _26343_ (.A(_03371_),
    .B(_03381_),
    .C(_03382_),
    .Y(_03386_));
 sky130_fd_sc_hd__nand4_1 _26344_ (.A(_03218_),
    .B(_03222_),
    .C(_03383_),
    .D(_03384_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand4_1 _26345_ (.A(_03218_),
    .B(_03222_),
    .C(_03381_),
    .D(_03382_),
    .Y(_03388_));
 sky130_fd_sc_hd__nand3_1 _26346_ (.A(_03371_),
    .B(_03383_),
    .C(_03384_),
    .Y(_03389_));
 sky130_fd_sc_hd__o211ai_2 _26347_ (.A1(_03368_),
    .A2(_03369_),
    .B1(_03386_),
    .C1(_03387_),
    .Y(_03390_));
 sky130_fd_sc_hd__nand3b_1 _26348_ (.A_N(_03370_),
    .B(_03386_),
    .C(_03387_),
    .Y(_03391_));
 sky130_fd_sc_hd__o211ai_1 _26349_ (.A1(_03368_),
    .A2(_03369_),
    .B1(_03388_),
    .C1(_03389_),
    .Y(_03392_));
 sky130_fd_sc_hd__nand4_1 _26350_ (.A(_03226_),
    .B(_03230_),
    .C(_03391_),
    .D(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__a22o_1 _26351_ (.A1(_03226_),
    .A2(_03230_),
    .B1(_03391_),
    .B2(_03392_),
    .X(_03394_));
 sky130_fd_sc_hd__o211a_1 _26352_ (.A1(_03365_),
    .A2(_03366_),
    .B1(_03393_),
    .C1(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__a21oi_1 _26353_ (.A1(_03393_),
    .A2(_03394_),
    .B1(_03367_),
    .Y(_03398_));
 sky130_fd_sc_hd__nor3_2 _26354_ (.A(_03268_),
    .B(_03395_),
    .C(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__o21a_1 _26355_ (.A1(_03395_),
    .A2(_03398_),
    .B1(_03268_),
    .X(_03400_));
 sky130_fd_sc_hd__nor3_1 _26356_ (.A(_02712_),
    .B(_03399_),
    .C(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__o32a_2 _26357_ (.A1(_11741_),
    .A2(_00360_),
    .A3(_02708_),
    .B1(_03399_),
    .B2(_03400_),
    .X(_03402_));
 sky130_fd_sc_hd__o21ai_1 _26358_ (.A1(_03268_),
    .A2(_03239_),
    .B1(_03258_),
    .Y(_03403_));
 sky130_fd_sc_hd__o21a_1 _26359_ (.A1(_03268_),
    .A2(_03239_),
    .B1(_03258_),
    .X(_03404_));
 sky130_fd_sc_hd__o21ai_1 _26360_ (.A1(_03401_),
    .A2(_03402_),
    .B1(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__o31ai_2 _26361_ (.A1(_02712_),
    .A2(_03399_),
    .A3(_03400_),
    .B1(_03403_),
    .Y(_03406_));
 sky130_fd_sc_hd__o21ai_2 _26362_ (.A1(_03402_),
    .A2(_03406_),
    .B1(_03405_),
    .Y(_03407_));
 sky130_fd_sc_hd__a21oi_1 _26363_ (.A1(_03321_),
    .A2(_00736_),
    .B1(_03317_),
    .Y(_03409_));
 sky130_fd_sc_hd__a21o_1 _26364_ (.A1(_03321_),
    .A2(_00736_),
    .B1(_03317_),
    .X(_03410_));
 sky130_fd_sc_hd__o21a_1 _26365_ (.A1(_09299_),
    .A2(_03291_),
    .B1(_03294_),
    .X(_03411_));
 sky130_fd_sc_hd__o21ai_1 _26366_ (.A1(_09299_),
    .A2(_03291_),
    .B1(_03294_),
    .Y(_03412_));
 sky130_fd_sc_hd__or3_1 _26367_ (.A(net57),
    .B(_04266_),
    .C(_04212_),
    .X(_03413_));
 sky130_fd_sc_hd__nand3_2 _26368_ (.A(_07072_),
    .B(net170),
    .C(_08657_),
    .Y(_03414_));
 sky130_fd_sc_hd__a21oi_1 _26369_ (.A1(_03413_),
    .A2(_03414_),
    .B1(net149),
    .Y(_03415_));
 sky130_fd_sc_hd__a21o_1 _26370_ (.A1(_03413_),
    .A2(_03414_),
    .B1(net149),
    .X(_03416_));
 sky130_fd_sc_hd__o311a_1 _26371_ (.A1(_04212_),
    .A2(_04266_),
    .A3(net57),
    .B1(net149),
    .C1(_03414_),
    .X(_03417_));
 sky130_fd_sc_hd__o211ai_2 _26372_ (.A1(_04212_),
    .A2(_08660_),
    .B1(net149),
    .C1(_03414_),
    .Y(_03418_));
 sky130_fd_sc_hd__o211ai_1 _26373_ (.A1(net237),
    .A2(_09297_),
    .B1(_03416_),
    .C1(_03418_),
    .Y(_03420_));
 sky130_fd_sc_hd__o21ai_1 _26374_ (.A1(_03415_),
    .A2(_03417_),
    .B1(_09299_),
    .Y(_03421_));
 sky130_fd_sc_hd__o22ai_2 _26375_ (.A1(net237),
    .A2(_09297_),
    .B1(_03415_),
    .B2(_03417_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand3_1 _26376_ (.A(_03416_),
    .B(_03418_),
    .C(_09299_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21oi_1 _26377_ (.A1(_03422_),
    .A2(_03423_),
    .B1(_03411_),
    .Y(_03424_));
 sky130_fd_sc_hd__nand3_1 _26378_ (.A(_03412_),
    .B(_03420_),
    .C(_03421_),
    .Y(_03425_));
 sky130_fd_sc_hd__nand3_1 _26379_ (.A(_03411_),
    .B(_03422_),
    .C(_03423_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand3_1 _26380_ (.A(_03412_),
    .B(_03422_),
    .C(_03423_),
    .Y(_03427_));
 sky130_fd_sc_hd__nand3_1 _26381_ (.A(_03421_),
    .B(_03411_),
    .C(_03420_),
    .Y(_03428_));
 sky130_fd_sc_hd__o211ai_4 _26382_ (.A1(net140),
    .A2(_10542_),
    .B1(_03427_),
    .C1(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__nand3_2 _26383_ (.A(_03425_),
    .B(_03426_),
    .C(_10545_),
    .Y(_03431_));
 sky130_fd_sc_hd__a31oi_2 _26384_ (.A1(_03288_),
    .A2(_03295_),
    .A3(_03296_),
    .B1(_10545_),
    .Y(_03432_));
 sky130_fd_sc_hd__a32oi_4 _26385_ (.A1(_03285_),
    .A2(_03297_),
    .A3(_03299_),
    .B1(_03302_),
    .B2(_10546_),
    .Y(_03433_));
 sky130_fd_sc_hd__o2bb2a_1 _26386_ (.A1_N(_03429_),
    .A2_N(_03431_),
    .B1(_03432_),
    .B2(_03301_),
    .X(_03434_));
 sky130_fd_sc_hd__o2bb2ai_4 _26387_ (.A1_N(_03429_),
    .A2_N(_03431_),
    .B1(_03432_),
    .B2(_03301_),
    .Y(_03435_));
 sky130_fd_sc_hd__and3_2 _26388_ (.A(_03433_),
    .B(_03431_),
    .C(_03429_),
    .X(_03436_));
 sky130_fd_sc_hd__nand3_4 _26389_ (.A(_03433_),
    .B(_03431_),
    .C(_03429_),
    .Y(_03437_));
 sky130_fd_sc_hd__a21oi_1 _26390_ (.A1(_03435_),
    .A2(_03437_),
    .B1(_12099_),
    .Y(_03438_));
 sky130_fd_sc_hd__a21o_1 _26391_ (.A1(_03435_),
    .A2(_03437_),
    .B1(_12099_),
    .X(_03439_));
 sky130_fd_sc_hd__o21ai_2 _26392_ (.A1(net141),
    .A2(_11742_),
    .B1(_03435_),
    .Y(_03440_));
 sky130_fd_sc_hd__o311a_1 _26393_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_03435_),
    .C1(_03437_),
    .X(_03442_));
 sky130_fd_sc_hd__o211ai_4 _26394_ (.A1(_11742_),
    .A2(net141),
    .B1(_03437_),
    .C1(_03435_),
    .Y(_03443_));
 sky130_fd_sc_hd__o21ai_1 _26395_ (.A1(_12098_),
    .A2(_03310_),
    .B1(_03308_),
    .Y(_03444_));
 sky130_fd_sc_hd__o221a_1 _26396_ (.A1(_03436_),
    .A2(_03440_),
    .B1(_03307_),
    .B2(_03314_),
    .C1(_03439_),
    .X(_03445_));
 sky130_fd_sc_hd__o221ai_4 _26397_ (.A1(_03436_),
    .A2(_03440_),
    .B1(_03307_),
    .B2(_03314_),
    .C1(_03439_),
    .Y(_03446_));
 sky130_fd_sc_hd__a21oi_1 _26398_ (.A1(_03439_),
    .A2(_03443_),
    .B1(_03444_),
    .Y(_03447_));
 sky130_fd_sc_hd__o221ai_2 _26399_ (.A1(_12098_),
    .A2(_03310_),
    .B1(_03438_),
    .B2(_03442_),
    .C1(_03308_),
    .Y(_03448_));
 sky130_fd_sc_hd__o22ai_1 _26400_ (.A1(net131),
    .A2(_00366_),
    .B1(_03445_),
    .B2(_03447_),
    .Y(_03449_));
 sky130_fd_sc_hd__o2111ai_1 _26401_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_03446_),
    .D1(_03448_),
    .Y(_03450_));
 sky130_fd_sc_hd__o211ai_1 _26402_ (.A1(net131),
    .A2(_00366_),
    .B1(_03446_),
    .C1(_03448_),
    .Y(_03451_));
 sky130_fd_sc_hd__o21ai_1 _26403_ (.A1(_03445_),
    .A2(_03447_),
    .B1(_00736_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand3_1 _26404_ (.A(_03453_),
    .B(_03409_),
    .C(_03451_),
    .Y(_03454_));
 sky130_fd_sc_hd__nand3_2 _26405_ (.A(_03410_),
    .B(_03449_),
    .C(_03450_),
    .Y(_03455_));
 sky130_fd_sc_hd__a21oi_2 _26406_ (.A1(_03454_),
    .A2(_03455_),
    .B1(_02948_),
    .Y(_03456_));
 sky130_fd_sc_hd__o2111a_1 _26407_ (.A1(_02944_),
    .A2(_02706_),
    .B1(_02712_),
    .C1(_03454_),
    .D1(_03455_),
    .X(_03457_));
 sky130_fd_sc_hd__nand3_1 _26408_ (.A(_03454_),
    .B(_03455_),
    .C(_02948_),
    .Y(_03458_));
 sky130_fd_sc_hd__o21ai_1 _26409_ (.A1(_02949_),
    .A2(_03326_),
    .B1(_03329_),
    .Y(_03459_));
 sky130_fd_sc_hd__a21oi_2 _26410_ (.A1(_03327_),
    .A2(_02948_),
    .B1(_03328_),
    .Y(_03460_));
 sky130_fd_sc_hd__o21ai_4 _26411_ (.A1(_03456_),
    .A2(_03457_),
    .B1(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__inv_2 _26412_ (.A(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand3b_2 _26413_ (.A_N(_03456_),
    .B(_03458_),
    .C(_03459_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_1 _26414_ (.A(_03461_),
    .B(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__nand3_1 _26415_ (.A(_03407_),
    .B(_03461_),
    .C(_03464_),
    .Y(_03466_));
 sky130_fd_sc_hd__a21o_1 _26416_ (.A1(_03461_),
    .A2(_03464_),
    .B1(_03407_),
    .X(_03467_));
 sky130_fd_sc_hd__o2111a_1 _26417_ (.A1(_03406_),
    .A2(_03402_),
    .B1(_03405_),
    .C1(_03461_),
    .D1(_03464_),
    .X(_03468_));
 sky130_fd_sc_hd__nand2_1 _26418_ (.A(_03465_),
    .B(_03407_),
    .Y(_03469_));
 sky130_fd_sc_hd__nand3b_1 _26419_ (.A_N(_03468_),
    .B(_03469_),
    .C(_03364_),
    .Y(_03470_));
 sky130_fd_sc_hd__o2111ai_2 _26420_ (.A1(_03280_),
    .A2(_03336_),
    .B1(_03338_),
    .C1(_03466_),
    .D1(_03467_),
    .Y(_03471_));
 sky130_fd_sc_hd__a31o_1 _26421_ (.A1(_03064_),
    .A2(_03272_),
    .A3(_03276_),
    .B1(_03274_),
    .X(_03472_));
 sky130_fd_sc_hd__a22o_1 _26422_ (.A1(_03273_),
    .A2(_03278_),
    .B1(_03470_),
    .B2(_03471_),
    .X(_03473_));
 sky130_fd_sc_hd__nand4_1 _26423_ (.A(_03273_),
    .B(_03278_),
    .C(_03470_),
    .D(_03471_),
    .Y(_03475_));
 sky130_fd_sc_hd__a21o_1 _26424_ (.A1(_03473_),
    .A2(_03475_),
    .B1(_03362_),
    .X(_03476_));
 sky130_fd_sc_hd__nand3_1 _26425_ (.A(_03362_),
    .B(_03473_),
    .C(_03475_),
    .Y(_03477_));
 sky130_fd_sc_hd__a21o_1 _26426_ (.A1(_03476_),
    .A2(_03477_),
    .B1(_03360_),
    .X(_03478_));
 sky130_fd_sc_hd__nand3_1 _26427_ (.A(_03360_),
    .B(_03476_),
    .C(_03477_),
    .Y(_03479_));
 sky130_fd_sc_hd__a21oi_1 _26428_ (.A1(_03478_),
    .A2(_03479_),
    .B1(_03359_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand3_1 _26429_ (.A(_03359_),
    .B(_03478_),
    .C(_03479_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand2b_2 _26430_ (.A_N(_03480_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__a21boi_2 _26431_ (.A1(_03356_),
    .A2(_03192_),
    .B1_N(_03355_),
    .Y(_03483_));
 sky130_fd_sc_hd__nand3_1 _26432_ (.A(_03193_),
    .B(_03355_),
    .C(_03356_),
    .Y(_03484_));
 sky130_fd_sc_hd__inv_2 _26433_ (.A(_03484_),
    .Y(_03486_));
 sky130_fd_sc_hd__a21boi_1 _26434_ (.A1(_03202_),
    .A2(_03486_),
    .B1_N(_03483_),
    .Y(_03487_));
 sky130_fd_sc_hd__xor2_1 _26435_ (.A(_03482_),
    .B(_03487_),
    .X(net118));
 sky130_fd_sc_hd__a21bo_1 _26436_ (.A1(_03360_),
    .A2(_03477_),
    .B1_N(_03476_),
    .X(_03488_));
 sky130_fd_sc_hd__a21bo_1 _26437_ (.A1(_03367_),
    .A2(_03393_),
    .B1_N(_03394_),
    .X(_03489_));
 sky130_fd_sc_hd__nand2_1 _26438_ (.A(_03455_),
    .B(_03458_),
    .Y(_03490_));
 sky130_fd_sc_hd__a21oi_1 _26439_ (.A1(_03426_),
    .A2(_10545_),
    .B1(_03424_),
    .Y(_03491_));
 sky130_fd_sc_hd__a21o_1 _26440_ (.A1(_03426_),
    .A2(_10545_),
    .B1(_03424_),
    .X(_03492_));
 sky130_fd_sc_hd__a21oi_1 _26441_ (.A1(net144),
    .A2(_03418_),
    .B1(_03415_),
    .Y(_03493_));
 sky130_fd_sc_hd__o21ai_2 _26442_ (.A1(_09299_),
    .A2(_03417_),
    .B1(_03416_),
    .Y(_03494_));
 sky130_fd_sc_hd__or3_1 _26443_ (.A(net57),
    .B(_04266_),
    .C(_04223_),
    .X(_03496_));
 sky130_fd_sc_hd__nand3_2 _26444_ (.A(_07499_),
    .B(_07503_),
    .C(_08657_),
    .Y(_03497_));
 sky130_fd_sc_hd__o311a_2 _26445_ (.A1(_08658_),
    .A2(_07502_),
    .A3(_07498_),
    .B1(_03496_),
    .C1(_08878_),
    .X(_03498_));
 sky130_fd_sc_hd__o221ai_4 _26446_ (.A1(_04223_),
    .A2(_08660_),
    .B1(net153),
    .B2(_03286_),
    .C1(_03497_),
    .Y(_03499_));
 sky130_fd_sc_hd__a21oi_1 _26447_ (.A1(_03496_),
    .A2(_03497_),
    .B1(net149),
    .Y(_03500_));
 sky130_fd_sc_hd__a21o_2 _26448_ (.A1(_03496_),
    .A2(_03497_),
    .B1(net149),
    .X(_03501_));
 sky130_fd_sc_hd__o211ai_4 _26449_ (.A1(net237),
    .A2(_09297_),
    .B1(_03499_),
    .C1(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__o21ai_2 _26450_ (.A1(_03498_),
    .A2(_03500_),
    .B1(_09299_),
    .Y(_03503_));
 sky130_fd_sc_hd__o22ai_2 _26451_ (.A1(net237),
    .A2(_09297_),
    .B1(_03498_),
    .B2(_03500_),
    .Y(_03504_));
 sky130_fd_sc_hd__nand3_1 _26452_ (.A(_03501_),
    .B(_09299_),
    .C(_03499_),
    .Y(_03505_));
 sky130_fd_sc_hd__a21oi_1 _26453_ (.A1(_03504_),
    .A2(_03505_),
    .B1(_03493_),
    .Y(_03508_));
 sky130_fd_sc_hd__nand3_4 _26454_ (.A(_03494_),
    .B(_03502_),
    .C(_03503_),
    .Y(_03509_));
 sky130_fd_sc_hd__nand3_2 _26455_ (.A(_03493_),
    .B(_03504_),
    .C(_03505_),
    .Y(_03510_));
 sky130_fd_sc_hd__nand3_1 _26456_ (.A(_03503_),
    .B(_03493_),
    .C(_03502_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand3_1 _26457_ (.A(_03494_),
    .B(_03504_),
    .C(_03505_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand3_4 _26458_ (.A(_03509_),
    .B(_03510_),
    .C(_10545_),
    .Y(_03513_));
 sky130_fd_sc_hd__o211ai_4 _26459_ (.A1(net140),
    .A2(_10542_),
    .B1(_03511_),
    .C1(_03512_),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2_1 _26460_ (.A(_03513_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__a21oi_2 _26461_ (.A1(_03513_),
    .A2(_03514_),
    .B1(_03492_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_2 _26462_ (.A(_03515_),
    .B(_03491_),
    .Y(_03517_));
 sky130_fd_sc_hd__and3_1 _26463_ (.A(_03492_),
    .B(_03513_),
    .C(_03514_),
    .X(_03519_));
 sky130_fd_sc_hd__nand3_4 _26464_ (.A(_03492_),
    .B(_03513_),
    .C(_03514_),
    .Y(_03520_));
 sky130_fd_sc_hd__a21o_1 _26465_ (.A1(_03517_),
    .A2(_03520_),
    .B1(_12099_),
    .X(_03521_));
 sky130_fd_sc_hd__a22o_2 _26466_ (.A1(net143),
    .A2(_11743_),
    .B1(_03515_),
    .B2(_03491_),
    .X(_03522_));
 sky130_fd_sc_hd__o2bb2ai_4 _26467_ (.A1_N(_03517_),
    .A2_N(_03520_),
    .B1(net141),
    .B2(_11742_),
    .Y(_03523_));
 sky130_fd_sc_hd__o2111ai_4 _26468_ (.A1(_11737_),
    .A2(_11740_),
    .B1(_03520_),
    .C1(net143),
    .D1(_03517_),
    .Y(_03524_));
 sky130_fd_sc_hd__a22oi_4 _26469_ (.A1(_03437_),
    .A2(_03443_),
    .B1(_03523_),
    .B2(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__o221ai_4 _26470_ (.A1(_03519_),
    .A2(_03522_),
    .B1(_03436_),
    .B2(_03442_),
    .C1(_03521_),
    .Y(_03526_));
 sky130_fd_sc_hd__o2111a_1 _26471_ (.A1(_12098_),
    .A2(_03434_),
    .B1(_03437_),
    .C1(_03523_),
    .D1(_03524_),
    .X(_03527_));
 sky130_fd_sc_hd__o2111ai_4 _26472_ (.A1(_12098_),
    .A2(_03434_),
    .B1(_03437_),
    .C1(_03523_),
    .D1(_03524_),
    .Y(_03528_));
 sky130_fd_sc_hd__o22ai_2 _26473_ (.A1(net131),
    .A2(_00366_),
    .B1(_03525_),
    .B2(_03527_),
    .Y(_03530_));
 sky130_fd_sc_hd__a41oi_2 _26474_ (.A1(_03437_),
    .A2(_03443_),
    .A3(_03523_),
    .A4(_03524_),
    .B1(net129),
    .Y(_03531_));
 sky130_fd_sc_hd__o2111ai_4 _26475_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_03526_),
    .D1(_03528_),
    .Y(_03532_));
 sky130_fd_sc_hd__o21ai_2 _26476_ (.A1(net129),
    .A2(_03447_),
    .B1(_03446_),
    .Y(_03533_));
 sky130_fd_sc_hd__a21oi_1 _26477_ (.A1(_03530_),
    .A2(_03532_),
    .B1(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__a21o_1 _26478_ (.A1(_03530_),
    .A2(_03532_),
    .B1(_03533_),
    .X(_03535_));
 sky130_fd_sc_hd__and3_1 _26479_ (.A(_03530_),
    .B(_03533_),
    .C(_03532_),
    .X(_03536_));
 sky130_fd_sc_hd__nand3_1 _26480_ (.A(_03530_),
    .B(_03533_),
    .C(_03532_),
    .Y(_03537_));
 sky130_fd_sc_hd__o22ai_1 _26481_ (.A1(_02711_),
    .A2(_02945_),
    .B1(_03534_),
    .B2(_03536_),
    .Y(_03538_));
 sky130_fd_sc_hd__o211a_1 _26482_ (.A1(_02944_),
    .A2(_02706_),
    .B1(_02712_),
    .C1(_03535_),
    .X(_03539_));
 sky130_fd_sc_hd__nand3_1 _26483_ (.A(_03535_),
    .B(_03537_),
    .C(_02948_),
    .Y(_03541_));
 sky130_fd_sc_hd__a21o_1 _26484_ (.A1(_03538_),
    .A2(_03541_),
    .B1(_03490_),
    .X(_03542_));
 sky130_fd_sc_hd__nand3_1 _26485_ (.A(_03490_),
    .B(_03538_),
    .C(_03541_),
    .Y(_03543_));
 sky130_fd_sc_hd__a31o_1 _26486_ (.A1(_03240_),
    .A2(_03255_),
    .A3(_03256_),
    .B1(_03399_),
    .X(_03544_));
 sky130_fd_sc_hd__o311a_1 _26487_ (.A1(net233),
    .A2(_05927_),
    .A3(_07767_),
    .B1(_07771_),
    .C1(net238),
    .X(_03545_));
 sky130_fd_sc_hd__and3_1 _26488_ (.A(_04266_),
    .B(net54),
    .C(net22),
    .X(_03546_));
 sky130_fd_sc_hd__a31o_1 _26489_ (.A1(net166),
    .A2(_07771_),
    .A3(net238),
    .B1(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__o311a_1 _26490_ (.A1(_05931_),
    .A2(_07074_),
    .A3(net268),
    .B1(_07642_),
    .C1(_08204_),
    .X(_03548_));
 sky130_fd_sc_hd__and3b_1 _26491_ (.A_N(net54),
    .B(net24),
    .C(net53),
    .X(_03549_));
 sky130_fd_sc_hd__a21oi_1 _26492_ (.A1(net24),
    .A2(_07643_),
    .B1(_03548_),
    .Y(_03550_));
 sky130_fd_sc_hd__a31o_1 _26493_ (.A1(_08204_),
    .A2(net163),
    .A3(_07642_),
    .B1(_03549_),
    .X(_03552_));
 sky130_fd_sc_hd__or3b_4 _26494_ (.A(net53),
    .B(net319),
    .C_N(net52),
    .X(_03553_));
 sky130_fd_sc_hd__a21oi_1 _26495_ (.A1(net153),
    .A2(net158),
    .B1(_07306_),
    .Y(_03554_));
 sky130_fd_sc_hd__o21ai_1 _26496_ (.A1(net160),
    .A2(_08666_),
    .B1(net239),
    .Y(_03555_));
 sky130_fd_sc_hd__a31oi_4 _26497_ (.A1(net319),
    .A2(net163),
    .A3(net269),
    .B1(_03376_),
    .Y(_03556_));
 sky130_fd_sc_hd__o221ai_2 _26498_ (.A1(net319),
    .A2(_06866_),
    .B1(net153),
    .B2(_06864_),
    .C1(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__a22o_1 _26499_ (.A1(_03375_),
    .A2(_03556_),
    .B1(_03555_),
    .B2(_03553_),
    .X(_03558_));
 sky130_fd_sc_hd__o2111ai_4 _26500_ (.A1(_07306_),
    .A2(_08669_),
    .B1(_03375_),
    .C1(_03553_),
    .D1(_03556_),
    .Y(_03559_));
 sky130_fd_sc_hd__nand2_1 _26501_ (.A(_03558_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__a221oi_4 _26502_ (.A1(_03372_),
    .A2(_03378_),
    .B1(_03558_),
    .B2(_03559_),
    .C1(_03379_),
    .Y(_03561_));
 sky130_fd_sc_hd__a221o_1 _26503_ (.A1(_03372_),
    .A2(_03378_),
    .B1(_03558_),
    .B2(_03559_),
    .C1(_03379_),
    .X(_03563_));
 sky130_fd_sc_hd__a21oi_1 _26504_ (.A1(_03380_),
    .A2(_03381_),
    .B1(_03560_),
    .Y(_03564_));
 sky130_fd_sc_hd__a21o_1 _26505_ (.A1(_03380_),
    .A2(_03381_),
    .B1(_03560_),
    .X(_03565_));
 sky130_fd_sc_hd__o22a_1 _26506_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_03561_),
    .B2(_03564_),
    .X(_03566_));
 sky130_fd_sc_hd__o21ai_1 _26507_ (.A1(_03561_),
    .A2(_03564_),
    .B1(_03552_),
    .Y(_03567_));
 sky130_fd_sc_hd__nor4_1 _26508_ (.A(_03548_),
    .B(_03549_),
    .C(_03561_),
    .D(_03564_),
    .Y(_03568_));
 sky130_fd_sc_hd__nand3_1 _26509_ (.A(_03563_),
    .B(_03565_),
    .C(_03550_),
    .Y(_03569_));
 sky130_fd_sc_hd__o2bb2ai_2 _26510_ (.A1_N(_03386_),
    .A2_N(_03390_),
    .B1(_03566_),
    .B2(_03568_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand4_2 _26511_ (.A(_03386_),
    .B(_03390_),
    .C(_03567_),
    .D(_03569_),
    .Y(_03571_));
 sky130_fd_sc_hd__o211a_1 _26512_ (.A1(_03545_),
    .A2(_03546_),
    .B1(_03570_),
    .C1(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__o211ai_2 _26513_ (.A1(_03545_),
    .A2(_03546_),
    .B1(_03570_),
    .C1(_03571_),
    .Y(_03574_));
 sky130_fd_sc_hd__a21oi_1 _26514_ (.A1(_03570_),
    .A2(_03571_),
    .B1(_03547_),
    .Y(_03575_));
 sky130_fd_sc_hd__a21o_1 _26515_ (.A1(_03570_),
    .A2(_03571_),
    .B1(_03547_),
    .X(_03576_));
 sky130_fd_sc_hd__o22ai_2 _26516_ (.A1(_03263_),
    .A2(_03265_),
    .B1(_03572_),
    .B2(_03575_),
    .Y(_03577_));
 sky130_fd_sc_hd__nand3b_2 _26517_ (.A_N(_03267_),
    .B(_03574_),
    .C(_03576_),
    .Y(_03578_));
 sky130_fd_sc_hd__a32o_1 _26518_ (.A1(_11740_),
    .A2(_00361_),
    .A3(_02709_),
    .B1(_03577_),
    .B2(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__o2111ai_4 _26519_ (.A1(_02706_),
    .A2(_01332_),
    .B1(net131),
    .C1(_03578_),
    .D1(_03577_),
    .Y(_03580_));
 sky130_fd_sc_hd__inv_2 _26520_ (.A(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__a21o_1 _26521_ (.A1(_03579_),
    .A2(_03580_),
    .B1(_03544_),
    .X(_03582_));
 sky130_fd_sc_hd__nand2_1 _26522_ (.A(_03544_),
    .B(_03579_),
    .Y(_03583_));
 sky130_fd_sc_hd__o21a_1 _26523_ (.A1(_03581_),
    .A2(_03583_),
    .B1(_03582_),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_1 _26524_ (.A1(_03542_),
    .A2(_03543_),
    .B1(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__o2111ai_2 _26525_ (.A1(_03581_),
    .A2(_03583_),
    .B1(_03582_),
    .C1(_03542_),
    .D1(_03543_),
    .Y(_03587_));
 sky130_fd_sc_hd__o31a_1 _26526_ (.A1(_03456_),
    .A2(_03457_),
    .A3(_03460_),
    .B1(_03407_),
    .X(_03588_));
 sky130_fd_sc_hd__nand2_1 _26527_ (.A(_03407_),
    .B(_03464_),
    .Y(_03589_));
 sky130_fd_sc_hd__o2bb2ai_1 _26528_ (.A1_N(_03586_),
    .A2_N(_03587_),
    .B1(_03588_),
    .B2(_03462_),
    .Y(_03590_));
 sky130_fd_sc_hd__nand4_2 _26529_ (.A(_03461_),
    .B(_03586_),
    .C(_03587_),
    .D(_03589_),
    .Y(_03591_));
 sky130_fd_sc_hd__o21bai_1 _26530_ (.A1(_03404_),
    .A2(_03402_),
    .B1_N(_03401_),
    .Y(_03592_));
 sky130_fd_sc_hd__a21oi_1 _26531_ (.A1(_03590_),
    .A2(_03591_),
    .B1(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_1 _26532_ (.A(_03590_),
    .B(_03592_),
    .Y(_03594_));
 sky130_fd_sc_hd__and3_1 _26533_ (.A(_03590_),
    .B(_03591_),
    .C(_03592_),
    .X(_03596_));
 sky130_fd_sc_hd__a21boi_1 _26534_ (.A1(_03471_),
    .A2(_03472_),
    .B1_N(_03470_),
    .Y(_03597_));
 sky130_fd_sc_hd__o21a_1 _26535_ (.A1(_03593_),
    .A2(_03596_),
    .B1(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__o21ai_1 _26536_ (.A1(_03593_),
    .A2(_03596_),
    .B1(_03597_),
    .Y(_03599_));
 sky130_fd_sc_hd__nor3_1 _26537_ (.A(_03593_),
    .B(_03597_),
    .C(_03596_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21o_1 _26538_ (.A1(_03599_),
    .A2(_03489_),
    .B1(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__o21bai_1 _26539_ (.A1(_03598_),
    .A2(_03600_),
    .B1_N(_03489_),
    .Y(_03602_));
 sky130_fd_sc_hd__nand3b_1 _26540_ (.A_N(_03600_),
    .B(_03489_),
    .C(_03599_),
    .Y(_03603_));
 sky130_fd_sc_hd__a21oi_1 _26541_ (.A1(_03602_),
    .A2(_03603_),
    .B1(_03488_),
    .Y(_03604_));
 sky130_fd_sc_hd__nand3_1 _26542_ (.A(_03488_),
    .B(_03602_),
    .C(_03603_),
    .Y(_03605_));
 sky130_fd_sc_hd__nand2b_2 _26543_ (.A_N(_03604_),
    .B(_03605_),
    .Y(_03607_));
 sky130_fd_sc_hd__a21oi_1 _26544_ (.A1(_03487_),
    .A2(_03481_),
    .B1(_03480_),
    .Y(_03608_));
 sky130_fd_sc_hd__xnor2_1 _26545_ (.A(_03607_),
    .B(_03608_),
    .Y(net119));
 sky130_fd_sc_hd__nand2_1 _26546_ (.A(_03570_),
    .B(_03574_),
    .Y(_03609_));
 sky130_fd_sc_hd__a21bo_1 _26547_ (.A1(_03585_),
    .A2(_03542_),
    .B1_N(_03543_),
    .X(_03610_));
 sky130_fd_sc_hd__a21oi_1 _26548_ (.A1(_03528_),
    .A2(_00736_),
    .B1(_03525_),
    .Y(_03611_));
 sky130_fd_sc_hd__a21o_1 _26549_ (.A1(_10545_),
    .A2(_03510_),
    .B1(_03508_),
    .X(_03612_));
 sky130_fd_sc_hd__o21ai_1 _26550_ (.A1(_09299_),
    .A2(_03498_),
    .B1(_03501_),
    .Y(_03613_));
 sky130_fd_sc_hd__or3_1 _26551_ (.A(net57),
    .B(_04266_),
    .C(_04245_),
    .X(_03614_));
 sky130_fd_sc_hd__o211ai_4 _26552_ (.A1(net170),
    .A2(_07765_),
    .B1(_08657_),
    .C1(_07771_),
    .Y(_03615_));
 sky130_fd_sc_hd__o311a_1 _26553_ (.A1(_04245_),
    .A2(_04266_),
    .A3(net57),
    .B1(_08878_),
    .C1(_03615_),
    .X(_03618_));
 sky130_fd_sc_hd__o221ai_4 _26554_ (.A1(_04245_),
    .A2(_08660_),
    .B1(net152),
    .B2(_03286_),
    .C1(_03615_),
    .Y(_03619_));
 sky130_fd_sc_hd__a21oi_1 _26555_ (.A1(_03614_),
    .A2(_03615_),
    .B1(_08878_),
    .Y(_03620_));
 sky130_fd_sc_hd__a21o_1 _26556_ (.A1(_03614_),
    .A2(_03615_),
    .B1(_08878_),
    .X(_03621_));
 sky130_fd_sc_hd__o211ai_2 _26557_ (.A1(net237),
    .A2(_09297_),
    .B1(_03619_),
    .C1(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__o21ai_1 _26558_ (.A1(_03618_),
    .A2(_03620_),
    .B1(_09299_),
    .Y(_03623_));
 sky130_fd_sc_hd__o22ai_2 _26559_ (.A1(net237),
    .A2(_09297_),
    .B1(_03618_),
    .B2(_03620_),
    .Y(_03624_));
 sky130_fd_sc_hd__o2111ai_4 _26560_ (.A1(_04495_),
    .A2(net152),
    .B1(_08882_),
    .C1(_03619_),
    .D1(_03621_),
    .Y(_03625_));
 sky130_fd_sc_hd__a22oi_2 _26561_ (.A1(_03501_),
    .A2(_03502_),
    .B1(_03624_),
    .B2(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand3_1 _26562_ (.A(_03613_),
    .B(_03622_),
    .C(_03623_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand4_2 _26563_ (.A(_03501_),
    .B(_03502_),
    .C(_03624_),
    .D(_03625_),
    .Y(_03629_));
 sky130_fd_sc_hd__o2111ai_2 _26564_ (.A1(_09299_),
    .A2(_03498_),
    .B1(_03501_),
    .C1(_03622_),
    .D1(_03623_),
    .Y(_03630_));
 sky130_fd_sc_hd__nand3_1 _26565_ (.A(_03613_),
    .B(_03624_),
    .C(_03625_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand4_1 _26566_ (.A(net139),
    .B(_10544_),
    .C(_03627_),
    .D(_03629_),
    .Y(_03632_));
 sky130_fd_sc_hd__o211ai_1 _26567_ (.A1(net140),
    .A2(_10542_),
    .B1(_03630_),
    .C1(_03631_),
    .Y(_03633_));
 sky130_fd_sc_hd__o211ai_2 _26568_ (.A1(net140),
    .A2(_10542_),
    .B1(_03627_),
    .C1(_03629_),
    .Y(_03634_));
 sky130_fd_sc_hd__nand3_2 _26569_ (.A(_03630_),
    .B(_03631_),
    .C(_10545_),
    .Y(_03635_));
 sky130_fd_sc_hd__nand4_4 _26570_ (.A(_03509_),
    .B(_03513_),
    .C(_03634_),
    .D(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__nand3_2 _26571_ (.A(_03612_),
    .B(_03632_),
    .C(_03633_),
    .Y(_03637_));
 sky130_fd_sc_hd__a41o_1 _26572_ (.A1(_03509_),
    .A2(_03513_),
    .A3(_03634_),
    .A4(_03635_),
    .B1(_12098_),
    .X(_03638_));
 sky130_fd_sc_hd__o2bb2ai_4 _26573_ (.A1_N(_03636_),
    .A2_N(_03637_),
    .B1(net141),
    .B2(_11742_),
    .Y(_03640_));
 sky130_fd_sc_hd__o2111ai_4 _26574_ (.A1(_11737_),
    .A2(_11740_),
    .B1(net143),
    .C1(_03636_),
    .D1(_03637_),
    .Y(_03641_));
 sky130_fd_sc_hd__a31oi_1 _26575_ (.A1(_03492_),
    .A2(_03513_),
    .A3(_03514_),
    .B1(_12099_),
    .Y(_03642_));
 sky130_fd_sc_hd__o211a_1 _26576_ (.A1(_03516_),
    .A2(_03642_),
    .B1(_03641_),
    .C1(_03640_),
    .X(_03643_));
 sky130_fd_sc_hd__o2111ai_4 _26577_ (.A1(_12098_),
    .A2(_03516_),
    .B1(_03520_),
    .C1(_03640_),
    .D1(_03641_),
    .Y(_03644_));
 sky130_fd_sc_hd__a22oi_4 _26578_ (.A1(_03520_),
    .A2(_03522_),
    .B1(_03640_),
    .B2(_03641_),
    .Y(_03645_));
 sky130_fd_sc_hd__a22o_1 _26579_ (.A1(_03520_),
    .A2(_03522_),
    .B1(_03640_),
    .B2(_03641_),
    .X(_03646_));
 sky130_fd_sc_hd__o22ai_1 _26580_ (.A1(net131),
    .A2(_00366_),
    .B1(_03643_),
    .B2(_03645_),
    .Y(_03647_));
 sky130_fd_sc_hd__o2111ai_1 _26581_ (.A1(_00365_),
    .A2(_00357_),
    .B1(_00364_),
    .C1(_03644_),
    .D1(_03646_),
    .Y(_03648_));
 sky130_fd_sc_hd__o21ai_1 _26582_ (.A1(_03643_),
    .A2(_03645_),
    .B1(_00736_),
    .Y(_03649_));
 sky130_fd_sc_hd__o211ai_1 _26583_ (.A1(net131),
    .A2(_00366_),
    .B1(_03644_),
    .C1(_03646_),
    .Y(_03651_));
 sky130_fd_sc_hd__o211ai_2 _26584_ (.A1(_03525_),
    .A2(_03531_),
    .B1(_03647_),
    .C1(_03648_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand3_1 _26585_ (.A(_03611_),
    .B(_03649_),
    .C(_03651_),
    .Y(_03653_));
 sky130_fd_sc_hd__o2111a_1 _26586_ (.A1(_02944_),
    .A2(_02706_),
    .B1(_02712_),
    .C1(_03652_),
    .D1(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__a21oi_1 _26587_ (.A1(_03652_),
    .A2(_03653_),
    .B1(_02948_),
    .Y(_03655_));
 sky130_fd_sc_hd__nor2_1 _26588_ (.A(_03654_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__o21ai_1 _26589_ (.A1(_03536_),
    .A2(_03539_),
    .B1(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__o211ai_2 _26590_ (.A1(_03654_),
    .A2(_03655_),
    .B1(_03537_),
    .C1(_03541_),
    .Y(_03658_));
 sky130_fd_sc_hd__a31o_1 _26591_ (.A1(_03266_),
    .A2(_03574_),
    .A3(_03576_),
    .B1(_03263_),
    .X(_03659_));
 sky130_fd_sc_hd__a32o_1 _26592_ (.A1(_08204_),
    .A2(net163),
    .A3(net238),
    .B1(_08006_),
    .B2(net24),
    .X(_03660_));
 sky130_fd_sc_hd__a22o_1 _26593_ (.A1(net25),
    .A2(_07643_),
    .B1(_08670_),
    .B2(_07642_),
    .X(_03661_));
 sky130_fd_sc_hd__o31a_1 _26594_ (.A1(net25),
    .A2(_07306_),
    .A3(_08207_),
    .B1(_03553_),
    .X(_03662_));
 sky130_fd_sc_hd__nand3_2 _26595_ (.A(_03375_),
    .B(_03556_),
    .C(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__o2111a_1 _26596_ (.A1(_07306_),
    .A2(net153),
    .B1(_03553_),
    .C1(_03554_),
    .D1(_03557_),
    .X(_03664_));
 sky130_fd_sc_hd__o2111ai_2 _26597_ (.A1(_07306_),
    .A2(net153),
    .B1(_03553_),
    .C1(_03554_),
    .D1(_03557_),
    .Y(_03665_));
 sky130_fd_sc_hd__a21o_1 _26598_ (.A1(_03663_),
    .A2(_03665_),
    .B1(_03661_),
    .X(_03666_));
 sky130_fd_sc_hd__nand2_1 _26599_ (.A(_03661_),
    .B(_03663_),
    .Y(_03667_));
 sky130_fd_sc_hd__o21a_1 _26600_ (.A1(_03664_),
    .A2(_03667_),
    .B1(_03666_),
    .X(_03668_));
 sky130_fd_sc_hd__o21ai_1 _26601_ (.A1(_03550_),
    .A2(_03561_),
    .B1(_03565_),
    .Y(_03669_));
 sky130_fd_sc_hd__a211o_1 _26602_ (.A1(_03552_),
    .A2(_03563_),
    .B1(_03564_),
    .C1(_03668_),
    .X(_03670_));
 sky130_fd_sc_hd__nand2_1 _26603_ (.A(_03669_),
    .B(_03668_),
    .Y(_03672_));
 sky130_fd_sc_hd__and3_1 _26604_ (.A(_03660_),
    .B(_03670_),
    .C(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__nand3_2 _26605_ (.A(_03660_),
    .B(_03670_),
    .C(_03672_),
    .Y(_03674_));
 sky130_fd_sc_hd__a21o_1 _26606_ (.A1(_03670_),
    .A2(_03672_),
    .B1(_03660_),
    .X(_03675_));
 sky130_fd_sc_hd__a211o_1 _26607_ (.A1(_03674_),
    .A2(_03675_),
    .B1(_02699_),
    .C1(_03260_),
    .X(_03676_));
 sky130_fd_sc_hd__o211ai_4 _26608_ (.A1(_02699_),
    .A2(_03260_),
    .B1(_03674_),
    .C1(_03675_),
    .Y(_03677_));
 sky130_fd_sc_hd__o2111ai_2 _26609_ (.A1(_01332_),
    .A2(_02706_),
    .B1(_03677_),
    .C1(net131),
    .D1(_03676_),
    .Y(_03678_));
 sky130_fd_sc_hd__a32o_1 _26610_ (.A1(_11740_),
    .A2(_00361_),
    .A3(_02709_),
    .B1(_03676_),
    .B2(_03677_),
    .X(_03679_));
 sky130_fd_sc_hd__a21o_1 _26611_ (.A1(_03678_),
    .A2(_03679_),
    .B1(_03659_),
    .X(_03680_));
 sky130_fd_sc_hd__nand3_1 _26612_ (.A(_03659_),
    .B(_03678_),
    .C(_03679_),
    .Y(_03681_));
 sky130_fd_sc_hd__nand2_1 _26613_ (.A(_03680_),
    .B(_03681_),
    .Y(_03683_));
 sky130_fd_sc_hd__a22o_1 _26614_ (.A1(_03657_),
    .A2(_03658_),
    .B1(_03680_),
    .B2(_03681_),
    .X(_03684_));
 sky130_fd_sc_hd__nand3b_1 _26615_ (.A_N(_03683_),
    .B(_03658_),
    .C(_03657_),
    .Y(_03685_));
 sky130_fd_sc_hd__a21oi_1 _26616_ (.A1(_03684_),
    .A2(_03685_),
    .B1(_03610_),
    .Y(_03686_));
 sky130_fd_sc_hd__and3_1 _26617_ (.A(_03610_),
    .B(_03684_),
    .C(_03685_),
    .X(_03687_));
 sky130_fd_sc_hd__a21oi_1 _26618_ (.A1(_03544_),
    .A2(_03579_),
    .B1(_03581_),
    .Y(_03688_));
 sky130_fd_sc_hd__o211a_1 _26619_ (.A1(_03686_),
    .A2(_03687_),
    .B1(_03580_),
    .C1(_03583_),
    .X(_03689_));
 sky130_fd_sc_hd__a211oi_1 _26620_ (.A1(_03580_),
    .A2(_03583_),
    .B1(_03686_),
    .C1(_03687_),
    .Y(_03690_));
 sky130_fd_sc_hd__o211ai_2 _26621_ (.A1(_03689_),
    .A2(_03690_),
    .B1(_03591_),
    .C1(_03594_),
    .Y(_03691_));
 sky130_fd_sc_hd__a211o_1 _26622_ (.A1(_03591_),
    .A2(_03594_),
    .B1(_03689_),
    .C1(_03690_),
    .X(_03692_));
 sky130_fd_sc_hd__a21o_1 _26623_ (.A1(_03691_),
    .A2(_03692_),
    .B1(_03609_),
    .X(_03694_));
 sky130_fd_sc_hd__nand3_1 _26624_ (.A(_03609_),
    .B(_03691_),
    .C(_03692_),
    .Y(_03695_));
 sky130_fd_sc_hd__and2_1 _26625_ (.A(_03694_),
    .B(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__nand2_1 _26626_ (.A(_03601_),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__a221o_1 _26627_ (.A1(_03489_),
    .A2(_03599_),
    .B1(_03694_),
    .B2(_03695_),
    .C1(_03600_),
    .X(_03698_));
 sky130_fd_sc_hd__inv_2 _26628_ (.A(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__and4bb_1 _26629_ (.A_N(_03480_),
    .B_N(_03607_),
    .C(_03481_),
    .D(_03486_),
    .X(_03700_));
 sky130_fd_sc_hd__or3_1 _26630_ (.A(_03482_),
    .B(_03484_),
    .C(_03607_),
    .X(_03701_));
 sky130_fd_sc_hd__a21oi_2 _26631_ (.A1(_03197_),
    .A2(_03201_),
    .B1(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__o21a_1 _26632_ (.A1(_03481_),
    .A2(_03604_),
    .B1(_03605_),
    .X(_03703_));
 sky130_fd_sc_hd__o31ai_4 _26633_ (.A1(_03482_),
    .A2(_03483_),
    .A3(_03607_),
    .B1(_03703_),
    .Y(_03705_));
 sky130_fd_sc_hd__a21oi_2 _26634_ (.A1(_03202_),
    .A2(_03700_),
    .B1(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__o221a_1 _26635_ (.A1(_03601_),
    .A2(_03696_),
    .B1(_03705_),
    .B2(_03702_),
    .C1(_03697_),
    .X(_03707_));
 sky130_fd_sc_hd__nand2_1 _26636_ (.A(_03697_),
    .B(_03698_),
    .Y(_03708_));
 sky130_fd_sc_hd__a21oi_1 _26637_ (.A1(_03706_),
    .A2(_03708_),
    .B1(_03707_),
    .Y(net121));
 sky130_fd_sc_hd__a21boi_1 _26638_ (.A1(_03657_),
    .A2(_03683_),
    .B1_N(_03658_),
    .Y(_03709_));
 sky130_fd_sc_hd__nor2_1 _26639_ (.A(net129),
    .B(_03643_),
    .Y(_03710_));
 sky130_fd_sc_hd__a31o_1 _26640_ (.A1(_00364_),
    .A2(_00367_),
    .A3(_03644_),
    .B1(_03645_),
    .X(_03711_));
 sky130_fd_sc_hd__a21oi_1 _26641_ (.A1(_03629_),
    .A2(_10545_),
    .B1(_03626_),
    .Y(_03712_));
 sky130_fd_sc_hd__a31o_1 _26642_ (.A1(net139),
    .A2(_10544_),
    .A3(_03629_),
    .B1(_03626_),
    .X(_03713_));
 sky130_fd_sc_hd__a21oi_1 _26643_ (.A1(net144),
    .A2(_03619_),
    .B1(_03620_),
    .Y(_03715_));
 sky130_fd_sc_hd__o21ai_1 _26644_ (.A1(_09299_),
    .A2(_03618_),
    .B1(_03621_),
    .Y(_03716_));
 sky130_fd_sc_hd__or3_1 _26645_ (.A(net57),
    .B(_04266_),
    .C(_04256_),
    .X(_03717_));
 sky130_fd_sc_hd__nand3_2 _26646_ (.A(net164),
    .B(net163),
    .C(_08657_),
    .Y(_03718_));
 sky130_fd_sc_hd__o311a_1 _26647_ (.A1(_04256_),
    .A2(_04266_),
    .A3(net57),
    .B1(_08878_),
    .C1(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__o221ai_4 _26648_ (.A1(_04256_),
    .A2(_08660_),
    .B1(net152),
    .B2(_03286_),
    .C1(_03718_),
    .Y(_03720_));
 sky130_fd_sc_hd__a21oi_1 _26649_ (.A1(_03717_),
    .A2(_03718_),
    .B1(_08878_),
    .Y(_03721_));
 sky130_fd_sc_hd__a21o_1 _26650_ (.A1(_03717_),
    .A2(_03718_),
    .B1(_08878_),
    .X(_03722_));
 sky130_fd_sc_hd__o211ai_1 _26651_ (.A1(net237),
    .A2(_09297_),
    .B1(_03720_),
    .C1(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__o21ai_1 _26652_ (.A1(_03719_),
    .A2(_03721_),
    .B1(_09299_),
    .Y(_03724_));
 sky130_fd_sc_hd__o21ai_1 _26653_ (.A1(_03719_),
    .A2(_03721_),
    .B1(net144),
    .Y(_03727_));
 sky130_fd_sc_hd__o2111ai_1 _26654_ (.A1(_04495_),
    .A2(net152),
    .B1(_08882_),
    .C1(_03720_),
    .D1(_03722_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand3_2 _26655_ (.A(_03716_),
    .B(_03723_),
    .C(_03724_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand3_2 _26656_ (.A(_03727_),
    .B(_03728_),
    .C(_03715_),
    .Y(_03730_));
 sky130_fd_sc_hd__nand3_2 _26657_ (.A(_03729_),
    .B(_03730_),
    .C(_10545_),
    .Y(_03731_));
 sky130_fd_sc_hd__a22o_1 _26658_ (.A1(net139),
    .A2(_10544_),
    .B1(_03729_),
    .B2(_03730_),
    .X(_03732_));
 sky130_fd_sc_hd__a21o_1 _26659_ (.A1(_03729_),
    .A2(_03730_),
    .B1(_10546_),
    .X(_03733_));
 sky130_fd_sc_hd__o211ai_1 _26660_ (.A1(net140),
    .A2(_10542_),
    .B1(_03729_),
    .C1(_03730_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand3_2 _26661_ (.A(_03713_),
    .B(_03731_),
    .C(_03732_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand3_2 _26662_ (.A(_03733_),
    .B(_03734_),
    .C(_03712_),
    .Y(_03736_));
 sky130_fd_sc_hd__o211a_1 _26663_ (.A1(_11742_),
    .A2(net141),
    .B1(_03736_),
    .C1(_03735_),
    .X(_03738_));
 sky130_fd_sc_hd__o211ai_2 _26664_ (.A1(_11742_),
    .A2(net141),
    .B1(_03736_),
    .C1(_03735_),
    .Y(_03739_));
 sky130_fd_sc_hd__a21oi_1 _26665_ (.A1(_03735_),
    .A2(_03736_),
    .B1(_12099_),
    .Y(_03740_));
 sky130_fd_sc_hd__a21o_1 _26666_ (.A1(_03735_),
    .A2(_03736_),
    .B1(_12099_),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_1 _26667_ (.A(_03637_),
    .B(_03638_),
    .Y(_03742_));
 sky130_fd_sc_hd__o21bai_2 _26668_ (.A1(_03738_),
    .A2(_03740_),
    .B1_N(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand3_2 _26669_ (.A(_03739_),
    .B(_03741_),
    .C(_03742_),
    .Y(_03744_));
 sky130_fd_sc_hd__a21oi_1 _26670_ (.A1(_03743_),
    .A2(_03744_),
    .B1(_00736_),
    .Y(_03745_));
 sky130_fd_sc_hd__a22o_1 _26671_ (.A1(_00364_),
    .A2(_00367_),
    .B1(_03743_),
    .B2(_03744_),
    .X(_03746_));
 sky130_fd_sc_hd__nand3_2 _26672_ (.A(_03743_),
    .B(_03744_),
    .C(_00736_),
    .Y(_03747_));
 sky130_fd_sc_hd__o21ai_1 _26673_ (.A1(_03645_),
    .A2(_03710_),
    .B1(_03747_),
    .Y(_03749_));
 sky130_fd_sc_hd__nor2_1 _26674_ (.A(_03745_),
    .B(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__o211ai_4 _26675_ (.A1(_03645_),
    .A2(_03710_),
    .B1(_03746_),
    .C1(_03747_),
    .Y(_03751_));
 sky130_fd_sc_hd__a21oi_2 _26676_ (.A1(_03746_),
    .A2(_03747_),
    .B1(_03711_),
    .Y(_03752_));
 sky130_fd_sc_hd__o21ai_1 _26677_ (.A1(_03750_),
    .A2(_03752_),
    .B1(_02949_),
    .Y(_03753_));
 sky130_fd_sc_hd__or3_1 _26678_ (.A(_02711_),
    .B(_02945_),
    .C(_03752_),
    .X(_03754_));
 sky130_fd_sc_hd__nand3b_1 _26679_ (.A_N(_03752_),
    .B(_02948_),
    .C(_03751_),
    .Y(_03755_));
 sky130_fd_sc_hd__a211o_1 _26680_ (.A1(_02712_),
    .A2(_02947_),
    .B1(_03750_),
    .C1(_03752_),
    .X(_03756_));
 sky130_fd_sc_hd__o21ai_1 _26681_ (.A1(_03750_),
    .A2(_03752_),
    .B1(_02948_),
    .Y(_03757_));
 sky130_fd_sc_hd__a32o_1 _26682_ (.A1(_03611_),
    .A2(_03649_),
    .A3(_03651_),
    .B1(_03652_),
    .B2(_02949_),
    .X(_03758_));
 sky130_fd_sc_hd__and3_1 _26683_ (.A(_03756_),
    .B(_03757_),
    .C(_03758_),
    .X(_03760_));
 sky130_fd_sc_hd__nand3_1 _26684_ (.A(_03756_),
    .B(_03757_),
    .C(_03758_),
    .Y(_03761_));
 sky130_fd_sc_hd__nand3b_2 _26685_ (.A_N(_03758_),
    .B(_03755_),
    .C(_03753_),
    .Y(_03762_));
 sky130_fd_sc_hd__o2bb2a_1 _26686_ (.A1_N(net238),
    .A2_N(_08670_),
    .B1(_08007_),
    .B2(net319),
    .X(_03763_));
 sky130_fd_sc_hd__a22oi_1 _26687_ (.A1(net25),
    .A2(_07643_),
    .B1(net160),
    .B2(_07642_),
    .Y(_03764_));
 sky130_fd_sc_hd__a221oi_4 _26688_ (.A1(net25),
    .A2(_07643_),
    .B1(net160),
    .B2(_07642_),
    .C1(_03663_),
    .Y(_03765_));
 sky130_fd_sc_hd__a31oi_2 _26689_ (.A1(_03375_),
    .A2(_03556_),
    .A3(_03662_),
    .B1(_03764_),
    .Y(_03766_));
 sky130_fd_sc_hd__a21oi_1 _26690_ (.A1(_03661_),
    .A2(_03663_),
    .B1(_03664_),
    .Y(_03767_));
 sky130_fd_sc_hd__a211oi_1 _26691_ (.A1(_03665_),
    .A2(_03667_),
    .B1(_03765_),
    .C1(_03766_),
    .Y(_03768_));
 sky130_fd_sc_hd__o21bai_2 _26692_ (.A1(_03766_),
    .A2(_03767_),
    .B1_N(_03765_),
    .Y(_03769_));
 sky130_fd_sc_hd__xnor2_2 _26693_ (.A(_03763_),
    .B(_03769_),
    .Y(_03771_));
 sky130_fd_sc_hd__a41o_1 _26694_ (.A1(_02700_),
    .A2(_02704_),
    .A3(_02857_),
    .A4(_03250_),
    .B1(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__xor2_2 _26695_ (.A(_03265_),
    .B(_03771_),
    .X(_03773_));
 sky130_fd_sc_hd__xor2_2 _26696_ (.A(_02712_),
    .B(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__a31oi_1 _26697_ (.A1(_03266_),
    .A2(_03674_),
    .A3(_03675_),
    .B1(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__and4_1 _26698_ (.A(_03266_),
    .B(_03674_),
    .C(_03675_),
    .D(_03774_),
    .X(_03776_));
 sky130_fd_sc_hd__xnor2_2 _26699_ (.A(_03677_),
    .B(_03774_),
    .Y(_03777_));
 sky130_fd_sc_hd__nand3_1 _26700_ (.A(_03761_),
    .B(_03762_),
    .C(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__o2bb2ai_1 _26701_ (.A1_N(_03761_),
    .A2_N(_03762_),
    .B1(_03775_),
    .B2(_03776_),
    .Y(_03779_));
 sky130_fd_sc_hd__a31o_1 _26702_ (.A1(_03756_),
    .A2(_03757_),
    .A3(_03758_),
    .B1(_03777_),
    .X(_03780_));
 sky130_fd_sc_hd__nand2_1 _26703_ (.A(_03778_),
    .B(_03779_),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _26704_ (.A(_03782_),
    .B(_03709_),
    .Y(_03783_));
 sky130_fd_sc_hd__xor2_1 _26705_ (.A(_03709_),
    .B(_03782_),
    .X(_03784_));
 sky130_fd_sc_hd__a21bo_1 _26706_ (.A1(_03659_),
    .A2(_03679_),
    .B1_N(_03678_),
    .X(_03785_));
 sky130_fd_sc_hd__or2_1 _26707_ (.A(_03784_),
    .B(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__nand2_1 _26708_ (.A(_03784_),
    .B(_03785_),
    .Y(_03787_));
 sky130_fd_sc_hd__o21bai_1 _26709_ (.A1(_03686_),
    .A2(_03688_),
    .B1_N(_03687_),
    .Y(_03788_));
 sky130_fd_sc_hd__a21o_1 _26710_ (.A1(_03786_),
    .A2(_03787_),
    .B1(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__nand3_1 _26711_ (.A(_03786_),
    .B(_03787_),
    .C(_03788_),
    .Y(_03790_));
 sky130_fd_sc_hd__a21o_1 _26712_ (.A1(_03668_),
    .A2(_03669_),
    .B1(_03673_),
    .X(_03791_));
 sky130_fd_sc_hd__a21oi_1 _26713_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03791_),
    .Y(_03793_));
 sky130_fd_sc_hd__and3_1 _26714_ (.A(_03789_),
    .B(_03790_),
    .C(_03791_),
    .X(_03794_));
 sky130_fd_sc_hd__a21boi_1 _26715_ (.A1(_03609_),
    .A2(_03691_),
    .B1_N(_03692_),
    .Y(_03795_));
 sky130_fd_sc_hd__o21ai_1 _26716_ (.A1(_03793_),
    .A2(_03794_),
    .B1(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__or3_1 _26717_ (.A(_03793_),
    .B(_03795_),
    .C(_03794_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_1 _26718_ (.A(_03796_),
    .B(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__o21ai_1 _26719_ (.A1(_03699_),
    .A2(_03706_),
    .B1(_03697_),
    .Y(_03799_));
 sky130_fd_sc_hd__xor2_1 _26720_ (.A(_03798_),
    .B(_03799_),
    .X(net122));
 sky130_fd_sc_hd__o2bb2a_1 _26721_ (.A1_N(_02711_),
    .A2_N(_03773_),
    .B1(_03774_),
    .B2(_03677_),
    .X(_03800_));
 sky130_fd_sc_hd__nand2_1 _26722_ (.A(_03729_),
    .B(_03731_),
    .Y(_03801_));
 sky130_fd_sc_hd__nor2_1 _26723_ (.A(net319),
    .B(_08660_),
    .Y(_03803_));
 sky130_fd_sc_hd__a21oi_1 _26724_ (.A1(net152),
    .A2(net158),
    .B1(_08658_),
    .Y(_03804_));
 sky130_fd_sc_hd__a221o_2 _26725_ (.A1(_08878_),
    .A2(_09299_),
    .B1(_08670_),
    .B2(_08657_),
    .C1(_03803_),
    .X(_03805_));
 sky130_fd_sc_hd__o221ai_4 _26726_ (.A1(_03286_),
    .A2(net152),
    .B1(_03803_),
    .B2(_03804_),
    .C1(_09299_),
    .Y(_03806_));
 sky130_fd_sc_hd__a21oi_1 _26727_ (.A1(net144),
    .A2(_03720_),
    .B1(_03721_),
    .Y(_03807_));
 sky130_fd_sc_hd__o21ai_1 _26728_ (.A1(_09299_),
    .A2(_03719_),
    .B1(_03722_),
    .Y(_03808_));
 sky130_fd_sc_hd__o2111ai_2 _26729_ (.A1(_09299_),
    .A2(_03719_),
    .B1(_03722_),
    .C1(_03805_),
    .D1(_03806_),
    .Y(_03809_));
 sky130_fd_sc_hd__a21o_1 _26730_ (.A1(_03805_),
    .A2(_03806_),
    .B1(_03807_),
    .X(_03810_));
 sky130_fd_sc_hd__nand3_1 _26731_ (.A(_03805_),
    .B(_03806_),
    .C(_03808_),
    .Y(_03811_));
 sky130_fd_sc_hd__a21o_1 _26732_ (.A1(_03805_),
    .A2(_03806_),
    .B1(_03808_),
    .X(_03812_));
 sky130_fd_sc_hd__o211ai_1 _26733_ (.A1(net140),
    .A2(_10542_),
    .B1(_03809_),
    .C1(_03810_),
    .Y(_03814_));
 sky130_fd_sc_hd__nand3_1 _26734_ (.A(_03812_),
    .B(_10545_),
    .C(_03811_),
    .Y(_03815_));
 sky130_fd_sc_hd__a22o_1 _26735_ (.A1(net139),
    .A2(_10544_),
    .B1(_03809_),
    .B2(_03810_),
    .X(_03816_));
 sky130_fd_sc_hd__a211o_1 _26736_ (.A1(_03811_),
    .A2(_03812_),
    .B1(net140),
    .C1(_10542_),
    .X(_03817_));
 sky130_fd_sc_hd__nand4_1 _26737_ (.A(_03729_),
    .B(_03731_),
    .C(_03814_),
    .D(_03815_),
    .Y(_03818_));
 sky130_fd_sc_hd__a22o_1 _26738_ (.A1(_03729_),
    .A2(_03731_),
    .B1(_03814_),
    .B2(_03815_),
    .X(_03819_));
 sky130_fd_sc_hd__a21oi_1 _26739_ (.A1(_03818_),
    .A2(_03819_),
    .B1(_12099_),
    .Y(_03820_));
 sky130_fd_sc_hd__o311a_1 _26740_ (.A1(_10566_),
    .A2(_11040_),
    .A3(_11742_),
    .B1(_03818_),
    .C1(_03819_),
    .X(_03821_));
 sky130_fd_sc_hd__o211ai_1 _26741_ (.A1(net141),
    .A2(_11742_),
    .B1(_03818_),
    .C1(_03819_),
    .Y(_03822_));
 sky130_fd_sc_hd__nand2_1 _26742_ (.A(_03735_),
    .B(_03739_),
    .Y(_03823_));
 sky130_fd_sc_hd__o211ai_2 _26743_ (.A1(_03820_),
    .A2(_03821_),
    .B1(_03735_),
    .C1(_03739_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand3b_1 _26744_ (.A_N(_03820_),
    .B(_03822_),
    .C(_03823_),
    .Y(_03826_));
 sky130_fd_sc_hd__a21oi_1 _26745_ (.A1(_03825_),
    .A2(_03826_),
    .B1(_00736_),
    .Y(_03827_));
 sky130_fd_sc_hd__and3_1 _26746_ (.A(_03825_),
    .B(_03826_),
    .C(_00736_),
    .X(_03828_));
 sky130_fd_sc_hd__a21boi_1 _26747_ (.A1(_03743_),
    .A2(_00736_),
    .B1_N(_03744_),
    .Y(_03829_));
 sky130_fd_sc_hd__nor3_1 _26748_ (.A(_03827_),
    .B(_03829_),
    .C(_03828_),
    .Y(_03830_));
 sky130_fd_sc_hd__o21a_1 _26749_ (.A1(_03827_),
    .A2(_03828_),
    .B1(_03829_),
    .X(_03831_));
 sky130_fd_sc_hd__nor3_2 _26750_ (.A(_02949_),
    .B(_03830_),
    .C(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__o22a_1 _26751_ (.A1(_02711_),
    .A2(_02945_),
    .B1(_03830_),
    .B2(_03831_),
    .X(_03833_));
 sky130_fd_sc_hd__o221a_1 _26752_ (.A1(_02949_),
    .A2(_03752_),
    .B1(_03832_),
    .B2(_03833_),
    .C1(_03751_),
    .X(_03834_));
 sky130_fd_sc_hd__o221ai_2 _26753_ (.A1(_02949_),
    .A2(_03752_),
    .B1(_03832_),
    .B2(_03833_),
    .C1(_03751_),
    .Y(_03837_));
 sky130_fd_sc_hd__a211oi_1 _26754_ (.A1(_03751_),
    .A2(_03754_),
    .B1(_03832_),
    .C1(_03833_),
    .Y(_03838_));
 sky130_fd_sc_hd__a211o_1 _26755_ (.A1(_03751_),
    .A2(_03754_),
    .B1(_03832_),
    .C1(_03833_),
    .X(_03839_));
 sky130_fd_sc_hd__a22oi_2 _26756_ (.A1(net25),
    .A2(_08006_),
    .B1(net160),
    .B2(net238),
    .Y(_03840_));
 sky130_fd_sc_hd__xnor2_1 _26757_ (.A(_03765_),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__nor2_1 _26758_ (.A(_03265_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__and3b_1 _26759_ (.A_N(_03260_),
    .B(_03841_),
    .C(_02700_),
    .X(_03843_));
 sky130_fd_sc_hd__o32a_1 _26760_ (.A1(_11741_),
    .A2(_00360_),
    .A3(_02708_),
    .B1(_03842_),
    .B2(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__nor4_1 _26761_ (.A(_00364_),
    .B(_02708_),
    .C(_03842_),
    .D(_03843_),
    .Y(_03845_));
 sky130_fd_sc_hd__or2_1 _26762_ (.A(_03844_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__xor2_1 _26763_ (.A(_03772_),
    .B(_03846_),
    .X(_03848_));
 sky130_fd_sc_hd__o21bai_1 _26764_ (.A1(_03834_),
    .A2(_03838_),
    .B1_N(_03848_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand3_1 _26765_ (.A(_03837_),
    .B(_03839_),
    .C(_03848_),
    .Y(_03850_));
 sky130_fd_sc_hd__nand2_1 _26766_ (.A(_03849_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__o211a_1 _26767_ (.A1(_03777_),
    .A2(_03760_),
    .B1(_03762_),
    .C1(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__o211ai_1 _26768_ (.A1(_03777_),
    .A2(_03760_),
    .B1(_03762_),
    .C1(_03851_),
    .Y(_03853_));
 sky130_fd_sc_hd__a21o_1 _26769_ (.A1(_03762_),
    .A2(_03780_),
    .B1(_03851_),
    .X(_03854_));
 sky130_fd_sc_hd__a21boi_1 _26770_ (.A1(_03853_),
    .A2(_03854_),
    .B1_N(_03800_),
    .Y(_03855_));
 sky130_fd_sc_hd__nor3b_1 _26771_ (.A(_03800_),
    .B(_03852_),
    .C_N(_03854_),
    .Y(_03856_));
 sky130_fd_sc_hd__o211ai_1 _26772_ (.A1(_03855_),
    .A2(_03856_),
    .B1(_03783_),
    .C1(_03787_),
    .Y(_03857_));
 sky130_fd_sc_hd__a211o_1 _26773_ (.A1(_03783_),
    .A2(_03787_),
    .B1(_03855_),
    .C1(_03856_),
    .X(_03859_));
 sky130_fd_sc_hd__nand2_1 _26774_ (.A(_03857_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__o21bai_2 _26775_ (.A1(_03763_),
    .A2(_03765_),
    .B1_N(_03768_),
    .Y(_03861_));
 sky130_fd_sc_hd__xnor2_1 _26776_ (.A(_03860_),
    .B(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__a21bo_1 _26777_ (.A1(_03789_),
    .A2(_03791_),
    .B1_N(_03790_),
    .X(_03863_));
 sky130_fd_sc_hd__and2_1 _26778_ (.A(_03862_),
    .B(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__xnor2_1 _26779_ (.A(_03862_),
    .B(_03863_),
    .Y(_03865_));
 sky130_fd_sc_hd__nand3b_1 _26780_ (.A_N(_03708_),
    .B(_03796_),
    .C(_03797_),
    .Y(_03866_));
 sky130_fd_sc_hd__o21bai_1 _26781_ (.A1(_03705_),
    .A2(_03702_),
    .B1_N(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__a21bo_1 _26782_ (.A1(_03697_),
    .A2(_03797_),
    .B1_N(_03796_),
    .X(_03868_));
 sky130_fd_sc_hd__o21ai_1 _26783_ (.A1(_03866_),
    .A2(_03706_),
    .B1(_03868_),
    .Y(_03870_));
 sky130_fd_sc_hd__a21oi_1 _26784_ (.A1(_03867_),
    .A2(_03868_),
    .B1(_03865_),
    .Y(_03871_));
 sky130_fd_sc_hd__a21o_1 _26785_ (.A1(_03867_),
    .A2(_03868_),
    .B1(_03865_),
    .X(_03872_));
 sky130_fd_sc_hd__xnor2_1 _26786_ (.A(_03865_),
    .B(_03870_),
    .Y(net123));
 sky130_fd_sc_hd__a21bo_1 _26787_ (.A1(_03857_),
    .A2(_03861_),
    .B1_N(_03859_),
    .X(_03873_));
 sky130_fd_sc_hd__o21ai_1 _26788_ (.A1(_03800_),
    .A2(_03852_),
    .B1(_03854_),
    .Y(_03874_));
 sky130_fd_sc_hd__o32a_1 _26789_ (.A1(_02712_),
    .A2(_03842_),
    .A3(_03843_),
    .B1(_03846_),
    .B2(_03772_),
    .X(_03875_));
 sky130_fd_sc_hd__a31o_1 _26790_ (.A1(_03801_),
    .A2(_03816_),
    .A3(_03817_),
    .B1(_03821_),
    .X(_03876_));
 sky130_fd_sc_hd__o22a_1 _26791_ (.A1(net319),
    .A2(_08660_),
    .B1(net152),
    .B2(_08658_),
    .X(_03877_));
 sky130_fd_sc_hd__a31o_1 _26792_ (.A1(_03805_),
    .A2(_03807_),
    .A3(_03806_),
    .B1(_10546_),
    .X(_03878_));
 sky130_fd_sc_hd__o21ai_1 _26793_ (.A1(net140),
    .A2(_10542_),
    .B1(_03810_),
    .Y(_03880_));
 sky130_fd_sc_hd__and4_1 _26794_ (.A(_03805_),
    .B(_03880_),
    .C(_03877_),
    .D(_03878_),
    .X(_03881_));
 sky130_fd_sc_hd__a22oi_1 _26795_ (.A1(_03877_),
    .A2(_03805_),
    .B1(_03880_),
    .B2(_03878_),
    .Y(_03882_));
 sky130_fd_sc_hd__a22o_1 _26796_ (.A1(net143),
    .A2(_11743_),
    .B1(_00364_),
    .B2(_00367_),
    .X(_03883_));
 sky130_fd_sc_hd__or4_1 _26797_ (.A(net141),
    .B(_11742_),
    .C(net131),
    .D(_00366_),
    .X(_03884_));
 sky130_fd_sc_hd__a211oi_1 _26798_ (.A1(_03883_),
    .A2(_03884_),
    .B1(_03881_),
    .C1(_03882_),
    .Y(_03885_));
 sky130_fd_sc_hd__o211a_1 _26799_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03883_),
    .C1(_03884_),
    .X(_03886_));
 sky130_fd_sc_hd__nor2_1 _26800_ (.A(_03885_),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__a21boi_1 _26801_ (.A1(_03825_),
    .A2(_00736_),
    .B1_N(_03826_),
    .Y(_03888_));
 sky130_fd_sc_hd__xnor2_1 _26802_ (.A(_03876_),
    .B(_03887_),
    .Y(_03889_));
 sky130_fd_sc_hd__xor2_1 _26803_ (.A(_02947_),
    .B(_03889_),
    .X(_03891_));
 sky130_fd_sc_hd__xor2_1 _26804_ (.A(_03843_),
    .B(_03888_),
    .X(_03892_));
 sky130_fd_sc_hd__xnor2_1 _26805_ (.A(_03891_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__nor3b_1 _26806_ (.A(_03765_),
    .B(_03840_),
    .C_N(_03875_),
    .Y(_03894_));
 sky130_fd_sc_hd__o21ba_1 _26807_ (.A1(_03765_),
    .A2(_03840_),
    .B1_N(_03875_),
    .X(_03895_));
 sky130_fd_sc_hd__nor2_1 _26808_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__or3_1 _26809_ (.A(_03830_),
    .B(_03832_),
    .C(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__o21ai_1 _26810_ (.A1(_03830_),
    .A2(_03832_),
    .B1(_03896_),
    .Y(_03898_));
 sky130_fd_sc_hd__and2_1 _26811_ (.A(_03897_),
    .B(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__xnor2_1 _26812_ (.A(_03893_),
    .B(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__a21oi_1 _26813_ (.A1(_03837_),
    .A2(_03848_),
    .B1(_03838_),
    .Y(_03902_));
 sky130_fd_sc_hd__xnor2_1 _26814_ (.A(_03900_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__xor2_1 _26815_ (.A(_03874_),
    .B(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__xnor2_1 _26816_ (.A(_03873_),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__nand3b_1 _26817_ (.A_N(_03864_),
    .B(_03872_),
    .C(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__o21bai_1 _26818_ (.A1(_03864_),
    .A2(_03871_),
    .B1_N(_03905_),
    .Y(_03907_));
 sky130_fd_sc_hd__nand2_1 _26819_ (.A(_03906_),
    .B(_03907_),
    .Y(net124));
 sky130_fd_sc_hd__a2bb2o_1 _26820_ (.A1_N(_07133_),
    .A2_N(_08174_),
    .B1(_10719_),
    .B2(_10796_),
    .X(_03908_));
 sky130_fd_sc_hd__a22o_1 _26821_ (.A1(_07045_),
    .A2(_08141_),
    .B1(_10828_),
    .B2(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__o31a_1 _26822_ (.A1(_07056_),
    .A2(_08130_),
    .A3(_09402_),
    .B1(_03909_),
    .X(net128));
 sky130_fd_sc_hd__o221a_1 _26823_ (.A1(net12),
    .A2(_03286_),
    .B1(_04484_),
    .B2(_04320_),
    .C1(net1),
    .X(_03911_));
 sky130_fd_sc_hd__o221a_1 _26824_ (.A1(_03176_),
    .A2(net44),
    .B1(_04298_),
    .B2(_04506_),
    .C1(net33),
    .X(_03912_));
 sky130_fd_sc_hd__or2_1 _26825_ (.A(_03911_),
    .B(_03912_),
    .X(net76));
 sky130_fd_sc_hd__a21oi_1 _26826_ (.A1(_04298_),
    .A2(_04320_),
    .B1(_04594_),
    .Y(_03913_));
 sky130_fd_sc_hd__nor2_1 _26827_ (.A(_04605_),
    .B(_03913_),
    .Y(net87));
 sky130_fd_sc_hd__clkbuf_16 input1 (.A(multiplicand[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_12 input2 (.A(multiplicand[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(multiplicand[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_12 input4 (.A(multiplicand[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(multiplicand[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input6 (.A(multiplicand[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input7 (.A(multiplicand[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_12 input8 (.A(multiplicand[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input9 (.A(multiplicand[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(multiplicand[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_12 input11 (.A(multiplicand[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(multiplicand[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input13 (.A(multiplicand[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_12 input14 (.A(multiplicand[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input15 (.A(multiplicand[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_12 input16 (.A(multiplicand[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input17 (.A(multiplicand[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_12 input18 (.A(multiplicand[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_12 input19 (.A(multiplicand[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_12 input20 (.A(multiplicand[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_12 input21 (.A(multiplicand[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_12 input22 (.A(multiplicand[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_12 input23 (.A(multiplicand[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_12 input24 (.A(multiplicand[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_12 input25 (.A(multiplicand[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_12 input26 (.A(multiplicand[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_12 input27 (.A(multiplicand[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_12 input28 (.A(multiplicand[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_12 input29 (.A(multiplicand[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_12 input30 (.A(multiplicand[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_12 input31 (.A(multiplicand[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_12 input32 (.A(multiplicand[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_16 input33 (.A(multiplier[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_12 input34 (.A(multiplier[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_12 input35 (.A(multiplier[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_12 input36 (.A(multiplier[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_12 input37 (.A(multiplier[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_8 input38 (.A(multiplier[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_12 input39 (.A(multiplier[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_12 input40 (.A(multiplier[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_12 input41 (.A(multiplier[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_12 input42 (.A(multiplier[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_12 input43 (.A(multiplier[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_12 input44 (.A(multiplier[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_12 input45 (.A(multiplier[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_12 input46 (.A(multiplier[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_12 input47 (.A(multiplier[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_12 input48 (.A(multiplier[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_12 input49 (.A(multiplier[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_8 input50 (.A(multiplier[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_12 input51 (.A(multiplier[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_12 input52 (.A(multiplier[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_8 input53 (.A(multiplier[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_12 input54 (.A(multiplier[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_16 input55 (.A(multiplier[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 input56 (.A(multiplier[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_16 input57 (.A(multiplier[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_12 input58 (.A(multiplier[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_12 input59 (.A(multiplier[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input60 (.A(multiplier[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_12 input61 (.A(multiplier[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_16 input62 (.A(multiplier[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_12 input63 (.A(multiplier[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_12 input64 (.A(multiplier[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(product[0]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(product[10]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(product[11]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(product[12]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(product[13]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(product[14]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(product[15]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(product[16]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(product[17]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(product[18]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(product[19]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(product[1]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(product[20]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(product[21]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(product[22]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(product[23]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(product[24]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(product[25]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(product[26]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(product[27]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(product[28]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(product[29]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(product[2]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(product[30]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(product[31]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(product[32]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(product[33]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(product[34]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(product[35]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(product[36]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(product[37]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(product[38]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(product[39]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(product[3]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(product[40]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(product[41]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(product[42]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(product[43]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(product[44]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(product[45]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(product[46]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(product[47]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(product[48]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(product[49]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(product[4]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(product[50]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(product[51]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(product[52]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(product[53]));
 sky130_fd_sc_hd__buf_1 output114 (.A(net114),
    .X(product[54]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(product[55]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(product[56]));
 sky130_fd_sc_hd__buf_1 output117 (.A(net117),
    .X(product[57]));
 sky130_fd_sc_hd__buf_1 output118 (.A(net118),
    .X(product[58]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(product[59]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(product[5]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(product[60]));
 sky130_fd_sc_hd__buf_1 output122 (.A(net122),
    .X(product[61]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(product[62]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(product[63]));
 sky130_fd_sc_hd__buf_1 output125 (.A(net125),
    .X(product[6]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(product[7]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(product[8]));
 sky130_fd_sc_hd__buf_1 output128 (.A(net128),
    .X(product[9]));
 sky130_fd_sc_hd__clkbuf_8 max_cap129 (.A(_00737_),
    .X(net129));
 sky130_fd_sc_hd__buf_8 max_cap130 (.A(_00363_),
    .X(net130));
 sky130_fd_sc_hd__buf_8 max_cap131 (.A(_00363_),
    .X(net131));
 sky130_fd_sc_hd__buf_8 max_cap132 (.A(_12098_),
    .X(net132));
 sky130_fd_sc_hd__buf_12 max_cap133 (.A(_10545_),
    .X(net133));
 sky130_fd_sc_hd__buf_12 max_cap134 (.A(_10544_),
    .X(net134));
 sky130_fd_sc_hd__buf_8 max_cap135 (.A(net137),
    .X(net135));
 sky130_fd_sc_hd__buf_8 max_cap136 (.A(_10542_),
    .X(net136));
 sky130_fd_sc_hd__buf_12 max_cap137 (.A(_10542_),
    .X(net137));
 sky130_fd_sc_hd__buf_8 wire138 (.A(_10541_),
    .X(net138));
 sky130_fd_sc_hd__buf_12 max_cap139 (.A(_10541_),
    .X(net139));
 sky130_fd_sc_hd__buf_12 max_cap140 (.A(_10540_),
    .X(net140));
 sky130_fd_sc_hd__buf_12 max_cap141 (.A(_11042_),
    .X(net141));
 sky130_fd_sc_hd__buf_8 max_cap142 (.A(_11041_),
    .X(net142));
 sky130_fd_sc_hd__buf_6 max_cap143 (.A(_11041_),
    .X(net143));
 sky130_fd_sc_hd__buf_12 max_cap144 (.A(_09300_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_16 max_cap145 (.A(_09299_),
    .X(net145));
 sky130_fd_sc_hd__buf_12 max_cap146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_12 max_cap147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_16 max_cap148 (.A(_09299_),
    .X(net148));
 sky130_fd_sc_hd__buf_12 max_cap149 (.A(_08878_),
    .X(net149));
 sky130_fd_sc_hd__buf_8 max_cap150 (.A(_08665_),
    .X(net150));
 sky130_fd_sc_hd__buf_12 max_cap151 (.A(_08665_),
    .X(net151));
 sky130_fd_sc_hd__buf_6 max_cap152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_12 max_cap153 (.A(_08665_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_8 max_cap154 (.A(_08207_),
    .X(net154));
 sky130_fd_sc_hd__buf_12 max_cap155 (.A(_05935_),
    .X(net155));
 sky130_fd_sc_hd__buf_4 wire156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 max_cap157 (.A(_08877_),
    .X(net157));
 sky130_fd_sc_hd__buf_12 max_cap158 (.A(_08668_),
    .X(net158));
 sky130_fd_sc_hd__buf_8 wire159 (.A(_08664_),
    .X(net159));
 sky130_fd_sc_hd__buf_6 max_cap160 (.A(_08664_),
    .X(net160));
 sky130_fd_sc_hd__buf_12 max_cap161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_16 max_cap162 (.A(_08208_),
    .X(net162));
 sky130_fd_sc_hd__buf_12 max_cap163 (.A(_08208_),
    .X(net163));
 sky130_fd_sc_hd__buf_12 max_cap164 (.A(_08204_),
    .X(net164));
 sky130_fd_sc_hd__buf_12 max_cap165 (.A(_07769_),
    .X(net165));
 sky130_fd_sc_hd__buf_8 max_cap166 (.A(_07769_),
    .X(net166));
 sky130_fd_sc_hd__buf_8 max_cap167 (.A(_07503_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_16 wire168 (.A(_07076_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_16 max_cap169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_12 max_cap170 (.A(_07076_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_16 max_cap171 (.A(_06762_),
    .X(net171));
 sky130_fd_sc_hd__buf_12 max_cap172 (.A(_06452_),
    .X(net172));
 sky130_fd_sc_hd__buf_12 max_cap173 (.A(_06221_),
    .X(net173));
 sky130_fd_sc_hd__buf_12 max_cap174 (.A(net176),
    .X(net174));
 sky130_fd_sc_hd__buf_12 max_cap175 (.A(_05931_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_16 max_cap176 (.A(_05931_),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_16 wire177 (.A(_05553_),
    .X(net177));
 sky130_fd_sc_hd__buf_12 max_cap178 (.A(_05549_),
    .X(net178));
 sky130_fd_sc_hd__buf_12 max_cap179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_12 max_cap180 (.A(_05292_),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_16 max_cap181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_12 max_cap182 (.A(_05290_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_16 max_cap183 (.A(_05074_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_16 max_cap184 (.A(_04789_),
    .X(net184));
 sky130_fd_sc_hd__buf_12 max_cap185 (.A(_04789_),
    .X(net185));
 sky130_fd_sc_hd__buf_12 max_cap186 (.A(_04559_),
    .X(net186));
 sky130_fd_sc_hd__buf_6 max_cap187 (.A(_04412_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_16 max_cap188 (.A(_04409_),
    .X(net188));
 sky130_fd_sc_hd__buf_4 wire189 (.A(_06761_),
    .X(net189));
 sky130_fd_sc_hd__buf_4 max_cap190 (.A(_06761_),
    .X(net190));
 sky130_fd_sc_hd__buf_4 max_cap191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_4 wire192 (.A(_06757_),
    .X(net192));
 sky130_fd_sc_hd__buf_4 max_cap193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_4 max_cap194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 max_cap195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__buf_4 max_cap196 (.A(_06757_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_8 max_cap197 (.A(_06449_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 wire198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 max_cap199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_6 max_cap200 (.A(_06449_),
    .X(net200));
 sky130_fd_sc_hd__buf_8 max_cap201 (.A(_06219_),
    .X(net201));
 sky130_fd_sc_hd__buf_8 max_cap202 (.A(_06219_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_8 max_cap203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__buf_6 max_cap204 (.A(_05930_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 max_cap205 (.A(_05930_),
    .X(net205));
 sky130_fd_sc_hd__buf_4 max_cap206 (.A(_05552_),
    .X(net206));
 sky130_fd_sc_hd__buf_4 max_cap207 (.A(_05552_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_16 wire208 (.A(_05073_),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 wire209 (.A(_05072_),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 wire210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 wire211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 max_cap212 (.A(_05072_),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_8 max_cap213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 max_cap214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_8 wire215 (.A(_04790_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_8 max_cap216 (.A(_04558_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 max_cap217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 wire218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_8 max_cap219 (.A(_04555_),
    .X(net219));
 sky130_fd_sc_hd__buf_6 max_cap220 (.A(_04555_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 wire221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 max_cap222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 wire223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_4 wire224 (.A(net226),
    .X(net224));
 sky130_fd_sc_hd__buf_4 wire225 (.A(_04411_),
    .X(net225));
 sky130_fd_sc_hd__buf_4 max_cap226 (.A(_04411_),
    .X(net226));
 sky130_fd_sc_hd__buf_8 max_cap227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_8 max_cap228 (.A(_04132_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_16 max_cap229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_16 max_cap230 (.A(_04130_),
    .X(net230));
 sky130_fd_sc_hd__buf_12 max_cap231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_12 max_cap232 (.A(_03958_),
    .X(net232));
 sky130_fd_sc_hd__buf_12 max_cap233 (.A(_03958_),
    .X(net233));
 sky130_fd_sc_hd__buf_8 max_cap234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_8 max_cap235 (.A(_12977_),
    .X(net235));
 sky130_fd_sc_hd__buf_8 max_cap236 (.A(_11453_),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_16 max_cap237 (.A(_08881_),
    .X(net237));
 sky130_fd_sc_hd__buf_12 max_cap238 (.A(_08005_),
    .X(net238));
 sky130_fd_sc_hd__buf_12 max_cap239 (.A(_07305_),
    .X(net239));
 sky130_fd_sc_hd__buf_12 max_cap240 (.A(_06863_),
    .X(net240));
 sky130_fd_sc_hd__buf_12 max_cap241 (.A(_05928_),
    .X(net241));
 sky130_fd_sc_hd__buf_12 max_cap242 (.A(_04985_),
    .X(net242));
 sky130_fd_sc_hd__buf_12 max_cap243 (.A(_04895_),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_16 max_cap244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_16 max_cap245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_6 max_cap246 (.A(_03956_),
    .X(net246));
 sky130_fd_sc_hd__buf_6 max_cap247 (.A(_03951_),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_16 max_cap248 (.A(_02453_),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_16 max_cap249 (.A(_02453_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_16 max_cap250 (.A(_00657_),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_16 wire251 (.A(_12999_),
    .X(net251));
 sky130_fd_sc_hd__buf_12 max_cap252 (.A(_11771_),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_16 max_cap253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_16 max_cap254 (.A(_11431_),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_16 max_cap255 (.A(_09676_),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_16 wire256 (.A(_08678_),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_16 max_cap257 (.A(_07253_),
    .X(net257));
 sky130_fd_sc_hd__buf_12 max_cap258 (.A(_07253_),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_16 max_cap259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_16 max_cap260 (.A(net263),
    .X(net260));
 sky130_fd_sc_hd__buf_12 max_cap261 (.A(net263),
    .X(net261));
 sky130_fd_sc_hd__buf_12 max_cap262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__buf_12 max_cap263 (.A(_06530_),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_16 max_cap264 (.A(_06508_),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_16 max_cap265 (.A(_05863_),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_16 max_cap266 (.A(_04998_),
    .X(net266));
 sky130_fd_sc_hd__buf_12 max_cap267 (.A(_04747_),
    .X(net267));
 sky130_fd_sc_hd__buf_12 max_cap268 (.A(_08206_),
    .X(net268));
 sky130_fd_sc_hd__buf_12 max_cap269 (.A(_07223_),
    .X(net269));
 sky130_fd_sc_hd__buf_4 max_cap270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_4 max_cap271 (.A(_07073_),
    .X(net271));
 sky130_fd_sc_hd__buf_4 max_cap272 (.A(_07073_),
    .X(net272));
 sky130_fd_sc_hd__buf_12 max_cap273 (.A(_06324_),
    .X(net273));
 sky130_fd_sc_hd__buf_12 wire274 (.A(_06026_),
    .X(net274));
 sky130_fd_sc_hd__buf_12 max_cap275 (.A(_05762_),
    .X(net275));
 sky130_fd_sc_hd__buf_12 max_cap276 (.A(_05225_),
    .X(net276));
 sky130_fd_sc_hd__buf_4 max_cap277 (.A(_04786_),
    .X(net277));
 sky130_fd_sc_hd__buf_4 max_cap278 (.A(_04786_),
    .X(net278));
 sky130_fd_sc_hd__buf_12 max_cap279 (.A(_04480_),
    .X(net279));
 sky130_fd_sc_hd__buf_12 max_cap280 (.A(_04267_),
    .X(net280));
 sky130_fd_sc_hd__buf_12 max_cap281 (.A(_04215_),
    .X(net281));
 sky130_fd_sc_hd__buf_4 max_cap282 (.A(_03953_),
    .X(net282));
 sky130_fd_sc_hd__buf_4 max_cap283 (.A(_03953_),
    .X(net283));
 sky130_fd_sc_hd__buf_4 max_cap284 (.A(_03953_),
    .X(net284));
 sky130_fd_sc_hd__buf_12 max_cap285 (.A(_03704_),
    .X(net285));
 sky130_fd_sc_hd__buf_4 max_cap286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_4 max_cap287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_4 max_cap288 (.A(_11376_),
    .X(net288));
 sky130_fd_sc_hd__buf_12 wire289 (.A(_10313_),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_8 max_cap290 (.A(_09654_),
    .X(net290));
 sky130_fd_sc_hd__buf_12 max_cap291 (.A(_08250_),
    .X(net291));
 sky130_fd_sc_hd__buf_12 wire292 (.A(_06826_),
    .X(net292));
 sky130_fd_sc_hd__buf_4 max_cap293 (.A(net296),
    .X(net293));
 sky130_fd_sc_hd__buf_4 wire294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_4 max_cap295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_4 max_cap296 (.A(_06497_),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_8 max_cap297 (.A(_05852_),
    .X(net297));
 sky130_fd_sc_hd__buf_12 max_cap298 (.A(_05720_),
    .X(net298));
 sky130_fd_sc_hd__buf_12 max_cap299 (.A(_05688_),
    .X(net299));
 sky130_fd_sc_hd__buf_4 max_cap300 (.A(_05009_),
    .X(net300));
 sky130_fd_sc_hd__buf_4 max_cap301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__buf_4 max_cap302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_4 max_cap303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_4 max_cap304 (.A(_05009_),
    .X(net304));
 sky130_fd_sc_hd__buf_12 max_cap305 (.A(_04889_),
    .X(net305));
 sky130_fd_sc_hd__buf_4 max_cap306 (.A(_04736_),
    .X(net306));
 sky130_fd_sc_hd__buf_4 max_cap307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__buf_4 max_cap308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_4 max_cap309 (.A(net312),
    .X(net309));
 sky130_fd_sc_hd__buf_4 max_cap310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__buf_4 max_cap311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_4 wire312 (.A(_04736_),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_8 wire313 (.A(net315),
    .X(net313));
 sky130_fd_sc_hd__buf_6 max_cap314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_8 max_cap315 (.A(_04714_),
    .X(net315));
 sky130_fd_sc_hd__buf_12 max_cap316 (.A(_04660_),
    .X(net316));
 sky130_fd_sc_hd__buf_12 max_cap317 (.A(_04627_),
    .X(net317));
 sky130_fd_sc_hd__buf_12 max_cap318 (.A(_04419_),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_16 load_slew319 (.A(_04277_),
    .X(net319));
endmodule
