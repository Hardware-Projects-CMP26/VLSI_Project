module ALU (select,
    A,
    B,
    result);
 input select;
 input [31:0] A;
 input [31:0] B;
 output [31:0] result;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire \adder_inst.fraction1[0] ;
 wire \adder_inst.fraction1_32neg[0] ;
 wire \adder_inst.fraction1_32neg[10] ;
 wire \adder_inst.fraction1_32neg[11] ;
 wire \adder_inst.fraction1_32neg[12] ;
 wire \adder_inst.fraction1_32neg[13] ;
 wire \adder_inst.fraction1_32neg[14] ;
 wire \adder_inst.fraction1_32neg[15] ;
 wire \adder_inst.fraction1_32neg[16] ;
 wire \adder_inst.fraction1_32neg[17] ;
 wire \adder_inst.fraction1_32neg[18] ;
 wire \adder_inst.fraction1_32neg[19] ;
 wire \adder_inst.fraction1_32neg[1] ;
 wire \adder_inst.fraction1_32neg[20] ;
 wire \adder_inst.fraction1_32neg[21] ;
 wire \adder_inst.fraction1_32neg[22] ;
 wire \adder_inst.fraction1_32neg[2] ;
 wire \adder_inst.fraction1_32neg[3] ;
 wire \adder_inst.fraction1_32neg[4] ;
 wire \adder_inst.fraction1_32neg[5] ;
 wire \adder_inst.fraction1_32neg[6] ;
 wire \adder_inst.fraction1_32neg[7] ;
 wire \adder_inst.fraction1_32neg[8] ;
 wire \adder_inst.fraction1_32neg[9] ;
 wire \adder_inst.fraction2[0] ;
 wire \adder_inst.fraction2_32neg[0] ;
 wire \adder_inst.fraction2_32neg[10] ;
 wire \adder_inst.fraction2_32neg[11] ;
 wire \adder_inst.fraction2_32neg[12] ;
 wire \adder_inst.fraction2_32neg[13] ;
 wire \adder_inst.fraction2_32neg[14] ;
 wire \adder_inst.fraction2_32neg[15] ;
 wire \adder_inst.fraction2_32neg[16] ;
 wire \adder_inst.fraction2_32neg[17] ;
 wire \adder_inst.fraction2_32neg[18] ;
 wire \adder_inst.fraction2_32neg[19] ;
 wire \adder_inst.fraction2_32neg[1] ;
 wire \adder_inst.fraction2_32neg[20] ;
 wire \adder_inst.fraction2_32neg[21] ;
 wire \adder_inst.fraction2_32neg[22] ;
 wire \adder_inst.fraction2_32neg[2] ;
 wire \adder_inst.fraction2_32neg[3] ;
 wire \adder_inst.fraction2_32neg[4] ;
 wire \adder_inst.fraction2_32neg[5] ;
 wire \adder_inst.fraction2_32neg[6] ;
 wire \adder_inst.fraction2_32neg[7] ;
 wire \adder_inst.fraction2_32neg[8] ;
 wire \adder_inst.fraction2_32neg[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;

 sky130_fd_sc_hd__inv_2 _05411_ (.A(net22),
    .Y(_00966_));
 sky130_fd_sc_hd__inv_2 _05412_ (.A(net20),
    .Y(_00977_));
 sky130_fd_sc_hd__inv_2 _05413_ (.A(net19),
    .Y(_00988_));
 sky130_fd_sc_hd__inv_2 _05414_ (.A(net49),
    .Y(_00999_));
 sky130_fd_sc_hd__inv_2 _05415_ (.A(net48),
    .Y(_01010_));
 sky130_fd_sc_hd__inv_2 _05416_ (.A(net16),
    .Y(_01021_));
 sky130_fd_sc_hd__inv_2 _05417_ (.A(net15),
    .Y(_01032_));
 sky130_fd_sc_hd__inv_6 _05418_ (.A(net47),
    .Y(_01043_));
 sky130_fd_sc_hd__inv_6 _05419_ (.A(net45),
    .Y(_01054_));
 sky130_fd_sc_hd__clkinv_4 _05420_ (.A(net43),
    .Y(_01065_));
 sky130_fd_sc_hd__inv_4 _05421_ (.A(net9),
    .Y(_01076_));
 sky130_fd_sc_hd__clkinv_4 _05422_ (.A(net38),
    .Y(_01087_));
 sky130_fd_sc_hd__inv_4 _05423_ (.A(net5),
    .Y(_01098_));
 sky130_fd_sc_hd__clkinv_4 _05424_ (.A(net35),
    .Y(_01109_));
 sky130_fd_sc_hd__inv_2 _05425_ (.A(net3),
    .Y(_01120_));
 sky130_fd_sc_hd__inv_4 _05426_ (.A(net2),
    .Y(_01131_));
 sky130_fd_sc_hd__inv_2 _05427_ (.A(net63),
    .Y(_01142_));
 sky130_fd_sc_hd__clkinv_4 _05428_ (.A(net31),
    .Y(_01153_));
 sky130_fd_sc_hd__inv_2 _05429_ (.A(net62),
    .Y(_01164_));
 sky130_fd_sc_hd__inv_4 _05430_ (.A(net30),
    .Y(_01175_));
 sky130_fd_sc_hd__inv_4 _05431_ (.A(net29),
    .Y(_01186_));
 sky130_fd_sc_hd__clkinv_4 _05432_ (.A(net60),
    .Y(_01197_));
 sky130_fd_sc_hd__clkinv_4 _05433_ (.A(net27),
    .Y(_01208_));
 sky130_fd_sc_hd__inv_2 _05434_ (.A(net26),
    .Y(_01219_));
 sky130_fd_sc_hd__clkinv_4 _05435_ (.A(net55),
    .Y(_01230_));
 sky130_fd_sc_hd__inv_2 _05436_ (.A(net12),
    .Y(_01241_));
 sky130_fd_sc_hd__inv_2 _05437_ (.A(net44),
    .Y(_01252_));
 sky130_fd_sc_hd__clkinv_4 _05438_ (.A(net1),
    .Y(_01263_));
 sky130_fd_sc_hd__inv_2 _05439_ (.A(\adder_inst.fraction2_32neg[0] ),
    .Y(_01274_));
 sky130_fd_sc_hd__inv_2 _05440_ (.A(\adder_inst.fraction1_32neg[1] ),
    .Y(_01285_));
 sky130_fd_sc_hd__inv_2 _05441_ (.A(\adder_inst.fraction1_32neg[3] ),
    .Y(_01296_));
 sky130_fd_sc_hd__inv_2 _05442_ (.A(\adder_inst.fraction1_32neg[5] ),
    .Y(_01307_));
 sky130_fd_sc_hd__inv_2 _05443_ (.A(\adder_inst.fraction1_32neg[7] ),
    .Y(_01318_));
 sky130_fd_sc_hd__inv_2 _05444_ (.A(\adder_inst.fraction1_32neg[8] ),
    .Y(_01329_));
 sky130_fd_sc_hd__inv_2 _05445_ (.A(\adder_inst.fraction1_32neg[10] ),
    .Y(_01340_));
 sky130_fd_sc_hd__inv_2 _05446_ (.A(\adder_inst.fraction1_32neg[11] ),
    .Y(_01351_));
 sky130_fd_sc_hd__inv_2 _05447_ (.A(\adder_inst.fraction1_32neg[14] ),
    .Y(_01362_));
 sky130_fd_sc_hd__inv_2 _05448_ (.A(\adder_inst.fraction1_32neg[15] ),
    .Y(_01373_));
 sky130_fd_sc_hd__inv_2 _05449_ (.A(\adder_inst.fraction1_32neg[20] ),
    .Y(_01384_));
 sky130_fd_sc_hd__inv_2 _05450_ (.A(\adder_inst.fraction1_32neg[21] ),
    .Y(_01395_));
 sky130_fd_sc_hd__inv_2 _05451_ (.A(\adder_inst.fraction2_32neg[1] ),
    .Y(_01406_));
 sky130_fd_sc_hd__inv_2 _05452_ (.A(\adder_inst.fraction2_32neg[4] ),
    .Y(_01417_));
 sky130_fd_sc_hd__inv_2 _05453_ (.A(\adder_inst.fraction2_32neg[5] ),
    .Y(_01428_));
 sky130_fd_sc_hd__inv_2 _05454_ (.A(\adder_inst.fraction2_32neg[6] ),
    .Y(_01439_));
 sky130_fd_sc_hd__inv_2 _05455_ (.A(\adder_inst.fraction2_32neg[7] ),
    .Y(_01450_));
 sky130_fd_sc_hd__inv_2 _05456_ (.A(\adder_inst.fraction2_32neg[15] ),
    .Y(_01461_));
 sky130_fd_sc_hd__inv_2 _05457_ (.A(\adder_inst.fraction2_32neg[16] ),
    .Y(_01472_));
 sky130_fd_sc_hd__inv_2 _05458_ (.A(\adder_inst.fraction2_32neg[18] ),
    .Y(_01483_));
 sky130_fd_sc_hd__inv_2 _05459_ (.A(\adder_inst.fraction2_32neg[20] ),
    .Y(_01494_));
 sky130_fd_sc_hd__nor2_4 _05460_ (.A(net54),
    .B(_00966_),
    .Y(_01505_));
 sky130_fd_sc_hd__inv_2 _05461_ (.A(_01505_),
    .Y(_01516_));
 sky130_fd_sc_hd__nor2_1 _05462_ (.A(net54),
    .B(net22),
    .Y(_01527_));
 sky130_fd_sc_hd__or2_2 _05463_ (.A(net54),
    .B(net22),
    .X(_01538_));
 sky130_fd_sc_hd__and2_2 _05464_ (.A(net54),
    .B(net22),
    .X(_01549_));
 sky130_fd_sc_hd__nand2_1 _05465_ (.A(net54),
    .B(net22),
    .Y(_01560_));
 sky130_fd_sc_hd__nor2_1 _05466_ (.A(_01527_),
    .B(_01549_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_1 _05467_ (.A(net49),
    .B(net17),
    .Y(_01582_));
 sky130_fd_sc_hd__and2_1 _05468_ (.A(net49),
    .B(net17),
    .X(_01593_));
 sky130_fd_sc_hd__nor2_1 _05469_ (.A(_01582_),
    .B(_01593_),
    .Y(_01604_));
 sky130_fd_sc_hd__o22a_2 _05470_ (.A1(_01010_),
    .A2(net16),
    .B1(_01582_),
    .B2(_01593_),
    .X(_01615_));
 sky130_fd_sc_hd__o22ai_2 _05471_ (.A1(_01010_),
    .A2(net16),
    .B1(_01582_),
    .B2(_01593_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _05472_ (.A(_00999_),
    .B(net17),
    .Y(_01637_));
 sky130_fd_sc_hd__nor2_2 _05473_ (.A(net51),
    .B(net19),
    .Y(_01648_));
 sky130_fd_sc_hd__and2_2 _05474_ (.A(net51),
    .B(net19),
    .X(_01659_));
 sky130_fd_sc_hd__nor2_1 _05475_ (.A(_01648_),
    .B(_01659_),
    .Y(_01670_));
 sky130_fd_sc_hd__nor2_1 _05476_ (.A(net50),
    .B(net18),
    .Y(_01681_));
 sky130_fd_sc_hd__and2_1 _05477_ (.A(net50),
    .B(net18),
    .X(_01692_));
 sky130_fd_sc_hd__nor2_2 _05478_ (.A(_01681_),
    .B(_01692_),
    .Y(_01703_));
 sky130_fd_sc_hd__o22ai_2 _05479_ (.A1(_01648_),
    .A2(_01659_),
    .B1(_01681_),
    .B2(_01692_),
    .Y(_01714_));
 sky130_fd_sc_hd__a21oi_2 _05480_ (.A1(_01626_),
    .A2(_01637_),
    .B1(_01714_),
    .Y(_01725_));
 sky130_fd_sc_hd__and2b_1 _05481_ (.A_N(net50),
    .B(net18),
    .X(_01736_));
 sky130_fd_sc_hd__o21a_1 _05482_ (.A1(_01648_),
    .A2(_01659_),
    .B1(_01736_),
    .X(_01747_));
 sky130_fd_sc_hd__o21ai_1 _05483_ (.A1(_01648_),
    .A2(_01659_),
    .B1(_01736_),
    .Y(_01758_));
 sky130_fd_sc_hd__o21ai_2 _05484_ (.A1(net51),
    .A2(_00988_),
    .B1(_01758_),
    .Y(_01769_));
 sky130_fd_sc_hd__nor2_2 _05485_ (.A(_01769_),
    .B(_01725_),
    .Y(_01780_));
 sky130_fd_sc_hd__or2_1 _05486_ (.A(net52),
    .B(net20),
    .X(_01791_));
 sky130_fd_sc_hd__nand2_1 _05487_ (.A(net52),
    .B(net20),
    .Y(_01802_));
 sky130_fd_sc_hd__and2_2 _05488_ (.A(_01791_),
    .B(_01802_),
    .X(_01813_));
 sky130_fd_sc_hd__nor2_1 _05489_ (.A(net53),
    .B(net21),
    .Y(_01824_));
 sky130_fd_sc_hd__or2_1 _05490_ (.A(net53),
    .B(net21),
    .X(_01835_));
 sky130_fd_sc_hd__nand2_1 _05491_ (.A(net53),
    .B(net21),
    .Y(_01846_));
 sky130_fd_sc_hd__and2b_2 _05492_ (.A_N(_01824_),
    .B(_01846_),
    .X(_01857_));
 sky130_fd_sc_hd__a22o_1 _05493_ (.A1(_01791_),
    .A2(_01802_),
    .B1(_01835_),
    .B2(_01846_),
    .X(_01868_));
 sky130_fd_sc_hd__o21bai_4 _05494_ (.A1(_01769_),
    .A2(_01725_),
    .B1_N(_01868_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand2b_1 _05495_ (.A_N(net53),
    .B(net21),
    .Y(_01890_));
 sky130_fd_sc_hd__or2_2 _05496_ (.A(net52),
    .B(_00977_),
    .X(_01901_));
 sky130_fd_sc_hd__o31a_2 _05497_ (.A1(net52),
    .A2(_00977_),
    .A3(_01857_),
    .B1(_01890_),
    .X(_01912_));
 sky130_fd_sc_hd__a22oi_4 _05498_ (.A1(_01538_),
    .A2(_01560_),
    .B1(_01879_),
    .B2(_01912_),
    .Y(_01923_));
 sky130_fd_sc_hd__o2bb2ai_4 _05499_ (.A1_N(_01912_),
    .A2_N(_01879_),
    .B1(_01549_),
    .B2(_01527_),
    .Y(_01934_));
 sky130_fd_sc_hd__nor2_2 _05500_ (.A(net24),
    .B(net56),
    .Y(_01945_));
 sky130_fd_sc_hd__and2_2 _05501_ (.A(net24),
    .B(net56),
    .X(_01956_));
 sky130_fd_sc_hd__or2_4 _05502_ (.A(_01945_),
    .B(_01956_),
    .X(_01967_));
 sky130_fd_sc_hd__inv_2 _05503_ (.A(_01967_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor3_4 _05504_ (.A(_01505_),
    .B(_01967_),
    .C(_01923_),
    .Y(_01989_));
 sky130_fd_sc_hd__o211ai_4 _05505_ (.A1(net54),
    .A2(_00966_),
    .B1(_01978_),
    .C1(_01934_),
    .Y(_02000_));
 sky130_fd_sc_hd__a21oi_4 _05506_ (.A1(_01516_),
    .A2(_01934_),
    .B1(_01978_),
    .Y(_02011_));
 sky130_fd_sc_hd__o21ai_4 _05507_ (.A1(_01505_),
    .A2(_01923_),
    .B1(_01967_),
    .Y(_02022_));
 sky130_fd_sc_hd__o221a_4 _05508_ (.A1(net54),
    .A2(_00966_),
    .B1(_01945_),
    .B2(_01956_),
    .C1(_01934_),
    .X(_02033_));
 sky130_fd_sc_hd__o221ai_4 _05509_ (.A1(net54),
    .A2(_00966_),
    .B1(_01945_),
    .B2(_01956_),
    .C1(_01934_),
    .Y(_02044_));
 sky130_fd_sc_hd__a21oi_4 _05510_ (.A1(_01516_),
    .A2(_01934_),
    .B1(_01967_),
    .Y(_02055_));
 sky130_fd_sc_hd__o21bai_4 _05511_ (.A1(_01505_),
    .A2(_01923_),
    .B1_N(_01967_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_8 _05512_ (.A(_02044_),
    .B(net105),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_8 _05513_ (.A(_02000_),
    .B(_02022_),
    .Y(_02088_));
 sky130_fd_sc_hd__xor2_4 _05514_ (.A(_01780_),
    .B(_01813_),
    .X(_02099_));
 sky130_fd_sc_hd__nor2_4 _05515_ (.A(net48),
    .B(net16),
    .Y(_02110_));
 sky130_fd_sc_hd__and2_4 _05516_ (.A(net48),
    .B(net16),
    .X(_02121_));
 sky130_fd_sc_hd__nor2_8 _05517_ (.A(_02110_),
    .B(_02121_),
    .Y(_02132_));
 sky130_fd_sc_hd__or2_4 _05518_ (.A(_02110_),
    .B(_02121_),
    .X(_02143_));
 sky130_fd_sc_hd__o21ai_4 _05519_ (.A1(net48),
    .A2(_01021_),
    .B1(_01615_),
    .Y(_02154_));
 sky130_fd_sc_hd__or3_4 _05520_ (.A(_01604_),
    .B(_02132_),
    .C(_01714_),
    .X(_02165_));
 sky130_fd_sc_hd__o311a_4 _05521_ (.A1(_01670_),
    .A2(_01703_),
    .A3(_02154_),
    .B1(_02099_),
    .C1(_02077_),
    .X(_02176_));
 sky130_fd_sc_hd__a21oi_4 _05522_ (.A1(_02077_),
    .A2(_02165_),
    .B1(_02099_),
    .Y(_02187_));
 sky130_fd_sc_hd__or2_2 _05523_ (.A(_02176_),
    .B(_02187_),
    .X(_02198_));
 sky130_fd_sc_hd__nor2_4 _05524_ (.A(_02176_),
    .B(_02187_),
    .Y(_02209_));
 sky130_fd_sc_hd__and3_4 _05525_ (.A(net108),
    .B(net15),
    .C(net111),
    .X(_02220_));
 sky130_fd_sc_hd__nand3_4 _05526_ (.A(net108),
    .B(net15),
    .C(net111),
    .Y(_02231_));
 sky130_fd_sc_hd__nand3_4 _05527_ (.A(net105),
    .B(net47),
    .C(net107),
    .Y(_02242_));
 sky130_fd_sc_hd__o31a_1 _05528_ (.A1(_01032_),
    .A2(_01989_),
    .A3(net110),
    .B1(_02242_),
    .X(_02253_));
 sky130_fd_sc_hd__nand2_8 _05529_ (.A(_02231_),
    .B(_02242_),
    .Y(_02264_));
 sky130_fd_sc_hd__a21o_2 _05530_ (.A1(_01626_),
    .A2(_01637_),
    .B1(_01703_),
    .X(_02275_));
 sky130_fd_sc_hd__a2111o_2 _05531_ (.A1(net17),
    .A2(_00999_),
    .B1(_01681_),
    .C1(_01615_),
    .D1(_01692_),
    .X(_02286_));
 sky130_fd_sc_hd__nand2_1 _05532_ (.A(_02275_),
    .B(_02286_),
    .Y(_02297_));
 sky130_fd_sc_hd__and4_4 _05533_ (.A(_02077_),
    .B(_02154_),
    .C(_02275_),
    .D(_02286_),
    .X(_02308_));
 sky130_fd_sc_hd__a22oi_4 _05534_ (.A1(_02275_),
    .A2(_02286_),
    .B1(_02077_),
    .B2(_02154_),
    .Y(_02319_));
 sky130_fd_sc_hd__and3_4 _05535_ (.A(_02077_),
    .B(_02154_),
    .C(_02297_),
    .X(_02330_));
 sky130_fd_sc_hd__a21oi_4 _05536_ (.A1(_02077_),
    .A2(_02154_),
    .B1(_02297_),
    .Y(_02341_));
 sky130_fd_sc_hd__nor2_4 _05537_ (.A(_02308_),
    .B(_02319_),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_4 _05538_ (.A(_02330_),
    .B(_02341_),
    .Y(_02363_));
 sky130_fd_sc_hd__o221a_1 _05539_ (.A1(_02077_),
    .A2(_01043_),
    .B1(_02341_),
    .B2(_02330_),
    .C1(_02231_),
    .X(_02374_));
 sky130_fd_sc_hd__a311o_1 _05540_ (.A1(net47),
    .A2(net107),
    .A3(net105),
    .B1(_02220_),
    .C1(_02363_),
    .X(_02385_));
 sky130_fd_sc_hd__and3_1 _05541_ (.A(net48),
    .B(_01604_),
    .C(_01021_),
    .X(_02396_));
 sky130_fd_sc_hd__nor2_2 _05542_ (.A(_01615_),
    .B(_02396_),
    .Y(_02407_));
 sky130_fd_sc_hd__and4_4 _05543_ (.A(net111),
    .B(net108),
    .C(_02132_),
    .D(_02407_),
    .X(_02418_));
 sky130_fd_sc_hd__nand4_4 _05544_ (.A(net111),
    .B(net108),
    .C(_02132_),
    .D(_02407_),
    .Y(_02429_));
 sky130_fd_sc_hd__a21oi_4 _05545_ (.A1(_02077_),
    .A2(_02132_),
    .B1(_02407_),
    .Y(_02440_));
 sky130_fd_sc_hd__a31o_1 _05546_ (.A1(net111),
    .A2(net108),
    .A3(_02132_),
    .B1(_02407_),
    .X(_02451_));
 sky130_fd_sc_hd__nand2_8 _05547_ (.A(_02429_),
    .B(_02451_),
    .Y(_02462_));
 sky130_fd_sc_hd__nor2_8 _05548_ (.A(_02418_),
    .B(_02440_),
    .Y(_02473_));
 sky130_fd_sc_hd__o21ai_1 _05549_ (.A1(_02033_),
    .A2(_02055_),
    .B1(net14),
    .Y(_02484_));
 sky130_fd_sc_hd__o21ai_1 _05550_ (.A1(net113),
    .A2(net110),
    .B1(net46),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _05551_ (.A(_02484_),
    .B(_02495_),
    .Y(_02506_));
 sky130_fd_sc_hd__o2111ai_4 _05552_ (.A1(_01857_),
    .A2(_01901_),
    .B1(_01571_),
    .C1(_01890_),
    .D1(_01879_),
    .Y(_02517_));
 sky130_fd_sc_hd__nand2_4 _05553_ (.A(_01934_),
    .B(_02517_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand3b_4 _05554_ (.A_N(_02528_),
    .B(net105),
    .C(net107),
    .Y(_02539_));
 sky130_fd_sc_hd__o311a_2 _05555_ (.A1(_01813_),
    .A2(_01857_),
    .A3(_02165_),
    .B1(_02517_),
    .C1(_01934_),
    .X(_02550_));
 sky130_fd_sc_hd__o211ai_4 _05556_ (.A1(_01868_),
    .A2(_02165_),
    .B1(_02517_),
    .C1(_01934_),
    .Y(_02561_));
 sky130_fd_sc_hd__nand3_4 _05557_ (.A(net111),
    .B(net108),
    .C(_02561_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand3_4 _05558_ (.A(net106),
    .B(net104),
    .C(_02528_),
    .Y(_02583_));
 sky130_fd_sc_hd__nand3_4 _05559_ (.A(_02550_),
    .B(net108),
    .C(net111),
    .Y(_02594_));
 sky130_fd_sc_hd__nand2_4 _05560_ (.A(_02583_),
    .B(_02594_),
    .Y(_02605_));
 sky130_fd_sc_hd__nand2_8 _05561_ (.A(_02539_),
    .B(_02572_),
    .Y(_02616_));
 sky130_fd_sc_hd__o2111ai_1 _05562_ (.A1(_02077_),
    .A2(_02528_),
    .B1(_02572_),
    .C1(_02143_),
    .D1(_02506_),
    .Y(_02627_));
 sky130_fd_sc_hd__a32o_1 _05563_ (.A1(_02143_),
    .A2(_02539_),
    .A3(_02572_),
    .B1(_02231_),
    .B2(_02242_),
    .X(_02638_));
 sky130_fd_sc_hd__nand3_4 _05564_ (.A(_02242_),
    .B(_02583_),
    .C(_02594_),
    .Y(_02649_));
 sky130_fd_sc_hd__a21o_1 _05565_ (.A1(_02539_),
    .A2(_02572_),
    .B1(_02264_),
    .X(_02660_));
 sky130_fd_sc_hd__nand4_1 _05566_ (.A(_02484_),
    .B(_02495_),
    .C(_02539_),
    .D(_02572_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand3_1 _05567_ (.A(_02627_),
    .B(_02638_),
    .C(_02462_),
    .Y(_02682_));
 sky130_fd_sc_hd__o21ai_1 _05568_ (.A1(_02264_),
    .A2(_02462_),
    .B1(_02682_),
    .Y(_02693_));
 sky130_fd_sc_hd__a21oi_1 _05569_ (.A1(_02363_),
    .A2(_02693_),
    .B1(_02374_),
    .Y(_02704_));
 sky130_fd_sc_hd__and2b_1 _05570_ (.A_N(_01736_),
    .B(_02275_),
    .X(_02715_));
 sky130_fd_sc_hd__a211o_1 _05571_ (.A1(_01670_),
    .A2(_02715_),
    .B1(_01747_),
    .C1(_01725_),
    .X(_02726_));
 sky130_fd_sc_hd__a211o_1 _05572_ (.A1(_01010_),
    .A2(net16),
    .B1(_01703_),
    .C1(_01626_),
    .X(_02737_));
 sky130_fd_sc_hd__nand4_4 _05573_ (.A(_02000_),
    .B(_02022_),
    .C(_02726_),
    .D(_02737_),
    .Y(_02748_));
 sky130_fd_sc_hd__a31o_4 _05574_ (.A1(_02000_),
    .A2(_02022_),
    .A3(_02737_),
    .B1(_02726_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_4 _05575_ (.A(_02748_),
    .B(_02759_),
    .X(_02770_));
 sky130_fd_sc_hd__nand2_8 _05576_ (.A(_02748_),
    .B(_02759_),
    .Y(_02781_));
 sky130_fd_sc_hd__o311a_2 _05577_ (.A1(_01032_),
    .A2(_01989_),
    .A3(net110),
    .B1(_02242_),
    .C1(_02781_),
    .X(_02792_));
 sky130_fd_sc_hd__a221o_2 _05578_ (.A1(_02088_),
    .A2(net47),
    .B1(_02759_),
    .B2(_02748_),
    .C1(_02220_),
    .X(_02803_));
 sky130_fd_sc_hd__o21ai_1 _05579_ (.A1(_02781_),
    .A2(_02704_),
    .B1(_02803_),
    .Y(_02814_));
 sky130_fd_sc_hd__nand2_1 _05580_ (.A(_02209_),
    .B(_02814_),
    .Y(_02825_));
 sky130_fd_sc_hd__o211a_1 _05581_ (.A1(_01780_),
    .A2(_01813_),
    .B1(_01857_),
    .C1(_01901_),
    .X(_02836_));
 sky130_fd_sc_hd__o21ai_1 _05582_ (.A1(_01857_),
    .A2(_01901_),
    .B1(_01879_),
    .Y(_02847_));
 sky130_fd_sc_hd__or2_2 _05583_ (.A(_02847_),
    .B(_02836_),
    .X(_02858_));
 sky130_fd_sc_hd__o21ai_4 _05584_ (.A1(_02165_),
    .A2(_02099_),
    .B1(_02077_),
    .Y(_02869_));
 sky130_fd_sc_hd__nor2_2 _05585_ (.A(_02858_),
    .B(_02869_),
    .Y(_02880_));
 sky130_fd_sc_hd__or2_4 _05586_ (.A(_02858_),
    .B(_02869_),
    .X(_02891_));
 sky130_fd_sc_hd__and2_2 _05587_ (.A(_02869_),
    .B(_02858_),
    .X(_02902_));
 sky130_fd_sc_hd__nand2_4 _05588_ (.A(_02869_),
    .B(_02858_),
    .Y(_02913_));
 sky130_fd_sc_hd__nand2_8 _05589_ (.A(_02891_),
    .B(_02913_),
    .Y(_02924_));
 sky130_fd_sc_hd__nor2_4 _05590_ (.A(_02880_),
    .B(_02902_),
    .Y(_02935_));
 sky130_fd_sc_hd__o21ai_4 _05591_ (.A1(_02264_),
    .A2(_02605_),
    .B1(_02132_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand3_1 _05592_ (.A(_01087_),
    .B(net106),
    .C(net104),
    .Y(_02957_));
 sky130_fd_sc_hd__o31a_1 _05593_ (.A1(net6),
    .A2(net113),
    .A3(net110),
    .B1(_02957_),
    .X(_02968_));
 sky130_fd_sc_hd__o221ai_4 _05594_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_02968_),
    .C1(_02132_),
    .Y(_02979_));
 sky130_fd_sc_hd__o22ai_4 _05595_ (.A1(_02110_),
    .A2(_02121_),
    .B1(_02264_),
    .B2(_02605_),
    .Y(_02990_));
 sky130_fd_sc_hd__nand3b_1 _05596_ (.A_N(net37),
    .B(net106),
    .C(net104),
    .Y(_03001_));
 sky130_fd_sc_hd__o31a_1 _05597_ (.A1(net5),
    .A2(net113),
    .A3(net110),
    .B1(_03001_),
    .X(_03012_));
 sky130_fd_sc_hd__nor2_1 _05598_ (.A(_02616_),
    .B(_03012_),
    .Y(_03022_));
 sky130_fd_sc_hd__a21oi_1 _05599_ (.A1(net111),
    .A2(net108),
    .B1(net40),
    .Y(_03033_));
 sky130_fd_sc_hd__a21oi_1 _05600_ (.A1(net106),
    .A2(net104),
    .B1(net8),
    .Y(_03044_));
 sky130_fd_sc_hd__o2bb2a_2 _05601_ (.A1_N(_02583_),
    .A2_N(_02594_),
    .B1(_03033_),
    .B2(_03044_),
    .X(_03055_));
 sky130_fd_sc_hd__a21o_1 _05602_ (.A1(net111),
    .A2(net108),
    .B1(net39),
    .X(_03066_));
 sky130_fd_sc_hd__a21o_1 _05603_ (.A1(net106),
    .A2(net104),
    .B1(net7),
    .X(_03077_));
 sky130_fd_sc_hd__a21oi_4 _05604_ (.A1(_03066_),
    .A2(_03077_),
    .B1(_02616_),
    .Y(_03088_));
 sky130_fd_sc_hd__o221ai_4 _05605_ (.A1(_03088_),
    .A2(_02990_),
    .B1(_02946_),
    .B2(_03055_),
    .C1(_02473_),
    .Y(_03099_));
 sky130_fd_sc_hd__o211ai_2 _05606_ (.A1(_02990_),
    .A2(_03022_),
    .B1(_02462_),
    .C1(_02979_),
    .Y(_03110_));
 sky130_fd_sc_hd__o211ai_2 _05607_ (.A1(_02308_),
    .A2(_02319_),
    .B1(_03099_),
    .C1(_03110_),
    .Y(_03121_));
 sky130_fd_sc_hd__nand3_1 _05608_ (.A(_01076_),
    .B(net111),
    .C(net108),
    .Y(_03132_));
 sky130_fd_sc_hd__o31a_1 _05609_ (.A1(net41),
    .A2(_02033_),
    .A3(_02055_),
    .B1(_03132_),
    .X(_03143_));
 sky130_fd_sc_hd__o221a_1 _05610_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03143_),
    .C1(_02143_),
    .X(_03154_));
 sky130_fd_sc_hd__o221ai_2 _05611_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03143_),
    .C1(_02143_),
    .Y(_03165_));
 sky130_fd_sc_hd__a21o_1 _05612_ (.A1(net111),
    .A2(net108),
    .B1(net42),
    .X(_03176_));
 sky130_fd_sc_hd__nand3b_1 _05613_ (.A_N(net10),
    .B(net111),
    .C(net108),
    .Y(_03187_));
 sky130_fd_sc_hd__a22oi_4 _05614_ (.A1(_02583_),
    .A2(_02594_),
    .B1(_03176_),
    .B2(_03187_),
    .Y(_03198_));
 sky130_fd_sc_hd__nor2_1 _05615_ (.A(_03198_),
    .B(_02946_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand3_1 _05616_ (.A(_01054_),
    .B(net106),
    .C(net104),
    .Y(_03220_));
 sky130_fd_sc_hd__o31a_1 _05617_ (.A1(net13),
    .A2(net113),
    .A3(net110),
    .B1(_03220_),
    .X(_03231_));
 sky130_fd_sc_hd__o221ai_2 _05618_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03231_),
    .C1(_02132_),
    .Y(_03242_));
 sky130_fd_sc_hd__nand3_1 _05619_ (.A(_01065_),
    .B(net106),
    .C(net104),
    .Y(_03253_));
 sky130_fd_sc_hd__nand3b_1 _05620_ (.A_N(net11),
    .B(net111),
    .C(net108),
    .Y(_03264_));
 sky130_fd_sc_hd__o31a_1 _05621_ (.A1(net11),
    .A2(net113),
    .A3(net110),
    .B1(_03253_),
    .X(_03275_));
 sky130_fd_sc_hd__a22oi_2 _05622_ (.A1(_02583_),
    .A2(_02594_),
    .B1(_03253_),
    .B2(_03264_),
    .Y(_03286_));
 sky130_fd_sc_hd__o221ai_1 _05623_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03275_),
    .C1(_02143_),
    .Y(_03297_));
 sky130_fd_sc_hd__o211ai_2 _05624_ (.A1(_03286_),
    .A2(_02990_),
    .B1(_02473_),
    .C1(_03242_),
    .Y(_03308_));
 sky130_fd_sc_hd__o211ai_2 _05625_ (.A1(_03198_),
    .A2(_02946_),
    .B1(_02462_),
    .C1(_03165_),
    .Y(_03319_));
 sky130_fd_sc_hd__o211ai_2 _05626_ (.A1(_02330_),
    .A2(_02341_),
    .B1(_03308_),
    .C1(_03319_),
    .Y(_03330_));
 sky130_fd_sc_hd__o21a_2 _05627_ (.A1(_02176_),
    .A2(_02187_),
    .B1(_02781_),
    .X(_03341_));
 sky130_fd_sc_hd__a2bb2o_2 _05628_ (.A1_N(_02176_),
    .A2_N(_02187_),
    .B1(_02748_),
    .B2(_02759_),
    .X(_03352_));
 sky130_fd_sc_hd__a31oi_2 _05629_ (.A1(_03121_),
    .A2(_03330_),
    .A3(_03341_),
    .B1(_02935_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand3b_1 _05630_ (.A_N(net64),
    .B(net106),
    .C(net104),
    .Y(_03374_));
 sky130_fd_sc_hd__o31a_1 _05631_ (.A1(net32),
    .A2(net113),
    .A3(net110),
    .B1(_03374_),
    .X(_03385_));
 sky130_fd_sc_hd__o221ai_2 _05632_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03385_),
    .C1(_02143_),
    .Y(_03396_));
 sky130_fd_sc_hd__nand3b_1 _05633_ (.A_N(net34),
    .B(net106),
    .C(net104),
    .Y(_03407_));
 sky130_fd_sc_hd__o21ai_1 _05634_ (.A1(_02033_),
    .A2(_02055_),
    .B1(_01131_),
    .Y(_03418_));
 sky130_fd_sc_hd__o31a_1 _05635_ (.A1(net2),
    .A2(net113),
    .A3(net110),
    .B1(_03407_),
    .X(_03429_));
 sky130_fd_sc_hd__a21oi_1 _05636_ (.A1(_03407_),
    .A2(_03418_),
    .B1(_02616_),
    .Y(_03440_));
 sky130_fd_sc_hd__nand3b_2 _05637_ (.A_N(net36),
    .B(net106),
    .C(net104),
    .Y(_03451_));
 sky130_fd_sc_hd__nand3b_1 _05638_ (.A_N(net4),
    .B(net111),
    .C(net108),
    .Y(_03462_));
 sky130_fd_sc_hd__o31a_1 _05639_ (.A1(net4),
    .A2(net113),
    .A3(net110),
    .B1(_03451_),
    .X(_03473_));
 sky130_fd_sc_hd__a22oi_4 _05640_ (.A1(_02583_),
    .A2(_02594_),
    .B1(_03451_),
    .B2(_03462_),
    .Y(_03484_));
 sky130_fd_sc_hd__o221ai_1 _05641_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03473_),
    .C1(_02132_),
    .Y(_03495_));
 sky130_fd_sc_hd__o21ai_1 _05642_ (.A1(net113),
    .A2(net110),
    .B1(_01109_),
    .Y(_03506_));
 sky130_fd_sc_hd__o21ai_1 _05643_ (.A1(_02033_),
    .A2(_02055_),
    .B1(_01120_),
    .Y(_03517_));
 sky130_fd_sc_hd__a22oi_4 _05644_ (.A1(_02583_),
    .A2(_02594_),
    .B1(_03506_),
    .B2(_03517_),
    .Y(_03528_));
 sky130_fd_sc_hd__o211ai_1 _05645_ (.A1(_03528_),
    .A2(_02990_),
    .B1(_02473_),
    .C1(_03495_),
    .Y(_03539_));
 sky130_fd_sc_hd__o211ai_1 _05646_ (.A1(_03440_),
    .A2(_02946_),
    .B1(_02462_),
    .C1(_03396_),
    .Y(_03550_));
 sky130_fd_sc_hd__and3_1 _05647_ (.A(_03550_),
    .B(_02352_),
    .C(_03539_),
    .X(_03561_));
 sky130_fd_sc_hd__and3_1 _05648_ (.A(_02198_),
    .B(_02748_),
    .C(_02759_),
    .X(_03572_));
 sky130_fd_sc_hd__o21ai_2 _05649_ (.A1(_02176_),
    .A2(_02187_),
    .B1(_02770_),
    .Y(_03583_));
 sky130_fd_sc_hd__a21o_1 _05650_ (.A1(net111),
    .A2(net108),
    .B1(net61),
    .X(_03594_));
 sky130_fd_sc_hd__nand3_1 _05651_ (.A(_01186_),
    .B(net111),
    .C(net108),
    .Y(_03605_));
 sky130_fd_sc_hd__a22oi_4 _05652_ (.A1(_02583_),
    .A2(_02594_),
    .B1(_03594_),
    .B2(_03605_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand3_1 _05653_ (.A(_01197_),
    .B(net106),
    .C(net104),
    .Y(_03627_));
 sky130_fd_sc_hd__o31a_1 _05654_ (.A1(net28),
    .A2(net113),
    .A3(net110),
    .B1(_03627_),
    .X(_03638_));
 sky130_fd_sc_hd__o221ai_4 _05655_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03638_),
    .C1(_02143_),
    .Y(_03649_));
 sky130_fd_sc_hd__o21ai_1 _05656_ (.A1(net113),
    .A2(net110),
    .B1(_01142_),
    .Y(_03660_));
 sky130_fd_sc_hd__o21ai_1 _05657_ (.A1(_02033_),
    .A2(_02055_),
    .B1(_01153_),
    .Y(_03671_));
 sky130_fd_sc_hd__a21oi_2 _05658_ (.A1(_03660_),
    .A2(_03671_),
    .B1(_02616_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand3_1 _05659_ (.A(_01164_),
    .B(net106),
    .C(net104),
    .Y(_03693_));
 sky130_fd_sc_hd__o31a_1 _05660_ (.A1(net30),
    .A2(net113),
    .A3(net110),
    .B1(_03693_),
    .X(_03704_));
 sky130_fd_sc_hd__o221ai_2 _05661_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03704_),
    .C1(_02143_),
    .Y(_03715_));
 sky130_fd_sc_hd__o21ai_1 _05662_ (.A1(_03682_),
    .A2(_02946_),
    .B1(_03715_),
    .Y(_03726_));
 sky130_fd_sc_hd__o211ai_1 _05663_ (.A1(_03682_),
    .A2(_02946_),
    .B1(_02473_),
    .C1(_03715_),
    .Y(_03737_));
 sky130_fd_sc_hd__o211ai_1 _05664_ (.A1(_03616_),
    .A2(_02946_),
    .B1(_02462_),
    .C1(_03649_),
    .Y(_03748_));
 sky130_fd_sc_hd__a31o_1 _05665_ (.A1(_02363_),
    .A2(_03737_),
    .A3(_03748_),
    .B1(_03583_),
    .X(_03759_));
 sky130_fd_sc_hd__o211ai_4 _05666_ (.A1(_03561_),
    .A2(_03759_),
    .B1(_03363_),
    .C1(_02825_),
    .Y(_03770_));
 sky130_fd_sc_hd__and3_1 _05667_ (.A(_02264_),
    .B(_02891_),
    .C(_02913_),
    .X(_03781_));
 sky130_fd_sc_hd__o32a_2 _05668_ (.A1(_02253_),
    .A2(_02880_),
    .A3(_02902_),
    .B1(net110),
    .B2(_01989_),
    .X(_03792_));
 sky130_fd_sc_hd__a31o_1 _05669_ (.A1(_02264_),
    .A2(_02891_),
    .A3(_02913_),
    .B1(_02077_),
    .X(_03803_));
 sky130_fd_sc_hd__o2bb2a_2 _05670_ (.A1_N(_03792_),
    .A2_N(_03770_),
    .B1(_02088_),
    .B2(net60),
    .X(_03814_));
 sky130_fd_sc_hd__inv_2 _05671_ (.A(_03814_),
    .Y(_03825_));
 sky130_fd_sc_hd__a21oi_1 _05672_ (.A1(net112),
    .A2(net109),
    .B1(net28),
    .Y(_03836_));
 sky130_fd_sc_hd__o32a_4 _05673_ (.A1(_02253_),
    .A2(_02880_),
    .A3(_02902_),
    .B1(_02055_),
    .B2(_02033_),
    .X(_03847_));
 sky130_fd_sc_hd__a31o_1 _05674_ (.A1(_02264_),
    .A2(_02891_),
    .A3(_02913_),
    .B1(_02088_),
    .X(_03858_));
 sky130_fd_sc_hd__o211a_1 _05675_ (.A1(_01032_),
    .A2(_02924_),
    .B1(_02077_),
    .C1(_03770_),
    .X(_03869_));
 sky130_fd_sc_hd__o2bb2a_2 _05676_ (.A1_N(_03847_),
    .A2_N(_03770_),
    .B1(_02077_),
    .B2(net28),
    .X(_03880_));
 sky130_fd_sc_hd__inv_2 _05677_ (.A(_03880_),
    .Y(_03891_));
 sky130_fd_sc_hd__o22a_2 _05678_ (.A1(_02033_),
    .A2(_02055_),
    .B1(_02264_),
    .B2(_02924_),
    .X(_03902_));
 sky130_fd_sc_hd__a31o_1 _05679_ (.A1(_01032_),
    .A2(_02242_),
    .A3(_02935_),
    .B1(_02088_),
    .X(_03913_));
 sky130_fd_sc_hd__o211ai_2 _05680_ (.A1(_02264_),
    .A2(_02605_),
    .B1(_02132_),
    .C1(_02671_),
    .Y(_03924_));
 sky130_fd_sc_hd__o221ai_4 _05681_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03231_),
    .C1(_02143_),
    .Y(_03935_));
 sky130_fd_sc_hd__o211ai_2 _05682_ (.A1(_02418_),
    .A2(_02440_),
    .B1(_03924_),
    .C1(_03935_),
    .Y(_03946_));
 sky130_fd_sc_hd__o31a_1 _05683_ (.A1(_02264_),
    .A2(_02418_),
    .A3(_02440_),
    .B1(_03946_),
    .X(_03956_));
 sky130_fd_sc_hd__o21ai_2 _05684_ (.A1(_02352_),
    .A2(_03956_),
    .B1(_02385_),
    .Y(_03965_));
 sky130_fd_sc_hd__o21a_1 _05685_ (.A1(_02264_),
    .A2(_02770_),
    .B1(_02209_),
    .X(_03975_));
 sky130_fd_sc_hd__a211o_1 _05686_ (.A1(_03965_),
    .A2(_02770_),
    .B1(_02198_),
    .C1(_02792_),
    .X(_03984_));
 sky130_fd_sc_hd__o221ai_1 _05687_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03012_),
    .C1(_02132_),
    .Y(_03993_));
 sky130_fd_sc_hd__o22a_1 _05688_ (.A1(_03484_),
    .A2(_02990_),
    .B1(_02946_),
    .B2(_03022_),
    .X(_04003_));
 sky130_fd_sc_hd__o221ai_2 _05689_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_02968_),
    .C1(_02143_),
    .Y(_04012_));
 sky130_fd_sc_hd__o211ai_1 _05690_ (.A1(_03088_),
    .A2(_02946_),
    .B1(_02473_),
    .C1(_04012_),
    .Y(_04021_));
 sky130_fd_sc_hd__o211ai_1 _05691_ (.A1(_03484_),
    .A2(_02990_),
    .B1(_02462_),
    .C1(_03993_),
    .Y(_04031_));
 sky130_fd_sc_hd__o221ai_2 _05692_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03143_),
    .C1(_02132_),
    .Y(_04040_));
 sky130_fd_sc_hd__o21ai_1 _05693_ (.A1(_02990_),
    .A2(_03055_),
    .B1(_04040_),
    .Y(_04050_));
 sky130_fd_sc_hd__o221ai_4 _05694_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03275_),
    .C1(_02132_),
    .Y(_04060_));
 sky130_fd_sc_hd__o211ai_2 _05695_ (.A1(_03198_),
    .A2(_02990_),
    .B1(_02473_),
    .C1(_04060_),
    .Y(_04069_));
 sky130_fd_sc_hd__o211ai_1 _05696_ (.A1(_02990_),
    .A2(_03055_),
    .B1(_02462_),
    .C1(_04040_),
    .Y(_04079_));
 sky130_fd_sc_hd__o221a_1 _05697_ (.A1(_02330_),
    .A2(_02341_),
    .B1(_02473_),
    .B2(_04050_),
    .C1(_04069_),
    .X(_04088_));
 sky130_fd_sc_hd__a31o_1 _05698_ (.A1(_02363_),
    .A2(_04021_),
    .A3(_04031_),
    .B1(_04088_),
    .X(_04099_));
 sky130_fd_sc_hd__nand2_1 _05699_ (.A(_04099_),
    .B(_03341_),
    .Y(_04110_));
 sky130_fd_sc_hd__o221ai_2 _05700_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03385_),
    .C1(_02132_),
    .Y(_04121_));
 sky130_fd_sc_hd__o221ai_2 _05701_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03429_),
    .C1(_02143_),
    .Y(_04132_));
 sky130_fd_sc_hd__o21ai_1 _05702_ (.A1(_03528_),
    .A2(_02946_),
    .B1(_04132_),
    .Y(_04143_));
 sky130_fd_sc_hd__o211ai_1 _05703_ (.A1(_03528_),
    .A2(_02946_),
    .B1(_02473_),
    .C1(_04132_),
    .Y(_04153_));
 sky130_fd_sc_hd__o211ai_2 _05704_ (.A1(_03682_),
    .A2(_02990_),
    .B1(_02462_),
    .C1(_04121_),
    .Y(_04164_));
 sky130_fd_sc_hd__o21ai_1 _05705_ (.A1(_02462_),
    .A2(_04143_),
    .B1(_04164_),
    .Y(_04175_));
 sky130_fd_sc_hd__o221ai_2 _05706_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03638_),
    .C1(_02132_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand3b_1 _05707_ (.A_N(net59),
    .B(net106),
    .C(net104),
    .Y(_04197_));
 sky130_fd_sc_hd__nand3_1 _05708_ (.A(_01208_),
    .B(net111),
    .C(net108),
    .Y(_04208_));
 sky130_fd_sc_hd__o31a_1 _05709_ (.A1(net27),
    .A2(net113),
    .A3(net110),
    .B1(_04197_),
    .X(_04219_));
 sky130_fd_sc_hd__a21oi_1 _05710_ (.A1(_04197_),
    .A2(_04208_),
    .B1(_02616_),
    .Y(_04230_));
 sky130_fd_sc_hd__o221ai_2 _05711_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_03704_),
    .C1(_02132_),
    .Y(_04241_));
 sky130_fd_sc_hd__o211ai_1 _05712_ (.A1(_03616_),
    .A2(_02990_),
    .B1(_02473_),
    .C1(_04241_),
    .Y(_04252_));
 sky130_fd_sc_hd__o211ai_1 _05713_ (.A1(_04230_),
    .A2(_02990_),
    .B1(_02462_),
    .C1(_04186_),
    .Y(_04262_));
 sky130_fd_sc_hd__a21oi_1 _05714_ (.A1(_04252_),
    .A2(_04262_),
    .B1(_02352_),
    .Y(_04273_));
 sky130_fd_sc_hd__a211o_1 _05715_ (.A1(_02352_),
    .A2(_04175_),
    .B1(_03583_),
    .C1(_04273_),
    .X(_04284_));
 sky130_fd_sc_hd__nand4_4 _05716_ (.A(_03984_),
    .B(_04110_),
    .C(_04284_),
    .D(_02924_),
    .Y(_04295_));
 sky130_fd_sc_hd__o2bb2a_1 _05717_ (.A1_N(_04295_),
    .A2_N(_03902_),
    .B1(_02077_),
    .B2(_01208_),
    .X(_04306_));
 sky130_fd_sc_hd__a32o_2 _05718_ (.A1(net27),
    .A2(net107),
    .A3(net105),
    .B1(_04295_),
    .B2(_03902_),
    .X(_04317_));
 sky130_fd_sc_hd__o311a_2 _05719_ (.A1(net47),
    .A2(_02220_),
    .A3(_02924_),
    .B1(net106),
    .C1(net104),
    .X(_04328_));
 sky130_fd_sc_hd__a32o_4 _05720_ (.A1(net59),
    .A2(net112),
    .A3(net109),
    .B1(_04295_),
    .B2(_04328_),
    .X(_04339_));
 sky130_fd_sc_hd__a21oi_1 _05721_ (.A1(_02627_),
    .A2(_02638_),
    .B1(_02462_),
    .Y(_04350_));
 sky130_fd_sc_hd__a21oi_1 _05722_ (.A1(_03242_),
    .A2(_03297_),
    .B1(_02473_),
    .Y(_04361_));
 sky130_fd_sc_hd__o31a_1 _05723_ (.A1(_02352_),
    .A2(_04350_),
    .A3(_04361_),
    .B1(_02385_),
    .X(_04371_));
 sky130_fd_sc_hd__o21ai_2 _05724_ (.A1(_02781_),
    .A2(_04371_),
    .B1(_02803_),
    .Y(_04382_));
 sky130_fd_sc_hd__o211ai_1 _05725_ (.A1(_03440_),
    .A2(_02946_),
    .B1(_02473_),
    .C1(_03396_),
    .Y(_04393_));
 sky130_fd_sc_hd__o21a_1 _05726_ (.A1(_02473_),
    .A2(_03726_),
    .B1(_04393_),
    .X(_04404_));
 sky130_fd_sc_hd__o221a_1 _05727_ (.A1(_02330_),
    .A2(_02341_),
    .B1(_02473_),
    .B2(_03726_),
    .C1(_04393_),
    .X(_04415_));
 sky130_fd_sc_hd__o211ai_1 _05728_ (.A1(_03616_),
    .A2(_02946_),
    .B1(_02473_),
    .C1(_03649_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand3b_1 _05729_ (.A_N(net58),
    .B(net106),
    .C(net104),
    .Y(_04437_));
 sky130_fd_sc_hd__o31a_1 _05730_ (.A1(net26),
    .A2(net113),
    .A3(net110),
    .B1(_04437_),
    .X(_04448_));
 sky130_fd_sc_hd__o31ai_1 _05731_ (.A1(net26),
    .A2(net113),
    .A3(net110),
    .B1(_04437_),
    .Y(_04459_));
 sky130_fd_sc_hd__o221ai_2 _05732_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_04448_),
    .C1(_02143_),
    .Y(_04470_));
 sky130_fd_sc_hd__o221ai_2 _05733_ (.A1(_02220_),
    .A2(_02649_),
    .B1(_02616_),
    .B2(_04219_),
    .C1(_02132_),
    .Y(_04481_));
 sky130_fd_sc_hd__o211ai_1 _05734_ (.A1(_02418_),
    .A2(_02440_),
    .B1(_04470_),
    .C1(_04481_),
    .Y(_04492_));
 sky130_fd_sc_hd__a31o_1 _05735_ (.A1(_02363_),
    .A2(_04426_),
    .A3(_04492_),
    .B1(_03583_),
    .X(_04503_));
 sky130_fd_sc_hd__o221ai_2 _05736_ (.A1(_03528_),
    .A2(_02990_),
    .B1(_03484_),
    .B2(_02946_),
    .C1(_02462_),
    .Y(_04514_));
 sky130_fd_sc_hd__o211ai_1 _05737_ (.A1(_02990_),
    .A2(_03022_),
    .B1(_02473_),
    .C1(_02979_),
    .Y(_04524_));
 sky130_fd_sc_hd__o211ai_1 _05738_ (.A1(_02308_),
    .A2(_02319_),
    .B1(_04514_),
    .C1(_04524_),
    .Y(_04535_));
 sky130_fd_sc_hd__o221ai_4 _05739_ (.A1(_03088_),
    .A2(_02990_),
    .B1(_02946_),
    .B2(_03055_),
    .C1(_02462_),
    .Y(_04546_));
 sky130_fd_sc_hd__o31a_1 _05740_ (.A1(_02462_),
    .A2(_03154_),
    .A3(_03209_),
    .B1(_04546_),
    .X(_04557_));
 sky130_fd_sc_hd__o311ai_2 _05741_ (.A1(_02462_),
    .A2(_03154_),
    .A3(_03209_),
    .B1(_04546_),
    .C1(_02352_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand4_1 _05742_ (.A(_02781_),
    .B(_04535_),
    .C(_04568_),
    .D(_02198_),
    .Y(_04579_));
 sky130_fd_sc_hd__o211ai_2 _05743_ (.A1(_04415_),
    .A2(_04503_),
    .B1(_02924_),
    .C1(_04579_),
    .Y(_04590_));
 sky130_fd_sc_hd__a21oi_4 _05744_ (.A1(_02209_),
    .A2(_04382_),
    .B1(_04590_),
    .Y(_04601_));
 sky130_fd_sc_hd__o22ai_4 _05745_ (.A1(net58),
    .A2(_02088_),
    .B1(_03803_),
    .B2(_04601_),
    .Y(_04612_));
 sky130_fd_sc_hd__inv_2 _05746_ (.A(_04612_),
    .Y(_04623_));
 sky130_fd_sc_hd__o32a_4 _05747_ (.A1(net26),
    .A2(_02033_),
    .A3(_02055_),
    .B1(_03858_),
    .B2(_04601_),
    .X(_04634_));
 sky130_fd_sc_hd__o22ai_4 _05748_ (.A1(net26),
    .A2(_02077_),
    .B1(_03858_),
    .B2(_04601_),
    .Y(_04645_));
 sky130_fd_sc_hd__nand3_1 _05749_ (.A(_03099_),
    .B(_03110_),
    .C(_02352_),
    .Y(_04655_));
 sky130_fd_sc_hd__o211ai_1 _05750_ (.A1(_02308_),
    .A2(_02319_),
    .B1(_03539_),
    .C1(_03550_),
    .Y(_04666_));
 sky130_fd_sc_hd__nand2_2 _05751_ (.A(_04655_),
    .B(_04666_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand3_1 _05752_ (.A(_01252_),
    .B(net106),
    .C(net104),
    .Y(_04688_));
 sky130_fd_sc_hd__o31ai_2 _05753_ (.A1(net12),
    .A2(net113),
    .A3(net110),
    .B1(_04688_),
    .Y(_04699_));
 sky130_fd_sc_hd__o2111ai_1 _05754_ (.A1(_02528_),
    .A2(_02077_),
    .B1(_02143_),
    .C1(_02572_),
    .D1(_04699_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand3_1 _05755_ (.A(_01230_),
    .B(net106),
    .C(net104),
    .Y(_04721_));
 sky130_fd_sc_hd__o31ai_2 _05756_ (.A1(net23),
    .A2(net113),
    .A3(net110),
    .B1(_04721_),
    .Y(_04732_));
 sky130_fd_sc_hd__nand2_1 _05757_ (.A(_04732_),
    .B(_02605_),
    .Y(_04743_));
 sky130_fd_sc_hd__o2111a_1 _05758_ (.A1(_02143_),
    .A2(_04743_),
    .B1(_04710_),
    .C1(_02660_),
    .D1(_02462_),
    .X(_04754_));
 sky130_fd_sc_hd__a21oi_1 _05759_ (.A1(_04470_),
    .A2(_04481_),
    .B1(_02462_),
    .Y(_04765_));
 sky130_fd_sc_hd__o21ai_1 _05760_ (.A1(_04754_),
    .A2(_04765_),
    .B1(_02363_),
    .Y(_04775_));
 sky130_fd_sc_hd__a31oi_1 _05761_ (.A1(_03737_),
    .A2(_03748_),
    .A3(_02352_),
    .B1(_03583_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2_1 _05762_ (.A(_04786_),
    .B(_04775_),
    .Y(_04797_));
 sky130_fd_sc_hd__o2bb2ai_1 _05763_ (.A1_N(_04775_),
    .A2_N(_04786_),
    .B1(_03352_),
    .B2(_04677_),
    .Y(_04808_));
 sky130_fd_sc_hd__o22a_4 _05764_ (.A1(_02176_),
    .A2(_02187_),
    .B1(_02880_),
    .B2(_02902_),
    .X(_04819_));
 sky130_fd_sc_hd__a2bb2o_2 _05765_ (.A1_N(_02176_),
    .A2_N(_02187_),
    .B1(_02891_),
    .B2(_02913_),
    .X(_04830_));
 sky130_fd_sc_hd__o211ai_2 _05766_ (.A1(_02308_),
    .A2(_02319_),
    .B1(_03308_),
    .C1(_03319_),
    .Y(_04841_));
 sky130_fd_sc_hd__o211ai_1 _05767_ (.A1(_02264_),
    .A2(_02462_),
    .B1(_02352_),
    .C1(_02682_),
    .Y(_04852_));
 sky130_fd_sc_hd__nand3_2 _05768_ (.A(_04841_),
    .B(_04852_),
    .C(_02770_),
    .Y(_04862_));
 sky130_fd_sc_hd__o22a_1 _05769_ (.A1(_02880_),
    .A2(_02902_),
    .B1(_02264_),
    .B2(_02770_),
    .X(_04873_));
 sky130_fd_sc_hd__nand2_1 _05770_ (.A(_04862_),
    .B(_04873_),
    .Y(_04884_));
 sky130_fd_sc_hd__o2bb2ai_1 _05771_ (.A1_N(_04873_),
    .A2_N(_04862_),
    .B1(_02935_),
    .B2(_02209_),
    .Y(_04895_));
 sky130_fd_sc_hd__a21oi_1 _05772_ (.A1(_02803_),
    .A2(_04862_),
    .B1(_02198_),
    .Y(_04906_));
 sky130_fd_sc_hd__o211ai_1 _05773_ (.A1(_03352_),
    .A2(_04677_),
    .B1(_02924_),
    .C1(_04797_),
    .Y(_04917_));
 sky130_fd_sc_hd__a21oi_1 _05774_ (.A1(_04830_),
    .A2(_04884_),
    .B1(_04808_),
    .Y(_04923_));
 sky130_fd_sc_hd__o211ai_4 _05775_ (.A1(_03352_),
    .A2(_04677_),
    .B1(_04797_),
    .C1(_04895_),
    .Y(_04930_));
 sky130_fd_sc_hd__o21ai_2 _05776_ (.A1(_03781_),
    .A2(_04923_),
    .B1(_02088_),
    .Y(_04936_));
 sky130_fd_sc_hd__or3_1 _05777_ (.A(_01252_),
    .B(_01989_),
    .C(net110),
    .X(_04943_));
 sky130_fd_sc_hd__a22oi_4 _05778_ (.A1(_01252_),
    .A2(_02077_),
    .B1(_04930_),
    .B2(_03792_),
    .Y(_04949_));
 sky130_fd_sc_hd__a32o_1 _05779_ (.A1(_01252_),
    .A2(net112),
    .A3(net109),
    .B1(_04930_),
    .B2(_03792_),
    .X(_04956_));
 sky130_fd_sc_hd__o21ai_1 _05780_ (.A1(_04906_),
    .A2(_04917_),
    .B1(_03847_),
    .Y(_04962_));
 sky130_fd_sc_hd__or3_1 _05781_ (.A(net12),
    .B(_02033_),
    .C(_02055_),
    .X(_04969_));
 sky130_fd_sc_hd__o22a_1 _05782_ (.A1(net12),
    .A2(_02077_),
    .B1(_03858_),
    .B2(_04923_),
    .X(_04975_));
 sky130_fd_sc_hd__a22o_2 _05783_ (.A1(_01241_),
    .A2(_02088_),
    .B1(_04930_),
    .B2(_03847_),
    .X(_04979_));
 sky130_fd_sc_hd__o221ai_4 _05784_ (.A1(_02330_),
    .A2(_02341_),
    .B1(_02462_),
    .B2(_02264_),
    .C1(_03946_),
    .Y(_04980_));
 sky130_fd_sc_hd__o211ai_2 _05785_ (.A1(_02308_),
    .A2(_02319_),
    .B1(_04069_),
    .C1(_04079_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand3_1 _05786_ (.A(_04981_),
    .B(_02770_),
    .C(_04980_),
    .Y(_04982_));
 sky130_fd_sc_hd__a31oi_2 _05787_ (.A1(_04981_),
    .A2(_02770_),
    .A3(_04980_),
    .B1(_02792_),
    .Y(_04983_));
 sky130_fd_sc_hd__a21oi_1 _05788_ (.A1(_02803_),
    .A2(_04982_),
    .B1(_02198_),
    .Y(_04984_));
 sky130_fd_sc_hd__o211ai_2 _05789_ (.A1(_02308_),
    .A2(_02319_),
    .B1(_04153_),
    .C1(_04164_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand3_1 _05790_ (.A(_04021_),
    .B(_04031_),
    .C(_02352_),
    .Y(_04986_));
 sky130_fd_sc_hd__o21ai_1 _05791_ (.A1(_02352_),
    .A2(_04175_),
    .B1(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__a22oi_4 _05792_ (.A1(_02748_),
    .A2(_02759_),
    .B1(_04985_),
    .B2(_04986_),
    .Y(_04988_));
 sky130_fd_sc_hd__a2bb2oi_1 _05793_ (.A1_N(_02330_),
    .A2_N(_02341_),
    .B1(_04252_),
    .B2(_04262_),
    .Y(_04989_));
 sky130_fd_sc_hd__o2111ai_2 _05794_ (.A1(_02077_),
    .A2(_02528_),
    .B1(_02572_),
    .C1(_02132_),
    .D1(_04459_),
    .Y(_04990_));
 sky130_fd_sc_hd__o211ai_1 _05795_ (.A1(_02110_),
    .A2(_02121_),
    .B1(_02605_),
    .C1(_04732_),
    .Y(_04991_));
 sky130_fd_sc_hd__nand3_1 _05796_ (.A(_02660_),
    .B(_04990_),
    .C(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__nand4_1 _05797_ (.A(_02473_),
    .B(_02660_),
    .C(_04990_),
    .D(_04991_),
    .Y(_04993_));
 sky130_fd_sc_hd__nand3b_1 _05798_ (.A_N(net33),
    .B(net106),
    .C(net104),
    .Y(_04994_));
 sky130_fd_sc_hd__o31ai_1 _05799_ (.A1(net1),
    .A2(net113),
    .A3(net110),
    .B1(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__o2111ai_1 _05800_ (.A1(_02528_),
    .A2(_02077_),
    .B1(_02143_),
    .C1(_02572_),
    .D1(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand3_1 _05801_ (.A(_04699_),
    .B(_02605_),
    .C(_02132_),
    .Y(_04997_));
 sky130_fd_sc_hd__nand4_1 _05802_ (.A(_02660_),
    .B(_04996_),
    .C(_04997_),
    .D(_02462_),
    .Y(_04998_));
 sky130_fd_sc_hd__a31o_1 _05803_ (.A1(_02363_),
    .A2(_04993_),
    .A3(_04998_),
    .B1(_02781_),
    .X(_04999_));
 sky130_fd_sc_hd__o22ai_4 _05804_ (.A1(_02176_),
    .A2(_02187_),
    .B1(_04989_),
    .B2(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__o22ai_1 _05805_ (.A1(_02880_),
    .A2(_02902_),
    .B1(_04988_),
    .B2(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__o221ai_4 _05806_ (.A1(_04988_),
    .A2(_05000_),
    .B1(_02198_),
    .B2(_04983_),
    .C1(_02924_),
    .Y(_05002_));
 sky130_fd_sc_hd__o2bb2ai_4 _05807_ (.A1_N(_03847_),
    .A2_N(_05002_),
    .B1(net1),
    .B2(_02077_),
    .Y(_05003_));
 sky130_fd_sc_hd__inv_2 _05808_ (.A(_05003_),
    .Y(\adder_inst.fraction1[0] ));
 sky130_fd_sc_hd__o21bai_2 _05809_ (.A1(_04984_),
    .A2(_05001_),
    .B1_N(_03803_),
    .Y(_05004_));
 sky130_fd_sc_hd__or3_1 _05810_ (.A(net33),
    .B(_01989_),
    .C(net110),
    .X(_05005_));
 sky130_fd_sc_hd__a2bb2o_1 _05811_ (.A1_N(net33),
    .A2_N(_02088_),
    .B1(_03792_),
    .B2(_05002_),
    .X(_05006_));
 sky130_fd_sc_hd__inv_2 _05812_ (.A(_05006_),
    .Y(\adder_inst.fraction2[0] ));
 sky130_fd_sc_hd__o22a_1 _05813_ (.A1(_05003_),
    .A2(\adder_inst.fraction2[0] ),
    .B1(_04949_),
    .B2(_04979_),
    .X(_05007_));
 sky130_fd_sc_hd__and3_1 _05814_ (.A(net105),
    .B(net23),
    .C(net107),
    .X(_05008_));
 sky130_fd_sc_hd__o21ai_1 _05815_ (.A1(_01989_),
    .A2(net110),
    .B1(net23),
    .Y(_05009_));
 sky130_fd_sc_hd__o211ai_1 _05816_ (.A1(_03198_),
    .A2(_02990_),
    .B1(_02462_),
    .C1(_04060_),
    .Y(_05010_));
 sky130_fd_sc_hd__nand3_1 _05817_ (.A(_02473_),
    .B(_03924_),
    .C(_03935_),
    .Y(_05011_));
 sky130_fd_sc_hd__a2bb2oi_1 _05818_ (.A1_N(_02308_),
    .A2_N(_02319_),
    .B1(_05010_),
    .B2(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__o21bai_1 _05819_ (.A1(_02374_),
    .A2(_05012_),
    .B1_N(_02781_),
    .Y(_05013_));
 sky130_fd_sc_hd__nand2_2 _05820_ (.A(_05013_),
    .B(_03975_),
    .Y(_05014_));
 sky130_fd_sc_hd__o21ai_2 _05821_ (.A1(_02418_),
    .A2(_02440_),
    .B1(_04143_),
    .Y(_05015_));
 sky130_fd_sc_hd__o221ai_4 _05822_ (.A1(_02308_),
    .A2(_02319_),
    .B1(_02462_),
    .B2(_04003_),
    .C1(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__o211ai_1 _05823_ (.A1(_03088_),
    .A2(_02946_),
    .B1(_02462_),
    .C1(_04012_),
    .Y(_05017_));
 sky130_fd_sc_hd__o21a_1 _05824_ (.A1(_02462_),
    .A2(_04050_),
    .B1(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__o21ai_2 _05825_ (.A1(_02363_),
    .A2(_05018_),
    .B1(_05016_),
    .Y(_05019_));
 sky130_fd_sc_hd__o211ai_4 _05826_ (.A1(_02363_),
    .A2(_05018_),
    .B1(_05016_),
    .C1(_03341_),
    .Y(_05020_));
 sky130_fd_sc_hd__o211a_1 _05827_ (.A1(_04230_),
    .A2(_02990_),
    .B1(_02473_),
    .C1(_04186_),
    .X(_05021_));
 sky130_fd_sc_hd__o2bb2ai_1 _05828_ (.A1_N(_02462_),
    .A2_N(_04992_),
    .B1(_02308_),
    .B2(_02319_),
    .Y(_05022_));
 sky130_fd_sc_hd__o211ai_1 _05829_ (.A1(_03616_),
    .A2(_02990_),
    .B1(_02462_),
    .C1(_04241_),
    .Y(_05023_));
 sky130_fd_sc_hd__o211ai_1 _05830_ (.A1(_03682_),
    .A2(_02990_),
    .B1(_02473_),
    .C1(_04121_),
    .Y(_05024_));
 sky130_fd_sc_hd__o211ai_1 _05831_ (.A1(_02330_),
    .A2(_02341_),
    .B1(_05023_),
    .C1(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__o21ai_2 _05832_ (.A1(_05021_),
    .A2(_05022_),
    .B1(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__a22oi_4 _05833_ (.A1(_02891_),
    .A2(_02913_),
    .B1(_05026_),
    .B2(_03572_),
    .Y(_05027_));
 sky130_fd_sc_hd__o211ai_4 _05834_ (.A1(_03352_),
    .A2(_05019_),
    .B1(_05027_),
    .C1(_05014_),
    .Y(_05028_));
 sky130_fd_sc_hd__a31oi_4 _05835_ (.A1(_05014_),
    .A2(_05027_),
    .A3(_05020_),
    .B1(_03913_),
    .Y(_05029_));
 sky130_fd_sc_hd__a31o_1 _05836_ (.A1(_05014_),
    .A2(_05027_),
    .A3(_05020_),
    .B1(_03913_),
    .X(_05030_));
 sky130_fd_sc_hd__a21oi_2 _05837_ (.A1(_05028_),
    .A2(_03902_),
    .B1(_05008_),
    .Y(_05031_));
 sky130_fd_sc_hd__a31o_1 _05838_ (.A1(net23),
    .A2(net107),
    .A3(net105),
    .B1(_05029_),
    .X(_05032_));
 sky130_fd_sc_hd__a22oi_2 _05839_ (.A1(net55),
    .A2(_02077_),
    .B1(_05028_),
    .B2(_04328_),
    .Y(_05033_));
 sky130_fd_sc_hd__a32o_1 _05840_ (.A1(net55),
    .A2(net112),
    .A3(net109),
    .B1(_05028_),
    .B2(_04328_),
    .X(_05034_));
 sky130_fd_sc_hd__a221o_1 _05841_ (.A1(_04949_),
    .A2(_04979_),
    .B1(_05031_),
    .B2(_05034_),
    .C1(_05007_),
    .X(_05035_));
 sky130_fd_sc_hd__o221a_1 _05842_ (.A1(_04623_),
    .A2(_04645_),
    .B1(_05031_),
    .B2(_05034_),
    .C1(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__a221oi_1 _05843_ (.A1(_04306_),
    .A2(_04339_),
    .B1(_04623_),
    .B2(_04645_),
    .C1(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nor2_1 _05844_ (.A(_04339_),
    .B(_04306_),
    .Y(_05038_));
 sky130_fd_sc_hd__a2bb2o_1 _05845_ (.A1_N(_05037_),
    .A2_N(_05038_),
    .B1(_03814_),
    .B2(_03891_),
    .X(_05039_));
 sky130_fd_sc_hd__o221a_4 _05846_ (.A1(_01043_),
    .A2(_02077_),
    .B1(_02209_),
    .B2(_02935_),
    .C1(_02231_),
    .X(_05040_));
 sky130_fd_sc_hd__a311o_2 _05847_ (.A1(net47),
    .A2(net107),
    .A3(net105),
    .B1(_02220_),
    .C1(_04819_),
    .X(_05041_));
 sky130_fd_sc_hd__o211a_1 _05848_ (.A1(_02462_),
    .A2(_04050_),
    .B1(_05017_),
    .C1(_02363_),
    .X(_05042_));
 sky130_fd_sc_hd__a31o_1 _05849_ (.A1(_02352_),
    .A2(_05010_),
    .A3(_05011_),
    .B1(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__nand2_1 _05850_ (.A(_05043_),
    .B(_02781_),
    .Y(_05044_));
 sky130_fd_sc_hd__a211o_1 _05851_ (.A1(_05023_),
    .A2(_05024_),
    .B1(_02330_),
    .C1(_02341_),
    .X(_05045_));
 sky130_fd_sc_hd__o221ai_1 _05852_ (.A1(_02330_),
    .A2(_02341_),
    .B1(_02462_),
    .B2(_04003_),
    .C1(_05015_),
    .Y(_05046_));
 sky130_fd_sc_hd__a311oi_1 _05853_ (.A1(_05045_),
    .A2(_05046_),
    .A3(_02770_),
    .B1(_02935_),
    .C1(_02209_),
    .Y(_05047_));
 sky130_fd_sc_hd__a21oi_1 _05854_ (.A1(_05047_),
    .A2(_05044_),
    .B1(_05040_),
    .Y(_05048_));
 sky130_fd_sc_hd__mux2_2 _05855_ (.A0(_05048_),
    .A1(net29),
    .S(_02088_),
    .X(_05049_));
 sky130_fd_sc_hd__inv_2 _05856_ (.A(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__mux2_4 _05857_ (.A0(_05048_),
    .A1(net61),
    .S(_02077_),
    .X(_05051_));
 sky130_fd_sc_hd__nor2_1 _05858_ (.A(_05051_),
    .B(_05050_),
    .Y(_05052_));
 sky130_fd_sc_hd__o221a_1 _05859_ (.A1(_03814_),
    .A2(_03891_),
    .B1(_05050_),
    .B2(_05051_),
    .C1(_05039_),
    .X(_05053_));
 sky130_fd_sc_hd__or4_1 _05860_ (.A(_02308_),
    .B(_02319_),
    .C(_04350_),
    .D(_04361_),
    .X(_05054_));
 sky130_fd_sc_hd__o21ai_1 _05861_ (.A1(_02352_),
    .A2(_04557_),
    .B1(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__o211ai_2 _05862_ (.A1(_04557_),
    .A2(_02352_),
    .B1(_02781_),
    .C1(_05054_),
    .Y(_05056_));
 sky130_fd_sc_hd__a211o_1 _05863_ (.A1(_04514_),
    .A2(_04524_),
    .B1(_02308_),
    .C1(_02319_),
    .X(_05057_));
 sky130_fd_sc_hd__o211ai_2 _05864_ (.A1(_02352_),
    .A2(_04404_),
    .B1(_02770_),
    .C1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__a31oi_4 _05865_ (.A1(_05056_),
    .A2(_05058_),
    .A3(_04819_),
    .B1(_05040_),
    .Y(_05059_));
 sky130_fd_sc_hd__and3_1 _05866_ (.A(_05059_),
    .B(net105),
    .C(net107),
    .X(_05060_));
 sky130_fd_sc_hd__and3_1 _05867_ (.A(net109),
    .B(net62),
    .C(net112),
    .X(_05061_));
 sky130_fd_sc_hd__a31o_1 _05868_ (.A1(_05059_),
    .A2(net105),
    .A3(net107),
    .B1(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__inv_2 _05869_ (.A(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__and3_1 _05870_ (.A(_05059_),
    .B(net109),
    .C(net112),
    .X(_05064_));
 sky130_fd_sc_hd__and3_1 _05871_ (.A(net105),
    .B(net30),
    .C(net107),
    .X(_05065_));
 sky130_fd_sc_hd__and3_1 _05872_ (.A(_01175_),
    .B(net107),
    .C(net105),
    .X(_05066_));
 sky130_fd_sc_hd__a21oi_1 _05873_ (.A1(net107),
    .A2(net105),
    .B1(_05059_),
    .Y(_05067_));
 sky130_fd_sc_hd__a31o_1 _05874_ (.A1(_01175_),
    .A2(net107),
    .A3(net105),
    .B1(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__a31o_1 _05875_ (.A1(_05059_),
    .A2(net109),
    .A3(net112),
    .B1(_05065_),
    .X(_05069_));
 sky130_fd_sc_hd__nand2_1 _05876_ (.A(_05050_),
    .B(_05051_),
    .Y(_05070_));
 sky130_fd_sc_hd__a221oi_1 _05877_ (.A1(_05050_),
    .A2(_05051_),
    .B1(_05062_),
    .B2(_05068_),
    .C1(_05053_),
    .Y(_05071_));
 sky130_fd_sc_hd__or3_1 _05878_ (.A(_02209_),
    .B(_02770_),
    .C(_02935_),
    .X(_05072_));
 sky130_fd_sc_hd__o221a_1 _05879_ (.A1(_02176_),
    .A2(_02187_),
    .B1(_02374_),
    .B2(_05012_),
    .C1(_02924_),
    .X(_05073_));
 sky130_fd_sc_hd__a32o_1 _05880_ (.A1(_02231_),
    .A2(_02242_),
    .A3(_04830_),
    .B1(_05073_),
    .B2(_02781_),
    .X(_05074_));
 sky130_fd_sc_hd__a31o_1 _05881_ (.A1(_02770_),
    .A2(_04819_),
    .A3(_05019_),
    .B1(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__and3_1 _05882_ (.A(_01131_),
    .B(net107),
    .C(net105),
    .X(_05076_));
 sky130_fd_sc_hd__a21oi_2 _05883_ (.A1(_05075_),
    .A2(_02077_),
    .B1(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__o21ai_1 _05884_ (.A1(_02033_),
    .A2(_02055_),
    .B1(net34),
    .Y(_05078_));
 sky130_fd_sc_hd__o21ai_2 _05885_ (.A1(_02077_),
    .A2(_05075_),
    .B1(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__inv_2 _05886_ (.A(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__o211a_1 _05887_ (.A1(_02077_),
    .A2(_01131_),
    .B1(_05078_),
    .C1(_05075_),
    .X(_05081_));
 sky130_fd_sc_hd__a311o_1 _05888_ (.A1(net112),
    .A2(net109),
    .A3(_05075_),
    .B1(_05076_),
    .C1(_05080_),
    .X(_05082_));
 sky130_fd_sc_hd__and2b_1 _05889_ (.A_N(_05081_),
    .B(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__nor2_1 _05890_ (.A(_05072_),
    .B(_04371_),
    .Y(_05084_));
 sky130_fd_sc_hd__and4_1 _05891_ (.A(_04568_),
    .B(_03572_),
    .C(_02924_),
    .D(_04535_),
    .X(_05085_));
 sky130_fd_sc_hd__or3_1 _05892_ (.A(_05040_),
    .B(_05084_),
    .C(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__and3_1 _05893_ (.A(_01120_),
    .B(net107),
    .C(net105),
    .X(_05087_));
 sky130_fd_sc_hd__a31o_1 _05894_ (.A1(net112),
    .A2(net109),
    .A3(_05086_),
    .B1(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__inv_2 _05895_ (.A(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__a21oi_1 _05896_ (.A1(net112),
    .A2(net109),
    .B1(_05086_),
    .Y(_05090_));
 sky130_fd_sc_hd__a31o_4 _05897_ (.A1(net35),
    .A2(net112),
    .A3(net109),
    .B1(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__inv_2 _05898_ (.A(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__a311o_1 _05899_ (.A1(net112),
    .A2(net109),
    .A3(_05086_),
    .B1(_05087_),
    .C1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__xnor2_2 _05900_ (.A(_05088_),
    .B(_05091_),
    .Y(_05094_));
 sky130_fd_sc_hd__a41oi_1 _05901_ (.A1(_04981_),
    .A2(_02924_),
    .A3(_04980_),
    .A4(_03341_),
    .B1(_05040_),
    .Y(_05095_));
 sky130_fd_sc_hd__o31a_1 _05902_ (.A1(_02781_),
    .A2(_04830_),
    .A3(_04987_),
    .B1(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__mux2_2 _05903_ (.A0(_05096_),
    .A1(net31),
    .S(_02088_),
    .X(_05097_));
 sky130_fd_sc_hd__inv_2 _05904_ (.A(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__mux2_4 _05905_ (.A0(_05096_),
    .A1(net63),
    .S(_02077_),
    .X(_05099_));
 sky130_fd_sc_hd__inv_2 _05906_ (.A(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _05907_ (.A(_05097_),
    .B(_05099_),
    .Y(_05101_));
 sky130_fd_sc_hd__or2_1 _05908_ (.A(_05097_),
    .B(_05099_),
    .X(_05102_));
 sky130_fd_sc_hd__and2_1 _05909_ (.A(_05101_),
    .B(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__o2111ai_1 _05910_ (.A1(_02363_),
    .A2(_02693_),
    .B1(_02781_),
    .C1(_04819_),
    .D1(_04841_),
    .Y(_05104_));
 sky130_fd_sc_hd__o311a_1 _05911_ (.A1(_02781_),
    .A2(_04677_),
    .A3(_04830_),
    .B1(_05041_),
    .C1(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__o21ai_1 _05912_ (.A1(_02033_),
    .A2(_02055_),
    .B1(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__o21ai_1 _05913_ (.A1(_01989_),
    .A2(net110),
    .B1(net32),
    .Y(_05107_));
 sky130_fd_sc_hd__a21oi_1 _05914_ (.A1(net112),
    .A2(net109),
    .B1(net32),
    .Y(_05108_));
 sky130_fd_sc_hd__a21oi_1 _05915_ (.A1(net107),
    .A2(net105),
    .B1(_05105_),
    .Y(_05109_));
 sky130_fd_sc_hd__or2_4 _05916_ (.A(_05108_),
    .B(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__mux2_4 _05917_ (.A0(_05105_),
    .A1(net64),
    .S(_02077_),
    .X(_05111_));
 sky130_fd_sc_hd__inv_2 _05918_ (.A(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__xnor2_1 _05919_ (.A(_05110_),
    .B(_05111_),
    .Y(_05113_));
 sky130_fd_sc_hd__or4_1 _05920_ (.A(_05094_),
    .B(_05103_),
    .C(_05113_),
    .D(_05083_),
    .X(_05114_));
 sky130_fd_sc_hd__nand2b_1 _05921_ (.A_N(_05052_),
    .B(_05070_),
    .Y(_05115_));
 sky130_fd_sc_hd__a211o_1 _05922_ (.A1(_05063_),
    .A2(_05069_),
    .B1(_05114_),
    .C1(_05071_),
    .X(_05116_));
 sky130_fd_sc_hd__o211a_1 _05923_ (.A1(_05111_),
    .A2(_05110_),
    .B1(_05099_),
    .C1(_05098_),
    .X(_05117_));
 sky130_fd_sc_hd__a21oi_1 _05924_ (.A1(_05110_),
    .A2(_05111_),
    .B1(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__a211o_1 _05925_ (.A1(_05089_),
    .A2(_05092_),
    .B1(_05077_),
    .C1(_05080_),
    .X(_05119_));
 sky130_fd_sc_hd__o32a_1 _05926_ (.A1(_05094_),
    .A2(_05118_),
    .A3(_05083_),
    .B1(_05089_),
    .B2(_05092_),
    .X(_05120_));
 sky130_fd_sc_hd__and3_1 _05927_ (.A(_05116_),
    .B(_05119_),
    .C(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__o2bb2a_1 _05928_ (.A1_N(_03965_),
    .A2_N(_03341_),
    .B1(_03583_),
    .B2(_04099_),
    .X(_05122_));
 sky130_fd_sc_hd__o21a_1 _05929_ (.A1(_02935_),
    .A2(_05122_),
    .B1(_05041_),
    .X(_05123_));
 sky130_fd_sc_hd__mux2_4 _05930_ (.A0(_05123_),
    .A1(net4),
    .S(_02088_),
    .X(_05124_));
 sky130_fd_sc_hd__mux2_4 _05931_ (.A0(_05123_),
    .A1(net36),
    .S(_02077_),
    .X(_05125_));
 sky130_fd_sc_hd__inv_2 _05932_ (.A(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__nor2_1 _05933_ (.A(_05124_),
    .B(_05125_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _05934_ (.A(_05124_),
    .B(_05125_),
    .Y(_05128_));
 sky130_fd_sc_hd__and2b_1 _05935_ (.A_N(_05127_),
    .B(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__a31o_1 _05936_ (.A1(_02198_),
    .A2(_02770_),
    .A3(_02924_),
    .B1(_02264_),
    .X(_05130_));
 sky130_fd_sc_hd__a31o_1 _05937_ (.A1(_02231_),
    .A2(_02242_),
    .A3(_04830_),
    .B1(_02792_),
    .X(_05131_));
 sky130_fd_sc_hd__o311a_1 _05938_ (.A1(_02781_),
    .A2(_04830_),
    .A3(_05043_),
    .B1(_05041_),
    .C1(_02803_),
    .X(_05132_));
 sky130_fd_sc_hd__mux2_4 _05939_ (.A0(_05132_),
    .A1(net38),
    .S(_02077_),
    .X(_05133_));
 sky130_fd_sc_hd__inv_2 _05940_ (.A(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__mux2_2 _05941_ (.A0(_05132_),
    .A1(net6),
    .S(_02088_),
    .X(_05135_));
 sky130_fd_sc_hd__nor2_1 _05942_ (.A(_05133_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__and2_1 _05943_ (.A(_05133_),
    .B(_05135_),
    .X(_05137_));
 sky130_fd_sc_hd__nor2_1 _05944_ (.A(_05136_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__a311oi_1 _05945_ (.A1(_02770_),
    .A2(_04819_),
    .A3(_05055_),
    .B1(_05040_),
    .C1(_02792_),
    .Y(_05139_));
 sky130_fd_sc_hd__mux2_4 _05946_ (.A0(_05139_),
    .A1(net39),
    .S(_02077_),
    .X(_05140_));
 sky130_fd_sc_hd__or3_1 _05947_ (.A(_01989_),
    .B(net110),
    .C(_05139_),
    .X(_05141_));
 sky130_fd_sc_hd__o21ai_4 _05948_ (.A1(net7),
    .A2(_02077_),
    .B1(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__o31a_2 _05949_ (.A1(net7),
    .A2(_02033_),
    .A3(_02055_),
    .B1(_05141_),
    .X(_05143_));
 sky130_fd_sc_hd__xnor2_1 _05950_ (.A(_05140_),
    .B(_05142_),
    .Y(_05144_));
 sky130_fd_sc_hd__or2_1 _05951_ (.A(_05138_),
    .B(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__o2111ai_1 _05952_ (.A1(_02176_),
    .A2(_02187_),
    .B1(_03330_),
    .C1(_02770_),
    .D1(_03121_),
    .Y(_05146_));
 sky130_fd_sc_hd__o221a_2 _05953_ (.A1(_05072_),
    .A2(_02704_),
    .B1(_02935_),
    .B2(_05146_),
    .C1(_05041_),
    .X(_05147_));
 sky130_fd_sc_hd__mux2_4 _05954_ (.A0(_05147_),
    .A1(net37),
    .S(_02077_),
    .X(_05148_));
 sky130_fd_sc_hd__inv_2 _05955_ (.A(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__o21ai_4 _05956_ (.A1(_02033_),
    .A2(_02055_),
    .B1(_05147_),
    .Y(_05150_));
 sky130_fd_sc_hd__or3_1 _05957_ (.A(_01098_),
    .B(_02033_),
    .C(_02055_),
    .X(_05151_));
 sky130_fd_sc_hd__a21oi_1 _05958_ (.A1(_02044_),
    .A2(net105),
    .B1(_05147_),
    .Y(_05152_));
 sky130_fd_sc_hd__and3_1 _05959_ (.A(_01098_),
    .B(_02044_),
    .C(net105),
    .X(_05153_));
 sky130_fd_sc_hd__a31o_1 _05960_ (.A1(_01098_),
    .A2(_02044_),
    .A3(net105),
    .B1(_05152_),
    .X(_05154_));
 sky130_fd_sc_hd__o21ai_4 _05961_ (.A1(_01098_),
    .A2(_02077_),
    .B1(_05150_),
    .Y(_05155_));
 sky130_fd_sc_hd__xor2_1 _05962_ (.A(_05148_),
    .B(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__or4_1 _05963_ (.A(_05145_),
    .B(_05156_),
    .C(_05121_),
    .D(_05129_),
    .X(_05157_));
 sky130_fd_sc_hd__o22a_1 _05964_ (.A1(_05149_),
    .A2(_05155_),
    .B1(_05124_),
    .B2(_05126_),
    .X(_05158_));
 sky130_fd_sc_hd__a2111oi_1 _05965_ (.A1(_05149_),
    .A2(_05155_),
    .B1(_05158_),
    .C1(_05138_),
    .D1(_05144_),
    .Y(_05159_));
 sky130_fd_sc_hd__o21ba_1 _05966_ (.A1(_05140_),
    .A2(_05142_),
    .B1_N(_05135_),
    .X(_05160_));
 sky130_fd_sc_hd__a221oi_1 _05967_ (.A1(_05140_),
    .A2(_05142_),
    .B1(_05160_),
    .B2(_05133_),
    .C1(_05159_),
    .Y(_05161_));
 sky130_fd_sc_hd__o221a_1 _05968_ (.A1(_02264_),
    .A2(_02770_),
    .B1(_04830_),
    .B2(_05013_),
    .C1(_05041_),
    .X(_05162_));
 sky130_fd_sc_hd__mux2_4 _05969_ (.A0(_05162_),
    .A1(net42),
    .S(_02077_),
    .X(_05163_));
 sky130_fd_sc_hd__mux2_2 _05970_ (.A0(_05162_),
    .A1(net10),
    .S(_02088_),
    .X(_05164_));
 sky130_fd_sc_hd__inv_2 _05971_ (.A(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__or2_1 _05972_ (.A(_05163_),
    .B(_05164_),
    .X(_05166_));
 sky130_fd_sc_hd__nand2_1 _05973_ (.A(_05163_),
    .B(_05164_),
    .Y(_05167_));
 sky130_fd_sc_hd__inv_2 _05974_ (.A(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand2_1 _05975_ (.A(_05166_),
    .B(_05167_),
    .Y(_05169_));
 sky130_fd_sc_hd__o31a_1 _05976_ (.A1(_02781_),
    .A2(_04830_),
    .A3(_04371_),
    .B1(_05130_),
    .X(_05170_));
 sky130_fd_sc_hd__mux2_8 _05977_ (.A0(_05170_),
    .A1(net43),
    .S(_02077_),
    .X(_05171_));
 sky130_fd_sc_hd__or3_2 _05978_ (.A(_01989_),
    .B(net110),
    .C(_05170_),
    .X(_05172_));
 sky130_fd_sc_hd__o21ai_4 _05979_ (.A1(net11),
    .A2(_02077_),
    .B1(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__o21a_2 _05980_ (.A1(net11),
    .A2(_02077_),
    .B1(_05172_),
    .X(_05174_));
 sky130_fd_sc_hd__xor2_2 _05981_ (.A(_05171_),
    .B(_05173_),
    .X(_05175_));
 sky130_fd_sc_hd__o311a_2 _05982_ (.A1(_02209_),
    .A2(_02935_),
    .A3(_04862_),
    .B1(_05130_),
    .C1(_02077_),
    .X(_05176_));
 sky130_fd_sc_hd__and3_1 _05983_ (.A(net105),
    .B(net9),
    .C(_02044_),
    .X(_05177_));
 sky130_fd_sc_hd__a21oi_4 _05984_ (.A1(net9),
    .A2(_02088_),
    .B1(_05176_),
    .Y(_05178_));
 sky130_fd_sc_hd__a31o_1 _05985_ (.A1(net9),
    .A2(_02044_),
    .A3(net105),
    .B1(_05176_),
    .X(_05179_));
 sky130_fd_sc_hd__o221a_1 _05986_ (.A1(_01989_),
    .A2(net110),
    .B1(_04830_),
    .B2(_04862_),
    .C1(_05130_),
    .X(_05180_));
 sky130_fd_sc_hd__a21oi_2 _05987_ (.A1(net41),
    .A2(_02077_),
    .B1(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__a31o_4 _05988_ (.A1(net41),
    .A2(net112),
    .A3(net109),
    .B1(_05180_),
    .X(_05182_));
 sky130_fd_sc_hd__xnor2_1 _05989_ (.A(_05178_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__o311a_1 _05990_ (.A1(_02209_),
    .A2(_02935_),
    .A3(_04982_),
    .B1(_05041_),
    .C1(_02803_),
    .X(_05184_));
 sky130_fd_sc_hd__mux2_4 _05991_ (.A0(_05184_),
    .A1(net8),
    .S(_02088_),
    .X(_05185_));
 sky130_fd_sc_hd__inv_2 _05992_ (.A(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__mux2_4 _05993_ (.A0(_05184_),
    .A1(net40),
    .S(_02077_),
    .X(_05187_));
 sky130_fd_sc_hd__nand2_1 _05994_ (.A(_05185_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__or2_1 _05995_ (.A(_05185_),
    .B(_05187_),
    .X(_05189_));
 sky130_fd_sc_hd__nand2_1 _05996_ (.A(_05188_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand3_1 _05997_ (.A(_05175_),
    .B(_05190_),
    .C(_05169_),
    .Y(_05191_));
 sky130_fd_sc_hd__a211o_1 _05998_ (.A1(_05157_),
    .A2(_05161_),
    .B1(_05183_),
    .C1(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__a22o_1 _05999_ (.A1(_05178_),
    .A2(_05182_),
    .B1(_05186_),
    .B2(_05187_),
    .X(_05193_));
 sky130_fd_sc_hd__o211a_1 _06000_ (.A1(_05178_),
    .A2(_05182_),
    .B1(_05193_),
    .C1(_05175_),
    .X(_05194_));
 sky130_fd_sc_hd__o21a_1 _06001_ (.A1(_05171_),
    .A2(_05173_),
    .B1(_05165_),
    .X(_05195_));
 sky130_fd_sc_hd__a22o_1 _06002_ (.A1(_05171_),
    .A2(_05173_),
    .B1(_05195_),
    .B2(_05163_),
    .X(_05196_));
 sky130_fd_sc_hd__a21oi_2 _06003_ (.A1(_05194_),
    .A2(_05169_),
    .B1(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__and4b_1 _06004_ (.A_N(_02704_),
    .B(_02770_),
    .C(_02924_),
    .D(_02198_),
    .X(_05198_));
 sky130_fd_sc_hd__o32a_1 _06005_ (.A1(_02792_),
    .A2(_05040_),
    .A3(_05198_),
    .B1(net110),
    .B2(_01989_),
    .X(_05199_));
 sky130_fd_sc_hd__a21oi_1 _06006_ (.A1(net107),
    .A2(net105),
    .B1(net46),
    .Y(_05200_));
 sky130_fd_sc_hd__o21ai_2 _06007_ (.A1(_02033_),
    .A2(_02055_),
    .B1(net46),
    .Y(_05201_));
 sky130_fd_sc_hd__a211o_2 _06008_ (.A1(_02814_),
    .A2(_04819_),
    .B1(_05040_),
    .C1(_02077_),
    .X(_05202_));
 sky130_fd_sc_hd__nand2_2 _06009_ (.A(_05201_),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__and3_2 _06010_ (.A(net105),
    .B(net14),
    .C(net107),
    .X(_05204_));
 sky130_fd_sc_hd__a21oi_4 _06011_ (.A1(net15),
    .A2(_02077_),
    .B1(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__xnor2_4 _06012_ (.A(_05203_),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__a31oi_4 _06013_ (.A1(_03965_),
    .A2(_04819_),
    .A3(_02770_),
    .B1(_05131_),
    .Y(_05207_));
 sky130_fd_sc_hd__and3_2 _06014_ (.A(net105),
    .B(net13),
    .C(net107),
    .X(_05208_));
 sky130_fd_sc_hd__and3_1 _06015_ (.A(_05207_),
    .B(net109),
    .C(net111),
    .X(_05209_));
 sky130_fd_sc_hd__a31o_1 _06016_ (.A1(_05207_),
    .A2(net109),
    .A3(net112),
    .B1(_05208_),
    .X(_05210_));
 sky130_fd_sc_hd__a21oi_4 _06017_ (.A1(_02077_),
    .A2(_05207_),
    .B1(_05208_),
    .Y(_05211_));
 sky130_fd_sc_hd__a21oi_1 _06018_ (.A1(net112),
    .A2(net109),
    .B1(_05207_),
    .Y(_05212_));
 sky130_fd_sc_hd__and3_1 _06019_ (.A(_01054_),
    .B(net112),
    .C(net109),
    .X(_05213_));
 sky130_fd_sc_hd__and3_1 _06020_ (.A(net108),
    .B(net45),
    .C(net111),
    .X(_05214_));
 sky130_fd_sc_hd__or3_1 _06021_ (.A(_01054_),
    .B(_01989_),
    .C(_02011_),
    .X(_05215_));
 sky130_fd_sc_hd__o21a_1 _06022_ (.A1(_01989_),
    .A2(net110),
    .B1(_05207_),
    .X(_05216_));
 sky130_fd_sc_hd__a311o_2 _06023_ (.A1(_03965_),
    .A2(_03572_),
    .A3(_02924_),
    .B1(_02077_),
    .C1(_05131_),
    .X(_05217_));
 sky130_fd_sc_hd__a31o_1 _06024_ (.A1(net45),
    .A2(net111),
    .A3(net108),
    .B1(_05216_),
    .X(_05218_));
 sky130_fd_sc_hd__a31o_2 _06025_ (.A1(_01054_),
    .A2(net112),
    .A3(net109),
    .B1(_05212_),
    .X(_05219_));
 sky130_fd_sc_hd__o311a_1 _06026_ (.A1(_01054_),
    .A2(_01989_),
    .A3(_02011_),
    .B1(_05211_),
    .C1(_05217_),
    .X(_05220_));
 sky130_fd_sc_hd__a21oi_2 _06027_ (.A1(_05215_),
    .A2(_05217_),
    .B1(_05211_),
    .Y(_05221_));
 sky130_fd_sc_hd__nor2_1 _06028_ (.A(_05220_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__or2_1 _06029_ (.A(_05220_),
    .B(_05221_),
    .X(_05223_));
 sky130_fd_sc_hd__a211oi_4 _06030_ (.A1(_05192_),
    .A2(_05197_),
    .B1(_05206_),
    .C1(_05222_),
    .Y(_05224_));
 sky130_fd_sc_hd__nor2_1 _06031_ (.A(net15),
    .B(net47),
    .Y(_05225_));
 sky130_fd_sc_hd__nor2_2 _06032_ (.A(_01032_),
    .B(_01043_),
    .Y(_05226_));
 sky130_fd_sc_hd__nor2_2 _06033_ (.A(_05225_),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__o211a_1 _06034_ (.A1(_05203_),
    .A2(_05205_),
    .B1(_05211_),
    .C1(_05218_),
    .X(_05228_));
 sky130_fd_sc_hd__a2bb2o_1 _06035_ (.A1_N(_05225_),
    .A2_N(_05226_),
    .B1(_05205_),
    .B2(_05203_),
    .X(_05229_));
 sky130_fd_sc_hd__o32a_4 _06036_ (.A1(_05229_),
    .A2(_05228_),
    .A3(_05224_),
    .B1(net15),
    .B2(_01043_),
    .X(_05230_));
 sky130_fd_sc_hd__o32ai_4 _06037_ (.A1(_05229_),
    .A2(_05228_),
    .A3(_05224_),
    .B1(net15),
    .B2(_01043_),
    .Y(_05231_));
 sky130_fd_sc_hd__xnor2_4 _06038_ (.A(net25),
    .B(net57),
    .Y(_05232_));
 sky130_fd_sc_hd__xor2_4 _06039_ (.A(net25),
    .B(net57),
    .X(_05233_));
 sky130_fd_sc_hd__nand2_8 _06040_ (.A(_05230_),
    .B(net115),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_4 _06041_ (.A(_05230_),
    .B(_05232_),
    .Y(_05234_));
 sky130_fd_sc_hd__inv_4 _06042_ (.A(_05234_),
    .Y(_00001_));
 sky130_fd_sc_hd__nor2_1 _06043_ (.A(_01032_),
    .B(_01065_),
    .Y(_05235_));
 sky130_fd_sc_hd__a21o_1 _06044_ (.A1(net15),
    .A2(net43),
    .B1(_01054_),
    .X(_05236_));
 sky130_fd_sc_hd__and3_1 _06045_ (.A(net46),
    .B(net15),
    .C(net47),
    .X(_05237_));
 sky130_fd_sc_hd__and3_2 _06046_ (.A(net46),
    .B(net14),
    .C(_05226_),
    .X(_05238_));
 sky130_fd_sc_hd__a22oi_2 _06047_ (.A1(net46),
    .A2(net15),
    .B1(net47),
    .B2(net14),
    .Y(_05239_));
 sky130_fd_sc_hd__nor3b_2 _06048_ (.A(_05238_),
    .B(_05239_),
    .C_N(net13),
    .Y(_05240_));
 sky130_fd_sc_hd__o21ba_1 _06049_ (.A1(_05238_),
    .A2(_05239_),
    .B1_N(net13),
    .X(_05241_));
 sky130_fd_sc_hd__nor2_1 _06050_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__xor2_2 _06051_ (.A(_05236_),
    .B(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__and4_1 _06052_ (.A(net46),
    .B(net47),
    .C(net14),
    .D(net13),
    .X(_05244_));
 sky130_fd_sc_hd__a22oi_1 _06053_ (.A1(net46),
    .A2(net14),
    .B1(net13),
    .B2(net47),
    .Y(_05245_));
 sky130_fd_sc_hd__nor2_1 _06054_ (.A(_05244_),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21oi_1 _06055_ (.A1(net11),
    .A2(_05246_),
    .B1(_05244_),
    .Y(_05247_));
 sky130_fd_sc_hd__and3_1 _06056_ (.A(net15),
    .B(net45),
    .C(net43),
    .X(_05248_));
 sky130_fd_sc_hd__a21oi_1 _06057_ (.A1(net15),
    .A2(net45),
    .B1(net43),
    .Y(_05249_));
 sky130_fd_sc_hd__or3b_2 _06058_ (.A(_01032_),
    .B(_01065_),
    .C_N(net42),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_1 _06059_ (.A1(net15),
    .A2(net43),
    .B1(net42),
    .X(_05251_));
 sky130_fd_sc_hd__nand4_2 _06060_ (.A(_05250_),
    .B(_05251_),
    .C(net14),
    .D(net45),
    .Y(_05252_));
 sky130_fd_sc_hd__a221oi_1 _06061_ (.A1(net45),
    .A2(_05235_),
    .B1(_05250_),
    .B2(_05252_),
    .C1(_05249_),
    .Y(_05253_));
 sky130_fd_sc_hd__a221o_1 _06062_ (.A1(net45),
    .A2(_05235_),
    .B1(_05250_),
    .B2(_05252_),
    .C1(_05249_),
    .X(_05254_));
 sky130_fd_sc_hd__xnor2_1 _06063_ (.A(net11),
    .B(_05246_),
    .Y(_05255_));
 sky130_fd_sc_hd__o211a_1 _06064_ (.A1(_05248_),
    .A2(_05249_),
    .B1(_05250_),
    .C1(_05252_),
    .X(_05256_));
 sky130_fd_sc_hd__or2_1 _06065_ (.A(_05253_),
    .B(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__o21ai_1 _06066_ (.A1(_05255_),
    .A2(_05257_),
    .B1(_05254_),
    .Y(_05258_));
 sky130_fd_sc_hd__xnor2_1 _06067_ (.A(_05255_),
    .B(_05257_),
    .Y(_05259_));
 sky130_fd_sc_hd__and2_1 _06068_ (.A(net15),
    .B(net40),
    .X(_05260_));
 sky130_fd_sc_hd__and3_1 _06069_ (.A(net15),
    .B(net41),
    .C(net40),
    .X(_05261_));
 sky130_fd_sc_hd__nand2_1 _06070_ (.A(net41),
    .B(_05260_),
    .Y(_05262_));
 sky130_fd_sc_hd__and4_1 _06071_ (.A(net46),
    .B(net47),
    .C(net13),
    .D(net11),
    .X(_05263_));
 sky130_fd_sc_hd__a22oi_1 _06072_ (.A1(net46),
    .A2(net13),
    .B1(net11),
    .B2(net47),
    .Y(_05264_));
 sky130_fd_sc_hd__nor2_1 _06073_ (.A(_05263_),
    .B(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__xnor2_1 _06074_ (.A(net10),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__and3_1 _06075_ (.A(net14),
    .B(net42),
    .C(_05235_),
    .X(_05267_));
 sky130_fd_sc_hd__a22oi_1 _06076_ (.A1(net14),
    .A2(net43),
    .B1(net42),
    .B2(net15),
    .Y(_05268_));
 sky130_fd_sc_hd__and4bb_1 _06077_ (.A_N(_05267_),
    .B_N(_05268_),
    .C(net45),
    .D(net13),
    .X(_05269_));
 sky130_fd_sc_hd__a22o_1 _06078_ (.A1(net14),
    .A2(net45),
    .B1(_05250_),
    .B2(_05251_),
    .X(_05270_));
 sky130_fd_sc_hd__a211o_1 _06079_ (.A1(_05252_),
    .A2(_05270_),
    .B1(_05269_),
    .C1(_05267_),
    .X(_05271_));
 sky130_fd_sc_hd__o211ai_2 _06080_ (.A1(_05267_),
    .A2(_05269_),
    .B1(_05270_),
    .C1(_05252_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand2_1 _06081_ (.A(_05271_),
    .B(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__or2_1 _06082_ (.A(_05266_),
    .B(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__nand2_1 _06083_ (.A(_05266_),
    .B(_05273_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_1 _06084_ (.A(_05274_),
    .B(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__or2_1 _06085_ (.A(_05262_),
    .B(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__nor2_1 _06086_ (.A(_05259_),
    .B(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__or4b_1 _06087_ (.A(_05259_),
    .B(_05262_),
    .C(_05276_),
    .D_N(_05258_),
    .X(_05279_));
 sky130_fd_sc_hd__or2_1 _06088_ (.A(_05258_),
    .B(_05278_),
    .X(_05280_));
 sky130_fd_sc_hd__nand2_1 _06089_ (.A(_05279_),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__xnor2_1 _06090_ (.A(_05247_),
    .B(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__o21a_1 _06091_ (.A1(_05235_),
    .A2(_05242_),
    .B1(net45),
    .X(_05283_));
 sky130_fd_sc_hd__o21ai_4 _06092_ (.A1(_05238_),
    .A2(_05240_),
    .B1(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__or3_1 _06093_ (.A(_05238_),
    .B(_05240_),
    .C(_05283_),
    .X(_05285_));
 sky130_fd_sc_hd__nand2_1 _06094_ (.A(_05284_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__a21oi_1 _06095_ (.A1(net15),
    .A2(net47),
    .B1(net46),
    .Y(_05287_));
 sky130_fd_sc_hd__or3b_2 _06096_ (.A(_05237_),
    .B(_05287_),
    .C_N(net14),
    .X(_05288_));
 sky130_fd_sc_hd__o21bai_1 _06097_ (.A1(_05237_),
    .A2(_05287_),
    .B1_N(net14),
    .Y(_05289_));
 sky130_fd_sc_hd__nand2_1 _06098_ (.A(_05288_),
    .B(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__or2_1 _06099_ (.A(_05286_),
    .B(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__a22o_1 _06100_ (.A1(_05284_),
    .A2(_05285_),
    .B1(_05288_),
    .B2(_05289_),
    .X(_05292_));
 sky130_fd_sc_hd__nand2_1 _06101_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__nor3_1 _06102_ (.A(_05243_),
    .B(_05282_),
    .C(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__o21ai_1 _06103_ (.A1(_05247_),
    .A2(_05281_),
    .B1(_05279_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_1 _06104_ (.A1(_05243_),
    .A2(_05282_),
    .B1(_05293_),
    .Y(_05296_));
 sky130_fd_sc_hd__nand2b_1 _06105_ (.A_N(_05294_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__a21o_1 _06106_ (.A1(_05295_),
    .A2(_05296_),
    .B1(_05294_),
    .X(_05298_));
 sky130_fd_sc_hd__o2bb2a_1 _06107_ (.A1_N(net46),
    .A2_N(net15),
    .B1(_05225_),
    .B2(_05226_),
    .X(_05299_));
 sky130_fd_sc_hd__a32oi_4 _06108_ (.A1(net46),
    .A2(net14),
    .A3(_05227_),
    .B1(_05288_),
    .B2(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__o21ai_1 _06109_ (.A1(_05286_),
    .A2(_05290_),
    .B1(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__or3_1 _06110_ (.A(_05300_),
    .B(_05290_),
    .C(_05286_),
    .X(_05302_));
 sky130_fd_sc_hd__a21bo_1 _06111_ (.A1(_05301_),
    .A2(_05302_),
    .B1_N(_05284_),
    .X(_05303_));
 sky130_fd_sc_hd__o21ai_1 _06112_ (.A1(_05284_),
    .A2(_05300_),
    .B1(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__and2_2 _06113_ (.A(_05298_),
    .B(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__a21oi_1 _06114_ (.A1(net10),
    .A2(_05265_),
    .B1(_05263_),
    .Y(_05306_));
 sky130_fd_sc_hd__a21bo_1 _06115_ (.A1(net15),
    .A2(net40),
    .B1_N(net41),
    .X(_05307_));
 sky130_fd_sc_hd__and3_1 _06116_ (.A(net15),
    .B(net40),
    .C(net39),
    .X(_05308_));
 sky130_fd_sc_hd__nand2_1 _06117_ (.A(net39),
    .B(_05260_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21oi_1 _06118_ (.A1(net15),
    .A2(net40),
    .B1(net39),
    .Y(_05310_));
 sky130_fd_sc_hd__or4bb_2 _06119_ (.A(_05308_),
    .B(_05310_),
    .C_N(net14),
    .D_N(net41),
    .X(_05311_));
 sky130_fd_sc_hd__a21oi_1 _06120_ (.A1(net15),
    .A2(net41),
    .B1(net40),
    .Y(_05312_));
 sky130_fd_sc_hd__a221o_1 _06121_ (.A1(net41),
    .A2(_05260_),
    .B1(_05309_),
    .B2(_05311_),
    .C1(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__xor2_1 _06122_ (.A(_05307_),
    .B(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__and4_1 _06123_ (.A(net46),
    .B(net47),
    .C(net11),
    .D(net10),
    .X(_05315_));
 sky130_fd_sc_hd__a22oi_1 _06124_ (.A1(net46),
    .A2(net11),
    .B1(net10),
    .B2(net47),
    .Y(_05316_));
 sky130_fd_sc_hd__o21a_1 _06125_ (.A1(_05315_),
    .A2(_05316_),
    .B1(_01076_),
    .X(_05317_));
 sky130_fd_sc_hd__nor3_1 _06126_ (.A(_05316_),
    .B(_01076_),
    .C(_05315_),
    .Y(_05318_));
 sky130_fd_sc_hd__and4_1 _06127_ (.A(net14),
    .B(net13),
    .C(net43),
    .D(net42),
    .X(_05319_));
 sky130_fd_sc_hd__a22oi_1 _06128_ (.A1(net13),
    .A2(net43),
    .B1(net42),
    .B2(net14),
    .Y(_05320_));
 sky130_fd_sc_hd__and4bb_1 _06129_ (.A_N(_05319_),
    .B_N(_05320_),
    .C(net45),
    .D(net11),
    .X(_05321_));
 sky130_fd_sc_hd__a41o_1 _06130_ (.A1(net14),
    .A2(net13),
    .A3(net43),
    .A4(net42),
    .B1(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__o2bb2a_1 _06131_ (.A1_N(net45),
    .A2_N(net13),
    .B1(_05267_),
    .B2(_05268_),
    .X(_05323_));
 sky130_fd_sc_hd__nor2_1 _06132_ (.A(_05269_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__xnor2_1 _06133_ (.A(_05322_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__nor3_1 _06134_ (.A(_05317_),
    .B(_05318_),
    .C(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__o21a_1 _06135_ (.A1(_05317_),
    .A2(_05318_),
    .B1(_05325_),
    .X(_05327_));
 sky130_fd_sc_hd__nor2_1 _06136_ (.A(_05326_),
    .B(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__nand2_1 _06137_ (.A(_05314_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__o21ai_1 _06138_ (.A1(_05307_),
    .A2(_05313_),
    .B1(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _06139_ (.A(_05262_),
    .B(_05276_),
    .Y(_05331_));
 sky130_fd_sc_hd__and2_1 _06140_ (.A(_05277_),
    .B(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__nand2_1 _06141_ (.A(_05330_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__a21oi_2 _06142_ (.A1(_05272_),
    .A2(_05274_),
    .B1(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__and3_1 _06143_ (.A(_05272_),
    .B(_05274_),
    .C(_05333_),
    .X(_05335_));
 sky130_fd_sc_hd__nor3_1 _06144_ (.A(_05306_),
    .B(_05334_),
    .C(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__o21a_1 _06145_ (.A1(_05334_),
    .A2(_05335_),
    .B1(_05306_),
    .X(_05337_));
 sky130_fd_sc_hd__or2_1 _06146_ (.A(_05336_),
    .B(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__o21a_1 _06147_ (.A1(_05262_),
    .A2(_05276_),
    .B1(_05259_),
    .X(_05339_));
 sky130_fd_sc_hd__or2_1 _06148_ (.A(_05278_),
    .B(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__xor2_1 _06149_ (.A(_05243_),
    .B(_05282_),
    .X(_05341_));
 sky130_fd_sc_hd__or3b_2 _06150_ (.A(_05338_),
    .B(_05340_),
    .C_N(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__o21bai_1 _06151_ (.A1(_05338_),
    .A2(_05340_),
    .B1_N(_05341_),
    .Y(_05343_));
 sky130_fd_sc_hd__o211ai_2 _06152_ (.A1(_05334_),
    .A2(_05336_),
    .B1(_05342_),
    .C1(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__xor2_1 _06153_ (.A(_05295_),
    .B(_05297_),
    .X(_05345_));
 sky130_fd_sc_hd__a21oi_1 _06154_ (.A1(_05342_),
    .A2(_05344_),
    .B1(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__and3_1 _06155_ (.A(_05342_),
    .B(_05344_),
    .C(_05345_),
    .X(_05347_));
 sky130_fd_sc_hd__or2_1 _06156_ (.A(_05346_),
    .B(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__inv_2 _06157_ (.A(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__a41o_1 _06158_ (.A1(net46),
    .A2(net47),
    .A3(net11),
    .A4(net10),
    .B1(_05318_),
    .X(_05350_));
 sky130_fd_sc_hd__a21o_1 _06159_ (.A1(_05322_),
    .A2(_05324_),
    .B1(_05326_),
    .X(_05351_));
 sky130_fd_sc_hd__xor2_1 _06160_ (.A(_05314_),
    .B(_05328_),
    .X(_05352_));
 sky130_fd_sc_hd__and3_1 _06161_ (.A(net14),
    .B(net39),
    .C(_05260_),
    .X(_05353_));
 sky130_fd_sc_hd__a22oi_1 _06162_ (.A1(net14),
    .A2(net40),
    .B1(net39),
    .B2(net15),
    .Y(_05354_));
 sky130_fd_sc_hd__and4bb_1 _06163_ (.A_N(_05353_),
    .B_N(_05354_),
    .C(net13),
    .D(net41),
    .X(_05355_));
 sky130_fd_sc_hd__a2bb2o_1 _06164_ (.A1_N(_05308_),
    .A2_N(_05310_),
    .B1(net14),
    .B2(net41),
    .X(_05356_));
 sky130_fd_sc_hd__o211ai_2 _06165_ (.A1(_05353_),
    .A2(_05355_),
    .B1(_05356_),
    .C1(_05311_),
    .Y(_05357_));
 sky130_fd_sc_hd__and4_1 _06166_ (.A(net46),
    .B(net47),
    .C(net10),
    .D(net9),
    .X(_05358_));
 sky130_fd_sc_hd__o2bb2a_1 _06167_ (.A1_N(net46),
    .A2_N(net10),
    .B1(_01076_),
    .B2(_01043_),
    .X(_05359_));
 sky130_fd_sc_hd__nor2_1 _06168_ (.A(_05358_),
    .B(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__xnor2_1 _06169_ (.A(net8),
    .B(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__and4_1 _06170_ (.A(net13),
    .B(net43),
    .C(net11),
    .D(net42),
    .X(_05362_));
 sky130_fd_sc_hd__a22oi_1 _06171_ (.A1(net43),
    .A2(net11),
    .B1(net42),
    .B2(net13),
    .Y(_05363_));
 sky130_fd_sc_hd__and4bb_1 _06172_ (.A_N(_05362_),
    .B_N(_05363_),
    .C(net45),
    .D(net10),
    .X(_05364_));
 sky130_fd_sc_hd__a41o_1 _06173_ (.A1(net13),
    .A2(net43),
    .A3(net11),
    .A4(net42),
    .B1(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__o2bb2a_1 _06174_ (.A1_N(net45),
    .A2_N(net11),
    .B1(_05319_),
    .B2(_05320_),
    .X(_05366_));
 sky130_fd_sc_hd__nor2_1 _06175_ (.A(_05321_),
    .B(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__xor2_1 _06176_ (.A(_05365_),
    .B(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__and2b_1 _06177_ (.A_N(_05361_),
    .B(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__xnor2_1 _06178_ (.A(_05361_),
    .B(_05368_),
    .Y(_05370_));
 sky130_fd_sc_hd__o211ai_1 _06179_ (.A1(_05261_),
    .A2(_05312_),
    .B1(_05311_),
    .C1(_05309_),
    .Y(_05371_));
 sky130_fd_sc_hd__and3_1 _06180_ (.A(_05313_),
    .B(_05357_),
    .C(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__a21bo_1 _06181_ (.A1(_05370_),
    .A2(_05372_),
    .B1_N(_05357_),
    .X(_05373_));
 sky130_fd_sc_hd__and2_1 _06182_ (.A(_05352_),
    .B(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__a221o_1 _06183_ (.A1(_05322_),
    .A2(_05324_),
    .B1(_05352_),
    .B2(_05373_),
    .C1(_05326_),
    .X(_05375_));
 sky130_fd_sc_hd__nand2_1 _06184_ (.A(_05374_),
    .B(_05351_),
    .Y(_05376_));
 sky130_fd_sc_hd__and3_1 _06185_ (.A(_05350_),
    .B(_05375_),
    .C(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__a21oi_1 _06186_ (.A1(_05375_),
    .A2(_05376_),
    .B1(_05350_),
    .Y(_05378_));
 sky130_fd_sc_hd__or2_1 _06187_ (.A(_05377_),
    .B(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__or2_1 _06188_ (.A(_05332_),
    .B(_05330_),
    .X(_05380_));
 sky130_fd_sc_hd__nand2_1 _06189_ (.A(_05333_),
    .B(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__nor2_1 _06190_ (.A(_05379_),
    .B(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__xnor2_1 _06191_ (.A(_05338_),
    .B(_05340_),
    .Y(_05383_));
 sky130_fd_sc_hd__or4_1 _06192_ (.A(_05377_),
    .B(_05378_),
    .C(_05381_),
    .D(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__a21oi_1 _06193_ (.A1(_05351_),
    .A2(_05374_),
    .B1(_05377_),
    .Y(_05385_));
 sky130_fd_sc_hd__o21ai_1 _06194_ (.A1(_05379_),
    .A2(_05381_),
    .B1(_05383_),
    .Y(_05386_));
 sky130_fd_sc_hd__nand2_1 _06195_ (.A(_05384_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__o21ai_1 _06196_ (.A1(_05385_),
    .A2(_05387_),
    .B1(_05384_),
    .Y(_05388_));
 sky130_fd_sc_hd__a211oi_1 _06197_ (.A1(_05342_),
    .A2(_05343_),
    .B1(_05334_),
    .C1(_05336_),
    .Y(_05389_));
 sky130_fd_sc_hd__inv_2 _06198_ (.A(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__nand2_1 _06199_ (.A(_05344_),
    .B(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__xnor2_1 _06200_ (.A(_05388_),
    .B(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__o21a_1 _06201_ (.A1(_05377_),
    .A2(_05378_),
    .B1(_05381_),
    .X(_05393_));
 sky130_fd_sc_hd__or2_1 _06202_ (.A(_05382_),
    .B(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__nor2_1 _06203_ (.A(_05373_),
    .B(_05352_),
    .Y(_05395_));
 sky130_fd_sc_hd__or2_2 _06204_ (.A(_05374_),
    .B(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__a21oi_1 _06205_ (.A1(net8),
    .A2(_05360_),
    .B1(_05358_),
    .Y(_05397_));
 sky130_fd_sc_hd__a21o_1 _06206_ (.A1(_05365_),
    .A2(_05367_),
    .B1(_05369_),
    .X(_05398_));
 sky130_fd_sc_hd__xnor2_1 _06207_ (.A(_05370_),
    .B(_05372_),
    .Y(_05399_));
 sky130_fd_sc_hd__and2_1 _06208_ (.A(net15),
    .B(net37),
    .X(_05400_));
 sky130_fd_sc_hd__and3_1 _06209_ (.A(net15),
    .B(net38),
    .C(net37),
    .X(_05401_));
 sky130_fd_sc_hd__o2bb2a_1 _06210_ (.A1_N(net13),
    .A2_N(net41),
    .B1(_05353_),
    .B2(_05354_),
    .X(_05402_));
 sky130_fd_sc_hd__and4bb_1 _06211_ (.A_N(_05355_),
    .B_N(_05402_),
    .C(_05400_),
    .D(net38),
    .X(_05403_));
 sky130_fd_sc_hd__and4_1 _06212_ (.A(net14),
    .B(net13),
    .C(net40),
    .D(net39),
    .X(_05404_));
 sky130_fd_sc_hd__a22oi_1 _06213_ (.A1(net13),
    .A2(net40),
    .B1(net39),
    .B2(net14),
    .Y(_05405_));
 sky130_fd_sc_hd__and4bb_1 _06214_ (.A_N(_05404_),
    .B_N(_05405_),
    .C(net11),
    .D(net41),
    .X(_05406_));
 sky130_fd_sc_hd__a41o_1 _06215_ (.A1(net14),
    .A2(net13),
    .A3(net40),
    .A4(net39),
    .B1(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__o2bb2a_1 _06216_ (.A1_N(net38),
    .A2_N(_05400_),
    .B1(_05402_),
    .B2(_05355_),
    .X(_05408_));
 sky130_fd_sc_hd__nor2_1 _06217_ (.A(_05403_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__a21o_1 _06218_ (.A1(_05409_),
    .A2(_05407_),
    .B1(_05403_),
    .X(_05410_));
 sky130_fd_sc_hd__a211o_1 _06219_ (.A1(_05311_),
    .A2(_05356_),
    .B1(_05355_),
    .C1(_05353_),
    .X(_00046_));
 sky130_fd_sc_hd__and3_1 _06220_ (.A(_05357_),
    .B(_05410_),
    .C(_00046_),
    .X(_00047_));
 sky130_fd_sc_hd__and4_1 _06221_ (.A(net43),
    .B(net11),
    .C(net42),
    .D(net10),
    .X(_00048_));
 sky130_fd_sc_hd__nand4_1 _06222_ (.A(net43),
    .B(net11),
    .C(net42),
    .D(net10),
    .Y(_00049_));
 sky130_fd_sc_hd__a22oi_1 _06223_ (.A1(net11),
    .A2(net42),
    .B1(net10),
    .B2(net43),
    .Y(_00050_));
 sky130_fd_sc_hd__or4_1 _06224_ (.A(_01054_),
    .B(_00050_),
    .C(_01076_),
    .D(_00048_),
    .X(_00051_));
 sky130_fd_sc_hd__o2bb2a_1 _06225_ (.A1_N(net45),
    .A2_N(net10),
    .B1(_05362_),
    .B2(_05363_),
    .X(_00052_));
 sky130_fd_sc_hd__o211a_1 _06226_ (.A1(_05364_),
    .A2(_00052_),
    .B1(_00051_),
    .C1(_00049_),
    .X(_00053_));
 sky130_fd_sc_hd__a211oi_2 _06227_ (.A1(_00049_),
    .A2(_00051_),
    .B1(_00052_),
    .C1(_05364_),
    .Y(_00054_));
 sky130_fd_sc_hd__and4_1 _06228_ (.A(net46),
    .B(net47),
    .C(net9),
    .D(net8),
    .X(_00055_));
 sky130_fd_sc_hd__nand4_1 _06229_ (.A(net46),
    .B(net47),
    .C(net9),
    .D(net8),
    .Y(_00056_));
 sky130_fd_sc_hd__a22o_1 _06230_ (.A1(net46),
    .A2(net9),
    .B1(net8),
    .B2(net47),
    .X(_00057_));
 sky130_fd_sc_hd__and3_1 _06231_ (.A(_00057_),
    .B(net7),
    .C(_00056_),
    .X(_00058_));
 sky130_fd_sc_hd__a21oi_1 _06232_ (.A1(_00056_),
    .A2(_00057_),
    .B1(net7),
    .Y(_00059_));
 sky130_fd_sc_hd__o22a_1 _06233_ (.A1(_00053_),
    .A2(_00054_),
    .B1(_00058_),
    .B2(_00059_),
    .X(_00060_));
 sky130_fd_sc_hd__nor4_1 _06234_ (.A(_00053_),
    .B(_00054_),
    .C(_00058_),
    .D(_00059_),
    .Y(_00061_));
 sky130_fd_sc_hd__nor2_1 _06235_ (.A(_00060_),
    .B(_00061_),
    .Y(_00062_));
 sky130_fd_sc_hd__a21oi_1 _06236_ (.A1(_05357_),
    .A2(_00046_),
    .B1(_05410_),
    .Y(_00063_));
 sky130_fd_sc_hd__nor2_1 _06237_ (.A(_00047_),
    .B(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__a21oi_1 _06238_ (.A1(_00062_),
    .A2(_00064_),
    .B1(_00047_),
    .Y(_00065_));
 sky130_fd_sc_hd__nor2_2 _06239_ (.A(_05399_),
    .B(_00065_),
    .Y(_00066_));
 sky130_fd_sc_hd__inv_2 _06240_ (.A(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__nor2_1 _06241_ (.A(_05398_),
    .B(_00066_),
    .Y(_00068_));
 sky130_fd_sc_hd__and2_1 _06242_ (.A(_00066_),
    .B(_05398_),
    .X(_00069_));
 sky130_fd_sc_hd__or2_1 _06243_ (.A(_00068_),
    .B(_00069_),
    .X(_00070_));
 sky130_fd_sc_hd__nor2_1 _06244_ (.A(_05397_),
    .B(_00070_),
    .Y(_00071_));
 sky130_fd_sc_hd__and2_1 _06245_ (.A(_00070_),
    .B(_05397_),
    .X(_00072_));
 sky130_fd_sc_hd__nor2_1 _06246_ (.A(_00071_),
    .B(_00072_),
    .Y(_00073_));
 sky130_fd_sc_hd__inv_2 _06247_ (.A(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__or2_1 _06248_ (.A(_05396_),
    .B(_00074_),
    .X(_00075_));
 sky130_fd_sc_hd__or3_2 _06249_ (.A(_05394_),
    .B(_05396_),
    .C(_00074_),
    .X(_00076_));
 sky130_fd_sc_hd__o21ai_2 _06250_ (.A1(_05396_),
    .A2(_00074_),
    .B1(_05394_),
    .Y(_00077_));
 sky130_fd_sc_hd__o211a_1 _06251_ (.A1(_00069_),
    .A2(_00071_),
    .B1(_00076_),
    .C1(_00077_),
    .X(_00078_));
 sky130_fd_sc_hd__o211ai_1 _06252_ (.A1(_00069_),
    .A2(_00071_),
    .B1(_00076_),
    .C1(_00077_),
    .Y(_00079_));
 sky130_fd_sc_hd__xnor2_1 _06253_ (.A(_05385_),
    .B(_05387_),
    .Y(_00080_));
 sky130_fd_sc_hd__a21oi_1 _06254_ (.A1(_00076_),
    .A2(_00079_),
    .B1(_00080_),
    .Y(_00081_));
 sky130_fd_sc_hd__o311a_1 _06255_ (.A1(_05394_),
    .A2(_05396_),
    .A3(_00074_),
    .B1(_00079_),
    .C1(_00080_),
    .X(_00082_));
 sky130_fd_sc_hd__nor2_1 _06256_ (.A(_00081_),
    .B(_00082_),
    .Y(_00083_));
 sky130_fd_sc_hd__or2_1 _06257_ (.A(_00054_),
    .B(_00061_),
    .X(_00084_));
 sky130_fd_sc_hd__xor2_1 _06258_ (.A(_00062_),
    .B(_00064_),
    .X(_00085_));
 sky130_fd_sc_hd__o2bb2a_1 _06259_ (.A1_N(net11),
    .A2_N(net41),
    .B1(_05404_),
    .B2(_05405_),
    .X(_00086_));
 sky130_fd_sc_hd__nand2_1 _06260_ (.A(net36),
    .B(_05400_),
    .Y(_00087_));
 sky130_fd_sc_hd__a21o_1 _06261_ (.A1(net15),
    .A2(net37),
    .B1(net36),
    .X(_00088_));
 sky130_fd_sc_hd__nand4_2 _06262_ (.A(_00087_),
    .B(_00088_),
    .C(net14),
    .D(net38),
    .Y(_00089_));
 sky130_fd_sc_hd__a211o_1 _06263_ (.A1(_00087_),
    .A2(_00089_),
    .B1(_05406_),
    .C1(_00086_),
    .X(_00090_));
 sky130_fd_sc_hd__and4_1 _06264_ (.A(net13),
    .B(net11),
    .C(net40),
    .D(net39),
    .X(_00091_));
 sky130_fd_sc_hd__a22oi_1 _06265_ (.A1(net11),
    .A2(net40),
    .B1(net39),
    .B2(net13),
    .Y(_00092_));
 sky130_fd_sc_hd__a22o_1 _06266_ (.A1(net11),
    .A2(net40),
    .B1(net39),
    .B2(net13),
    .X(_00093_));
 sky130_fd_sc_hd__and4b_1 _06267_ (.A_N(_00091_),
    .B(_00093_),
    .C(net10),
    .D(net41),
    .X(_00094_));
 sky130_fd_sc_hd__o211ai_1 _06268_ (.A1(_05406_),
    .A2(_00086_),
    .B1(_00087_),
    .C1(_00089_),
    .Y(_00095_));
 sky130_fd_sc_hd__and2_1 _06269_ (.A(_00090_),
    .B(_00095_),
    .X(_00096_));
 sky130_fd_sc_hd__o21ai_1 _06270_ (.A1(_00091_),
    .A2(_00094_),
    .B1(_00096_),
    .Y(_00097_));
 sky130_fd_sc_hd__xnor2_1 _06271_ (.A(_05407_),
    .B(_05409_),
    .Y(_00098_));
 sky130_fd_sc_hd__a21o_1 _06272_ (.A1(_00090_),
    .A2(_00097_),
    .B1(_00098_),
    .X(_00099_));
 sky130_fd_sc_hd__and4_1 _06273_ (.A(net43),
    .B(net42),
    .C(net10),
    .D(net9),
    .X(_00100_));
 sky130_fd_sc_hd__o2bb2a_1 _06274_ (.A1_N(net42),
    .A2_N(net10),
    .B1(_01076_),
    .B2(_01065_),
    .X(_00101_));
 sky130_fd_sc_hd__and4bb_1 _06275_ (.A_N(_00100_),
    .B_N(_00101_),
    .C(net45),
    .D(net8),
    .X(_00102_));
 sky130_fd_sc_hd__a2bb2o_1 _06276_ (.A1_N(_00048_),
    .A2_N(_00050_),
    .B1(net45),
    .B2(net9),
    .X(_00103_));
 sky130_fd_sc_hd__and2_1 _06277_ (.A(_00051_),
    .B(_00103_),
    .X(_00104_));
 sky130_fd_sc_hd__nor3_1 _06278_ (.A(_00100_),
    .B(_00102_),
    .C(_00104_),
    .Y(_00105_));
 sky130_fd_sc_hd__o21a_1 _06279_ (.A1(_00100_),
    .A2(_00102_),
    .B1(_00104_),
    .X(_00106_));
 sky130_fd_sc_hd__nor2_1 _06280_ (.A(_00105_),
    .B(_00106_),
    .Y(_00107_));
 sky130_fd_sc_hd__and4_1 _06281_ (.A(net46),
    .B(net47),
    .C(net8),
    .D(net7),
    .X(_00108_));
 sky130_fd_sc_hd__nand4_1 _06282_ (.A(net46),
    .B(net47),
    .C(net8),
    .D(net7),
    .Y(_00109_));
 sky130_fd_sc_hd__a22o_1 _06283_ (.A1(net46),
    .A2(net8),
    .B1(net7),
    .B2(net47),
    .X(_00110_));
 sky130_fd_sc_hd__and3_1 _06284_ (.A(_00110_),
    .B(net6),
    .C(_00109_),
    .X(_00111_));
 sky130_fd_sc_hd__a21oi_1 _06285_ (.A1(_00109_),
    .A2(_00110_),
    .B1(net6),
    .Y(_00112_));
 sky130_fd_sc_hd__nor2_1 _06286_ (.A(_00111_),
    .B(_00112_),
    .Y(_00113_));
 sky130_fd_sc_hd__xnor2_1 _06287_ (.A(_00107_),
    .B(_00113_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand3_1 _06288_ (.A(_00090_),
    .B(_00097_),
    .C(_00098_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_1 _06289_ (.A(_00099_),
    .B(_00115_),
    .Y(_00116_));
 sky130_fd_sc_hd__o21a_1 _06290_ (.A1(_00114_),
    .A2(_00116_),
    .B1(_00099_),
    .X(_00117_));
 sky130_fd_sc_hd__and2b_1 _06291_ (.A_N(_00117_),
    .B(_00085_),
    .X(_00118_));
 sky130_fd_sc_hd__nor2_1 _06292_ (.A(_00084_),
    .B(_00118_),
    .Y(_00119_));
 sky130_fd_sc_hd__o21a_1 _06293_ (.A1(_00054_),
    .A2(_00061_),
    .B1(_00118_),
    .X(_00120_));
 sky130_fd_sc_hd__nor2_1 _06294_ (.A(_00119_),
    .B(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__o21a_1 _06295_ (.A1(_00055_),
    .A2(_00058_),
    .B1(_00121_),
    .X(_00122_));
 sky130_fd_sc_hd__a211oi_1 _06296_ (.A1(_00057_),
    .A2(net7),
    .B1(_00055_),
    .C1(_00121_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _06297_ (.A(_00065_),
    .B(_05399_),
    .Y(_00124_));
 sky130_fd_sc_hd__nor4b_2 _06298_ (.A(_00066_),
    .B(_00122_),
    .C(_00123_),
    .D_N(_00124_),
    .Y(_00125_));
 sky130_fd_sc_hd__inv_2 _06299_ (.A(_00125_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _06300_ (.A(_05396_),
    .B(_00074_),
    .Y(_00127_));
 sky130_fd_sc_hd__nand3_2 _06301_ (.A(_00075_),
    .B(_00125_),
    .C(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__a21o_1 _06302_ (.A1(_00075_),
    .A2(_00127_),
    .B1(_00125_),
    .X(_00129_));
 sky130_fd_sc_hd__o211ai_2 _06303_ (.A1(_00120_),
    .A2(_00122_),
    .B1(_00128_),
    .C1(_00129_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _06304_ (.A(_00128_),
    .B(_00130_),
    .Y(_00131_));
 sky130_fd_sc_hd__a221oi_2 _06305_ (.A1(_05398_),
    .A2(_00066_),
    .B1(_00076_),
    .B2(_00077_),
    .C1(_00071_),
    .Y(_00132_));
 sky130_fd_sc_hd__nor2_1 _06306_ (.A(_00078_),
    .B(_00132_),
    .Y(_00133_));
 sky130_fd_sc_hd__a211oi_1 _06307_ (.A1(_00128_),
    .A2(_00130_),
    .B1(_00132_),
    .C1(_00078_),
    .Y(_00134_));
 sky130_fd_sc_hd__o211a_1 _06308_ (.A1(_00078_),
    .A2(_00132_),
    .B1(_00130_),
    .C1(_00128_),
    .X(_00135_));
 sky130_fd_sc_hd__or2_1 _06309_ (.A(_00134_),
    .B(_00135_),
    .X(_00136_));
 sky130_fd_sc_hd__a221o_1 _06310_ (.A1(_00118_),
    .A2(_00084_),
    .B1(_00129_),
    .B2(_00128_),
    .C1(_00122_),
    .X(_00137_));
 sky130_fd_sc_hd__and2_1 _06311_ (.A(_00130_),
    .B(_00137_),
    .X(_00138_));
 sky130_fd_sc_hd__and2b_1 _06312_ (.A_N(_00085_),
    .B(_00117_),
    .X(_00139_));
 sky130_fd_sc_hd__nor2_1 _06313_ (.A(_00118_),
    .B(_00139_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand4_2 _06314_ (.A(net15),
    .B(net14),
    .C(net37),
    .D(net36),
    .Y(_00141_));
 sky130_fd_sc_hd__a22o_1 _06315_ (.A1(net14),
    .A2(net37),
    .B1(net36),
    .B2(net15),
    .X(_00142_));
 sky130_fd_sc_hd__nand4_2 _06316_ (.A(_00142_),
    .B(net38),
    .C(net13),
    .D(_00141_),
    .Y(_00143_));
 sky130_fd_sc_hd__o2bb2a_1 _06317_ (.A1_N(net10),
    .A2_N(net41),
    .B1(_00091_),
    .B2(_00092_),
    .X(_00144_));
 sky130_fd_sc_hd__a211oi_1 _06318_ (.A1(_00141_),
    .A2(_00143_),
    .B1(_00144_),
    .C1(_00094_),
    .Y(_00145_));
 sky130_fd_sc_hd__and4_1 _06319_ (.A(net11),
    .B(net10),
    .C(net40),
    .D(net39),
    .X(_00146_));
 sky130_fd_sc_hd__a22oi_1 _06320_ (.A1(net10),
    .A2(net40),
    .B1(net39),
    .B2(net11),
    .Y(_00147_));
 sky130_fd_sc_hd__and4bb_1 _06321_ (.A_N(_00146_),
    .B_N(_00147_),
    .C(net41),
    .D(net9),
    .X(_00148_));
 sky130_fd_sc_hd__a41o_1 _06322_ (.A1(net11),
    .A2(net10),
    .A3(net40),
    .A4(net39),
    .B1(_00148_),
    .X(_00149_));
 sky130_fd_sc_hd__o211a_1 _06323_ (.A1(_00094_),
    .A2(_00144_),
    .B1(_00143_),
    .C1(_00141_),
    .X(_00150_));
 sky130_fd_sc_hd__nor2_1 _06324_ (.A(_00145_),
    .B(_00150_),
    .Y(_00151_));
 sky130_fd_sc_hd__o21a_1 _06325_ (.A1(_00146_),
    .A2(_00148_),
    .B1(_00151_),
    .X(_00152_));
 sky130_fd_sc_hd__a311o_1 _06326_ (.A1(net10),
    .A2(_00093_),
    .A3(net41),
    .B1(_00091_),
    .C1(_00096_),
    .X(_00153_));
 sky130_fd_sc_hd__and2_1 _06327_ (.A(_00097_),
    .B(_00153_),
    .X(_00154_));
 sky130_fd_sc_hd__o21ai_1 _06328_ (.A1(_00145_),
    .A2(_00152_),
    .B1(_00154_),
    .Y(_00155_));
 sky130_fd_sc_hd__and4_1 _06329_ (.A(net43),
    .B(net42),
    .C(net9),
    .D(net8),
    .X(_00156_));
 sky130_fd_sc_hd__nand4_1 _06330_ (.A(net43),
    .B(net42),
    .C(net9),
    .D(net8),
    .Y(_00157_));
 sky130_fd_sc_hd__a22oi_1 _06331_ (.A1(net42),
    .A2(net9),
    .B1(net8),
    .B2(net43),
    .Y(_00158_));
 sky130_fd_sc_hd__or4b_2 _06332_ (.A(_00158_),
    .B(_01054_),
    .C(_00156_),
    .D_N(net7),
    .X(_00159_));
 sky130_fd_sc_hd__o2bb2a_1 _06333_ (.A1_N(net45),
    .A2_N(net8),
    .B1(_00100_),
    .B2(_00101_),
    .X(_00160_));
 sky130_fd_sc_hd__o211a_1 _06334_ (.A1(_00102_),
    .A2(_00160_),
    .B1(_00159_),
    .C1(_00157_),
    .X(_00161_));
 sky130_fd_sc_hd__a211oi_2 _06335_ (.A1(_00157_),
    .A2(_00159_),
    .B1(_00160_),
    .C1(_00102_),
    .Y(_00162_));
 sky130_fd_sc_hd__and4_1 _06336_ (.A(net46),
    .B(net47),
    .C(net7),
    .D(net6),
    .X(_00163_));
 sky130_fd_sc_hd__a22oi_1 _06337_ (.A1(net46),
    .A2(net7),
    .B1(net6),
    .B2(net47),
    .Y(_00164_));
 sky130_fd_sc_hd__nor3_1 _06338_ (.A(_00164_),
    .B(_01098_),
    .C(_00163_),
    .Y(_00165_));
 sky130_fd_sc_hd__o21ai_1 _06339_ (.A1(_00163_),
    .A2(_00164_),
    .B1(_01098_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand2b_1 _06340_ (.A_N(_00165_),
    .B(_00166_),
    .Y(_00167_));
 sky130_fd_sc_hd__o21a_1 _06341_ (.A1(_00161_),
    .A2(_00162_),
    .B1(_00167_),
    .X(_00168_));
 sky130_fd_sc_hd__nor3_1 _06342_ (.A(_00167_),
    .B(_00162_),
    .C(_00161_),
    .Y(_00169_));
 sky130_fd_sc_hd__or2_1 _06343_ (.A(_00168_),
    .B(_00169_),
    .X(_00170_));
 sky130_fd_sc_hd__or3_1 _06344_ (.A(_00145_),
    .B(_00152_),
    .C(_00154_),
    .X(_00171_));
 sky130_fd_sc_hd__nand2_1 _06345_ (.A(_00155_),
    .B(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__o31a_1 _06346_ (.A1(_00168_),
    .A2(_00169_),
    .A3(_00172_),
    .B1(_00155_),
    .X(_00173_));
 sky130_fd_sc_hd__xnor2_1 _06347_ (.A(_00114_),
    .B(_00116_),
    .Y(_00174_));
 sky130_fd_sc_hd__nor2_1 _06348_ (.A(_00173_),
    .B(_00174_),
    .Y(_00175_));
 sky130_fd_sc_hd__o311a_1 _06349_ (.A1(_00168_),
    .A2(_00172_),
    .A3(_00169_),
    .B1(_00155_),
    .C1(_00174_),
    .X(_00176_));
 sky130_fd_sc_hd__or2_1 _06350_ (.A(_00175_),
    .B(_00176_),
    .X(_00177_));
 sky130_fd_sc_hd__nor2_1 _06351_ (.A(_01087_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__and2_1 _06352_ (.A(_00140_),
    .B(_00178_),
    .X(_00179_));
 sky130_fd_sc_hd__a21o_1 _06353_ (.A1(_00107_),
    .A2(_00113_),
    .B1(_00106_),
    .X(_00180_));
 sky130_fd_sc_hd__or2_1 _06354_ (.A(_00180_),
    .B(_00175_),
    .X(_00181_));
 sky130_fd_sc_hd__or3b_1 _06355_ (.A(_00173_),
    .B(_00174_),
    .C_N(_00180_),
    .X(_00182_));
 sky130_fd_sc_hd__o211a_1 _06356_ (.A1(_00108_),
    .A2(_00111_),
    .B1(_00181_),
    .C1(_00182_),
    .X(_00183_));
 sky130_fd_sc_hd__a211oi_1 _06357_ (.A1(_00181_),
    .A2(_00182_),
    .B1(_00108_),
    .C1(_00111_),
    .Y(_00184_));
 sky130_fd_sc_hd__or2_1 _06358_ (.A(_00140_),
    .B(_00178_),
    .X(_00185_));
 sky130_fd_sc_hd__inv_2 _06359_ (.A(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__nor4_1 _06360_ (.A(_00179_),
    .B(_00183_),
    .C(_00184_),
    .D(_00186_),
    .Y(_00187_));
 sky130_fd_sc_hd__a21o_1 _06361_ (.A1(_00140_),
    .A2(_00178_),
    .B1(_00187_),
    .X(_00188_));
 sky130_fd_sc_hd__a2bb2o_1 _06362_ (.A1_N(_00122_),
    .A2_N(_00123_),
    .B1(_00124_),
    .B2(_00067_),
    .X(_00189_));
 sky130_fd_sc_hd__and3_1 _06363_ (.A(_00126_),
    .B(_00188_),
    .C(_00189_),
    .X(_00190_));
 sky130_fd_sc_hd__a21oi_1 _06364_ (.A1(_00126_),
    .A2(_00189_),
    .B1(_00188_),
    .Y(_00191_));
 sky130_fd_sc_hd__or2_1 _06365_ (.A(_00190_),
    .B(_00191_),
    .X(_00192_));
 sky130_fd_sc_hd__a21oi_1 _06366_ (.A1(_00175_),
    .A2(_00180_),
    .B1(_00183_),
    .Y(_00193_));
 sky130_fd_sc_hd__nor2_1 _06367_ (.A(_00193_),
    .B(_00192_),
    .Y(_00194_));
 sky130_fd_sc_hd__o21ai_1 _06368_ (.A1(_00190_),
    .A2(_00194_),
    .B1(_00138_),
    .Y(_00195_));
 sky130_fd_sc_hd__a311o_1 _06369_ (.A1(_00126_),
    .A2(_00188_),
    .A3(_00189_),
    .B1(_00194_),
    .C1(_00138_),
    .X(_00196_));
 sky130_fd_sc_hd__nand2_1 _06370_ (.A(_00195_),
    .B(_00196_),
    .Y(_00197_));
 sky130_fd_sc_hd__xnor2_1 _06371_ (.A(_00192_),
    .B(_00193_),
    .Y(_00198_));
 sky130_fd_sc_hd__o2bb2a_1 _06372_ (.A1_N(net41),
    .A2_N(net9),
    .B1(_00146_),
    .B2(_00147_),
    .X(_00199_));
 sky130_fd_sc_hd__and4_1 _06373_ (.A(net14),
    .B(net13),
    .C(net37),
    .D(net36),
    .X(_00200_));
 sky130_fd_sc_hd__a22oi_2 _06374_ (.A1(net13),
    .A2(net37),
    .B1(net36),
    .B2(net14),
    .Y(_00201_));
 sky130_fd_sc_hd__a21oi_1 _06375_ (.A1(net11),
    .A2(net38),
    .B1(_00200_),
    .Y(_00202_));
 sky130_fd_sc_hd__or2_1 _06376_ (.A(_00201_),
    .B(_00202_),
    .X(_00203_));
 sky130_fd_sc_hd__or4_1 _06377_ (.A(_00148_),
    .B(_00199_),
    .C(_00201_),
    .D(_00202_),
    .X(_00204_));
 sky130_fd_sc_hd__and4_1 _06378_ (.A(net10),
    .B(net9),
    .C(net40),
    .D(net39),
    .X(_00205_));
 sky130_fd_sc_hd__a22oi_1 _06379_ (.A1(net9),
    .A2(net40),
    .B1(net39),
    .B2(net10),
    .Y(_00206_));
 sky130_fd_sc_hd__a22o_1 _06380_ (.A1(net9),
    .A2(net40),
    .B1(net39),
    .B2(net10),
    .X(_00207_));
 sky130_fd_sc_hd__and4b_1 _06381_ (.A_N(_00205_),
    .B(_00207_),
    .C(net41),
    .D(net8),
    .X(_00208_));
 sky130_fd_sc_hd__o21ai_1 _06382_ (.A1(_00148_),
    .A2(_00199_),
    .B1(_00203_),
    .Y(_00209_));
 sky130_fd_sc_hd__and2_1 _06383_ (.A(_00204_),
    .B(_00209_),
    .X(_00210_));
 sky130_fd_sc_hd__o21ai_2 _06384_ (.A1(_00205_),
    .A2(_00208_),
    .B1(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__nor2_1 _06385_ (.A(_00149_),
    .B(_00151_),
    .Y(_00212_));
 sky130_fd_sc_hd__or2_1 _06386_ (.A(_00152_),
    .B(_00212_),
    .X(_00213_));
 sky130_fd_sc_hd__a21oi_1 _06387_ (.A1(_00204_),
    .A2(_00211_),
    .B1(_00213_),
    .Y(_00214_));
 sky130_fd_sc_hd__a21o_1 _06388_ (.A1(_00204_),
    .A2(_00211_),
    .B1(_00213_),
    .X(_00215_));
 sky130_fd_sc_hd__and4_1 _06389_ (.A(net43),
    .B(net42),
    .C(net8),
    .D(net7),
    .X(_00216_));
 sky130_fd_sc_hd__a22oi_1 _06390_ (.A1(net42),
    .A2(net8),
    .B1(net7),
    .B2(net43),
    .Y(_00217_));
 sky130_fd_sc_hd__and4bb_1 _06391_ (.A_N(_00216_),
    .B_N(_00217_),
    .C(net45),
    .D(net6),
    .X(_00218_));
 sky130_fd_sc_hd__a2bb2o_1 _06392_ (.A1_N(_00156_),
    .A2_N(_00158_),
    .B1(net45),
    .B2(net7),
    .X(_00219_));
 sky130_fd_sc_hd__o211ai_1 _06393_ (.A1(_00216_),
    .A2(_00218_),
    .B1(_00219_),
    .C1(_00159_),
    .Y(_00220_));
 sky130_fd_sc_hd__a211o_1 _06394_ (.A1(_00159_),
    .A2(_00219_),
    .B1(_00218_),
    .C1(_00216_),
    .X(_00221_));
 sky130_fd_sc_hd__and4_1 _06395_ (.A(net46),
    .B(net47),
    .C(net6),
    .D(net5),
    .X(_00222_));
 sky130_fd_sc_hd__o2bb2a_1 _06396_ (.A1_N(net46),
    .A2_N(net6),
    .B1(_01098_),
    .B2(_01043_),
    .X(_00223_));
 sky130_fd_sc_hd__nor2_1 _06397_ (.A(_00222_),
    .B(_00223_),
    .Y(_00224_));
 sky130_fd_sc_hd__xor2_1 _06398_ (.A(net4),
    .B(_00224_),
    .X(_00225_));
 sky130_fd_sc_hd__and3_1 _06399_ (.A(_00220_),
    .B(_00221_),
    .C(_00225_),
    .X(_00226_));
 sky130_fd_sc_hd__a21o_1 _06400_ (.A1(_00220_),
    .A2(_00221_),
    .B1(_00225_),
    .X(_00227_));
 sky130_fd_sc_hd__nand2b_1 _06401_ (.A_N(_00226_),
    .B(_00227_),
    .Y(_00228_));
 sky130_fd_sc_hd__o311a_1 _06402_ (.A1(_00148_),
    .A2(_00199_),
    .A3(_00203_),
    .B1(_00211_),
    .C1(_00213_),
    .X(_00229_));
 sky130_fd_sc_hd__nor2_1 _06403_ (.A(_00214_),
    .B(_00229_),
    .Y(_00230_));
 sky130_fd_sc_hd__o21ai_1 _06404_ (.A1(_00228_),
    .A2(_00229_),
    .B1(_00215_),
    .Y(_00231_));
 sky130_fd_sc_hd__a22o_1 _06405_ (.A1(net14),
    .A2(net38),
    .B1(_00087_),
    .B2(_00088_),
    .X(_00232_));
 sky130_fd_sc_hd__and2_2 _06406_ (.A(net15),
    .B(net34),
    .X(_00233_));
 sky130_fd_sc_hd__and3_1 _06407_ (.A(net15),
    .B(net35),
    .C(net34),
    .X(_00234_));
 sky130_fd_sc_hd__a22o_1 _06408_ (.A1(net13),
    .A2(net38),
    .B1(_00141_),
    .B2(_00142_),
    .X(_00235_));
 sky130_fd_sc_hd__and4b_1 _06409_ (.A_N(_00233_),
    .B(net35),
    .C(_00143_),
    .D(_00235_),
    .X(_00236_));
 sky130_fd_sc_hd__o211ai_1 _06410_ (.A1(_00234_),
    .A2(_00236_),
    .B1(_00089_),
    .C1(_00232_),
    .Y(_00237_));
 sky130_fd_sc_hd__xnor2_1 _06411_ (.A(_00170_),
    .B(_00172_),
    .Y(_00238_));
 sky130_fd_sc_hd__or2_1 _06412_ (.A(_00237_),
    .B(_00238_),
    .X(_00239_));
 sky130_fd_sc_hd__nand2_1 _06413_ (.A(_00237_),
    .B(_00238_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _06414_ (.A(_00239_),
    .B(_00240_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2b_1 _06415_ (.A_N(_00241_),
    .B(_00231_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2b_1 _06416_ (.A_N(_00231_),
    .B(_00241_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _06417_ (.A(_00242_),
    .B(_00243_),
    .Y(_00244_));
 sky130_fd_sc_hd__a21oi_1 _06418_ (.A1(net15),
    .A2(net38),
    .B1(net37),
    .Y(_00245_));
 sky130_fd_sc_hd__or3_1 _06419_ (.A(_05401_),
    .B(_00245_),
    .C(_00244_),
    .X(_00246_));
 sky130_fd_sc_hd__and2_1 _06420_ (.A(_01087_),
    .B(_00177_),
    .X(_00247_));
 sky130_fd_sc_hd__or2_1 _06421_ (.A(_00178_),
    .B(_00247_),
    .X(_00248_));
 sky130_fd_sc_hd__or4_1 _06422_ (.A(_05401_),
    .B(_00244_),
    .C(_00245_),
    .D(_00248_),
    .X(_00249_));
 sky130_fd_sc_hd__or4bb_1 _06423_ (.A(_00162_),
    .B(_00169_),
    .C_N(_00239_),
    .D_N(_00242_),
    .X(_00250_));
 sky130_fd_sc_hd__a2bb2o_1 _06424_ (.A1_N(_00162_),
    .A2_N(_00169_),
    .B1(_00239_),
    .B2(_00242_),
    .X(_00251_));
 sky130_fd_sc_hd__o211ai_2 _06425_ (.A1(_00163_),
    .A2(_00165_),
    .B1(_00250_),
    .C1(_00251_),
    .Y(_00252_));
 sky130_fd_sc_hd__a211o_1 _06426_ (.A1(_00250_),
    .A2(_00251_),
    .B1(_00163_),
    .C1(_00165_),
    .X(_00253_));
 sky130_fd_sc_hd__nand2_1 _06427_ (.A(_00252_),
    .B(_00253_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _06428_ (.A(_00246_),
    .B(_00248_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _06429_ (.A(_00249_),
    .B(_00255_),
    .Y(_00256_));
 sky130_fd_sc_hd__o21ai_1 _06430_ (.A1(_00254_),
    .A2(_00256_),
    .B1(_00249_),
    .Y(_00257_));
 sky130_fd_sc_hd__o22a_1 _06431_ (.A1(_00183_),
    .A2(_00184_),
    .B1(_00186_),
    .B2(_00179_),
    .X(_00258_));
 sky130_fd_sc_hd__nor2_1 _06432_ (.A(_00187_),
    .B(_00258_),
    .Y(_00259_));
 sky130_fd_sc_hd__xnor2_1 _06433_ (.A(_00257_),
    .B(_00259_),
    .Y(_00260_));
 sky130_fd_sc_hd__a21oi_1 _06434_ (.A1(_00251_),
    .A2(_00252_),
    .B1(_00260_),
    .Y(_00261_));
 sky130_fd_sc_hd__a21oi_1 _06435_ (.A1(_00257_),
    .A2(_00259_),
    .B1(_00261_),
    .Y(_00262_));
 sky130_fd_sc_hd__nor2_1 _06436_ (.A(_00262_),
    .B(_00198_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _06437_ (.A(_00198_),
    .B(_00262_),
    .Y(_00264_));
 sky130_fd_sc_hd__and4_1 _06438_ (.A(net13),
    .B(net11),
    .C(net37),
    .D(net36),
    .X(_00265_));
 sky130_fd_sc_hd__a22oi_1 _06439_ (.A1(net11),
    .A2(net37),
    .B1(net36),
    .B2(net13),
    .Y(_00266_));
 sky130_fd_sc_hd__a22o_1 _06440_ (.A1(net11),
    .A2(net37),
    .B1(net36),
    .B2(net13),
    .X(_00267_));
 sky130_fd_sc_hd__a31oi_1 _06441_ (.A1(_00267_),
    .A2(net38),
    .A3(net10),
    .B1(_00265_),
    .Y(_00268_));
 sky130_fd_sc_hd__o2bb2a_1 _06442_ (.A1_N(net41),
    .A2_N(net8),
    .B1(_00205_),
    .B2(_00206_),
    .X(_00269_));
 sky130_fd_sc_hd__nor3_1 _06443_ (.A(_00208_),
    .B(_00268_),
    .C(_00269_),
    .Y(_00270_));
 sky130_fd_sc_hd__and4_1 _06444_ (.A(net9),
    .B(net40),
    .C(net8),
    .D(net39),
    .X(_00271_));
 sky130_fd_sc_hd__a22oi_1 _06445_ (.A1(net40),
    .A2(net8),
    .B1(net39),
    .B2(net9),
    .Y(_00272_));
 sky130_fd_sc_hd__a22o_1 _06446_ (.A1(net40),
    .A2(net8),
    .B1(net39),
    .B2(net9),
    .X(_00273_));
 sky130_fd_sc_hd__and4b_1 _06447_ (.A_N(_00271_),
    .B(_00273_),
    .C(net41),
    .D(net7),
    .X(_00274_));
 sky130_fd_sc_hd__a31o_1 _06448_ (.A1(_00273_),
    .A2(net7),
    .A3(net41),
    .B1(_00271_),
    .X(_00275_));
 sky130_fd_sc_hd__o21a_1 _06449_ (.A1(_00208_),
    .A2(_00269_),
    .B1(_00268_),
    .X(_00276_));
 sky130_fd_sc_hd__nor2_1 _06450_ (.A(_00270_),
    .B(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__o21a_1 _06451_ (.A1(_00271_),
    .A2(_00274_),
    .B1(_00277_),
    .X(_00278_));
 sky130_fd_sc_hd__a311o_1 _06452_ (.A1(net41),
    .A2(_00207_),
    .A3(net8),
    .B1(_00205_),
    .C1(_00210_),
    .X(_00279_));
 sky130_fd_sc_hd__o211ai_2 _06453_ (.A1(_00270_),
    .A2(_00278_),
    .B1(_00279_),
    .C1(_00211_),
    .Y(_00280_));
 sky130_fd_sc_hd__and4_1 _06454_ (.A(net43),
    .B(net42),
    .C(net7),
    .D(net6),
    .X(_00281_));
 sky130_fd_sc_hd__nand4_2 _06455_ (.A(net43),
    .B(net42),
    .C(net7),
    .D(net6),
    .Y(_00282_));
 sky130_fd_sc_hd__a22oi_2 _06456_ (.A1(net42),
    .A2(net7),
    .B1(net6),
    .B2(net43),
    .Y(_00283_));
 sky130_fd_sc_hd__and4b_1 _06457_ (.A_N(_00283_),
    .B(net5),
    .C(net45),
    .D(_00282_),
    .X(_00284_));
 sky130_fd_sc_hd__or4_1 _06458_ (.A(_01054_),
    .B(_00283_),
    .C(_01098_),
    .D(_00281_),
    .X(_00285_));
 sky130_fd_sc_hd__o2bb2a_1 _06459_ (.A1_N(net45),
    .A2_N(net6),
    .B1(_00216_),
    .B2(_00217_),
    .X(_00286_));
 sky130_fd_sc_hd__o211a_1 _06460_ (.A1(_00218_),
    .A2(_00286_),
    .B1(_00285_),
    .C1(_00282_),
    .X(_00287_));
 sky130_fd_sc_hd__a211oi_2 _06461_ (.A1(_00282_),
    .A2(_00285_),
    .B1(_00286_),
    .C1(_00218_),
    .Y(_00288_));
 sky130_fd_sc_hd__and4_1 _06462_ (.A(net46),
    .B(net47),
    .C(net5),
    .D(net4),
    .X(_00289_));
 sky130_fd_sc_hd__a22oi_2 _06463_ (.A1(net46),
    .A2(net5),
    .B1(net4),
    .B2(net47),
    .Y(_00290_));
 sky130_fd_sc_hd__o21ai_1 _06464_ (.A1(_00289_),
    .A2(_00290_),
    .B1(net3),
    .Y(_00291_));
 sky130_fd_sc_hd__or3_1 _06465_ (.A(net3),
    .B(_00289_),
    .C(_00290_),
    .X(_00292_));
 sky130_fd_sc_hd__o211ai_1 _06466_ (.A1(_00287_),
    .A2(_00288_),
    .B1(_00291_),
    .C1(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__a211oi_1 _06467_ (.A1(_00291_),
    .A2(_00292_),
    .B1(_00287_),
    .C1(_00288_),
    .Y(_00294_));
 sky130_fd_sc_hd__a211o_1 _06468_ (.A1(_00291_),
    .A2(_00292_),
    .B1(_00287_),
    .C1(_00288_),
    .X(_00295_));
 sky130_fd_sc_hd__a221o_1 _06469_ (.A1(_00275_),
    .A2(_00277_),
    .B1(_00279_),
    .B2(_00211_),
    .C1(_00270_),
    .X(_00296_));
 sky130_fd_sc_hd__and2_1 _06470_ (.A(_00280_),
    .B(_00296_),
    .X(_00297_));
 sky130_fd_sc_hd__nand3_1 _06471_ (.A(_00297_),
    .B(_00295_),
    .C(_00293_),
    .Y(_00298_));
 sky130_fd_sc_hd__a2bb2o_1 _06472_ (.A1_N(_00233_),
    .A2_N(_01109_),
    .B1(_00143_),
    .B2(_00235_),
    .X(_00299_));
 sky130_fd_sc_hd__nand2b_1 _06473_ (.A_N(_00236_),
    .B(_00299_),
    .Y(_00300_));
 sky130_fd_sc_hd__a21oi_1 _06474_ (.A1(net15),
    .A2(net35),
    .B1(net34),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _06475_ (.A(net64),
    .B(_00233_),
    .Y(_00302_));
 sky130_fd_sc_hd__a21o_1 _06476_ (.A1(net15),
    .A2(net34),
    .B1(net64),
    .X(_00303_));
 sky130_fd_sc_hd__nand4_2 _06477_ (.A(_00302_),
    .B(_00303_),
    .C(net14),
    .D(net35),
    .Y(_00304_));
 sky130_fd_sc_hd__a221o_1 _06478_ (.A1(net35),
    .A2(_00233_),
    .B1(_00302_),
    .B2(_00304_),
    .C1(_00301_),
    .X(_00305_));
 sky130_fd_sc_hd__o211ai_1 _06479_ (.A1(_00234_),
    .A2(_00301_),
    .B1(_00302_),
    .C1(_00304_),
    .Y(_00306_));
 sky130_fd_sc_hd__and2_1 _06480_ (.A(_00305_),
    .B(_00306_),
    .X(_00307_));
 sky130_fd_sc_hd__o211a_1 _06481_ (.A1(_00200_),
    .A2(_00201_),
    .B1(net11),
    .C1(net38),
    .X(_00308_));
 sky130_fd_sc_hd__a211oi_1 _06482_ (.A1(net11),
    .A2(net38),
    .B1(_00200_),
    .C1(_00201_),
    .Y(_00309_));
 sky130_fd_sc_hd__o21ai_1 _06483_ (.A1(_00308_),
    .A2(_00309_),
    .B1(_00307_),
    .Y(_00310_));
 sky130_fd_sc_hd__and2_1 _06484_ (.A(_00305_),
    .B(_00310_),
    .X(_00311_));
 sky130_fd_sc_hd__a21oi_1 _06485_ (.A1(_00305_),
    .A2(_00310_),
    .B1(_00300_),
    .Y(_00312_));
 sky130_fd_sc_hd__xor2_1 _06486_ (.A(_00228_),
    .B(_00230_),
    .X(_00313_));
 sky130_fd_sc_hd__xor2_1 _06487_ (.A(_00312_),
    .B(_00313_),
    .X(_00314_));
 sky130_fd_sc_hd__a21o_1 _06488_ (.A1(_00280_),
    .A2(_00298_),
    .B1(_00314_),
    .X(_00315_));
 sky130_fd_sc_hd__nand3_1 _06489_ (.A(_00280_),
    .B(_00298_),
    .C(_00314_),
    .Y(_00316_));
 sky130_fd_sc_hd__and2_1 _06490_ (.A(_00315_),
    .B(_00316_),
    .X(_00317_));
 sky130_fd_sc_hd__a221o_1 _06491_ (.A1(_00089_),
    .A2(_00232_),
    .B1(_00233_),
    .B2(net35),
    .C1(_00236_),
    .X(_00318_));
 sky130_fd_sc_hd__and2_1 _06492_ (.A(_00237_),
    .B(_00318_),
    .X(_00319_));
 sky130_fd_sc_hd__nand2_1 _06493_ (.A(_00317_),
    .B(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__o21ai_1 _06494_ (.A1(_05401_),
    .A2(_00245_),
    .B1(_00244_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _06495_ (.A(_00246_),
    .B(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__or2_1 _06496_ (.A(_00320_),
    .B(_00322_),
    .X(_00323_));
 sky130_fd_sc_hd__a21oi_1 _06497_ (.A1(net4),
    .A2(_00224_),
    .B1(_00222_),
    .Y(_00324_));
 sky130_fd_sc_hd__a21bo_1 _06498_ (.A1(_00221_),
    .A2(_00225_),
    .B1_N(_00220_),
    .X(_00325_));
 sky130_fd_sc_hd__o31ai_2 _06499_ (.A1(_00300_),
    .A2(_00311_),
    .A3(_00313_),
    .B1(_00315_),
    .Y(_00326_));
 sky130_fd_sc_hd__xnor2_1 _06500_ (.A(_00325_),
    .B(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__nor2_1 _06501_ (.A(_00324_),
    .B(_00327_),
    .Y(_00328_));
 sky130_fd_sc_hd__and2_1 _06502_ (.A(_00327_),
    .B(_00324_),
    .X(_00329_));
 sky130_fd_sc_hd__nand2_1 _06503_ (.A(_00320_),
    .B(_00322_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _06504_ (.A(_00323_),
    .B(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__or3_1 _06505_ (.A(_00328_),
    .B(_00329_),
    .C(_00331_),
    .X(_00332_));
 sky130_fd_sc_hd__xnor2_1 _06506_ (.A(_00254_),
    .B(_00256_),
    .Y(_00333_));
 sky130_fd_sc_hd__a21oi_1 _06507_ (.A1(_00323_),
    .A2(_00332_),
    .B1(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__a21o_1 _06508_ (.A1(_00325_),
    .A2(_00326_),
    .B1(_00328_),
    .X(_00335_));
 sky130_fd_sc_hd__o311a_1 _06509_ (.A1(_00328_),
    .A2(_00331_),
    .A3(_00329_),
    .B1(_00323_),
    .C1(_00333_),
    .X(_00336_));
 sky130_fd_sc_hd__nor2_1 _06510_ (.A(_00334_),
    .B(_00336_),
    .Y(_00337_));
 sky130_fd_sc_hd__a21oi_1 _06511_ (.A1(_00337_),
    .A2(_00335_),
    .B1(_00334_),
    .Y(_00338_));
 sky130_fd_sc_hd__and3_1 _06512_ (.A(_00251_),
    .B(_00252_),
    .C(_00260_),
    .X(_00339_));
 sky130_fd_sc_hd__nor2_1 _06513_ (.A(_00261_),
    .B(_00339_),
    .Y(_00340_));
 sky130_fd_sc_hd__and2b_1 _06514_ (.A_N(_00338_),
    .B(_00340_),
    .X(_00341_));
 sky130_fd_sc_hd__and4_1 _06515_ (.A(net11),
    .B(net10),
    .C(net37),
    .D(net36),
    .X(_00342_));
 sky130_fd_sc_hd__nand4_1 _06516_ (.A(net11),
    .B(net10),
    .C(net37),
    .D(net36),
    .Y(_00343_));
 sky130_fd_sc_hd__a22oi_1 _06517_ (.A1(net10),
    .A2(net37),
    .B1(net36),
    .B2(net11),
    .Y(_00344_));
 sky130_fd_sc_hd__or4_2 _06518_ (.A(_01076_),
    .B(_00344_),
    .C(_01087_),
    .D(_00342_),
    .X(_00345_));
 sky130_fd_sc_hd__o2bb2a_1 _06519_ (.A1_N(net41),
    .A2_N(net7),
    .B1(_00271_),
    .B2(_00272_),
    .X(_00346_));
 sky130_fd_sc_hd__a211oi_2 _06520_ (.A1(_00343_),
    .A2(_00345_),
    .B1(_00346_),
    .C1(_00274_),
    .Y(_00347_));
 sky130_fd_sc_hd__and4_1 _06521_ (.A(net40),
    .B(net8),
    .C(net39),
    .D(net7),
    .X(_00348_));
 sky130_fd_sc_hd__a22oi_1 _06522_ (.A1(net8),
    .A2(net39),
    .B1(net7),
    .B2(net40),
    .Y(_00349_));
 sky130_fd_sc_hd__a22o_1 _06523_ (.A1(net8),
    .A2(net39),
    .B1(net7),
    .B2(net40),
    .X(_00350_));
 sky130_fd_sc_hd__and4b_1 _06524_ (.A_N(_00348_),
    .B(_00350_),
    .C(net41),
    .D(net6),
    .X(_00351_));
 sky130_fd_sc_hd__a31o_1 _06525_ (.A1(_00350_),
    .A2(net6),
    .A3(net41),
    .B1(_00348_),
    .X(_00352_));
 sky130_fd_sc_hd__o211a_1 _06526_ (.A1(_00274_),
    .A2(_00346_),
    .B1(_00345_),
    .C1(_00343_),
    .X(_00353_));
 sky130_fd_sc_hd__nor2_1 _06527_ (.A(_00347_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__o21a_1 _06528_ (.A1(_00348_),
    .A2(_00351_),
    .B1(_00354_),
    .X(_00355_));
 sky130_fd_sc_hd__nor2_1 _06529_ (.A(_00275_),
    .B(_00277_),
    .Y(_00356_));
 sky130_fd_sc_hd__nor2_1 _06530_ (.A(_00278_),
    .B(_00356_),
    .Y(_00357_));
 sky130_fd_sc_hd__o21ai_2 _06531_ (.A1(_00347_),
    .A2(_00355_),
    .B1(_00357_),
    .Y(_00358_));
 sky130_fd_sc_hd__and4_1 _06532_ (.A(net43),
    .B(net42),
    .C(net6),
    .D(net5),
    .X(_00359_));
 sky130_fd_sc_hd__nand4_2 _06533_ (.A(net43),
    .B(net42),
    .C(net6),
    .D(net5),
    .Y(_00360_));
 sky130_fd_sc_hd__o2bb2a_1 _06534_ (.A1_N(net42),
    .A2_N(net6),
    .B1(_01098_),
    .B2(_01065_),
    .X(_00361_));
 sky130_fd_sc_hd__and4b_1 _06535_ (.A_N(_00361_),
    .B(net4),
    .C(net45),
    .D(_00360_),
    .X(_00362_));
 sky130_fd_sc_hd__or4b_1 _06536_ (.A(_01054_),
    .B(_00359_),
    .C(_00361_),
    .D_N(net4),
    .X(_00363_));
 sky130_fd_sc_hd__o22a_1 _06537_ (.A1(_01054_),
    .A2(_01098_),
    .B1(_00281_),
    .B2(_00283_),
    .X(_00364_));
 sky130_fd_sc_hd__o211a_1 _06538_ (.A1(_00284_),
    .A2(_00364_),
    .B1(_00363_),
    .C1(_00360_),
    .X(_00365_));
 sky130_fd_sc_hd__a211oi_2 _06539_ (.A1(_00360_),
    .A2(_00363_),
    .B1(_00364_),
    .C1(_00284_),
    .Y(_00366_));
 sky130_fd_sc_hd__nor2_1 _06540_ (.A(_00365_),
    .B(_00366_),
    .Y(_00367_));
 sky130_fd_sc_hd__and4_1 _06541_ (.A(net46),
    .B(net47),
    .C(net4),
    .D(net3),
    .X(_00368_));
 sky130_fd_sc_hd__o2bb2a_1 _06542_ (.A1_N(net46),
    .A2_N(net4),
    .B1(_01120_),
    .B2(_01043_),
    .X(_00369_));
 sky130_fd_sc_hd__nor3_1 _06543_ (.A(_01131_),
    .B(_00368_),
    .C(_00369_),
    .Y(_00370_));
 sky130_fd_sc_hd__o21ai_1 _06544_ (.A1(_00368_),
    .A2(_00369_),
    .B1(_01131_),
    .Y(_00371_));
 sky130_fd_sc_hd__nand2b_1 _06545_ (.A_N(_00370_),
    .B(_00371_),
    .Y(_00372_));
 sky130_fd_sc_hd__nor3_1 _06546_ (.A(_00365_),
    .B(_00372_),
    .C(_00366_),
    .Y(_00373_));
 sky130_fd_sc_hd__xor2_1 _06547_ (.A(_00367_),
    .B(_00372_),
    .X(_00374_));
 sky130_fd_sc_hd__or3_1 _06548_ (.A(_00347_),
    .B(_00355_),
    .C(_00357_),
    .X(_00375_));
 sky130_fd_sc_hd__nand2_1 _06549_ (.A(_00358_),
    .B(_00375_),
    .Y(_00376_));
 sky130_fd_sc_hd__or2_1 _06550_ (.A(_00374_),
    .B(_00376_),
    .X(_00377_));
 sky130_fd_sc_hd__and3_1 _06551_ (.A(net14),
    .B(net64),
    .C(_00233_),
    .X(_00378_));
 sky130_fd_sc_hd__a22oi_1 _06552_ (.A1(net14),
    .A2(net34),
    .B1(net64),
    .B2(net15),
    .Y(_00379_));
 sky130_fd_sc_hd__and4bb_1 _06553_ (.A_N(_00378_),
    .B_N(_00379_),
    .C(net13),
    .D(net35),
    .X(_00380_));
 sky130_fd_sc_hd__a31o_1 _06554_ (.A1(net14),
    .A2(net64),
    .A3(_00233_),
    .B1(_00380_),
    .X(_00381_));
 sky130_fd_sc_hd__a22o_1 _06555_ (.A1(net14),
    .A2(net35),
    .B1(_00302_),
    .B2(_00303_),
    .X(_00382_));
 sky130_fd_sc_hd__and3_1 _06556_ (.A(_00304_),
    .B(_00381_),
    .C(_00382_),
    .X(_00383_));
 sky130_fd_sc_hd__a21oi_1 _06557_ (.A1(_00304_),
    .A2(_00382_),
    .B1(_00381_),
    .Y(_00384_));
 sky130_fd_sc_hd__nor2_1 _06558_ (.A(_00383_),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__a211o_1 _06559_ (.A1(net10),
    .A2(net38),
    .B1(_00265_),
    .C1(_00266_),
    .X(_00386_));
 sky130_fd_sc_hd__o211ai_1 _06560_ (.A1(_00265_),
    .A2(_00266_),
    .B1(net10),
    .C1(net38),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _06561_ (.A(_00386_),
    .B(_00387_),
    .Y(_00388_));
 sky130_fd_sc_hd__and2_1 _06562_ (.A(_00385_),
    .B(_00388_),
    .X(_00389_));
 sky130_fd_sc_hd__a31o_1 _06563_ (.A1(_00304_),
    .A2(_00381_),
    .A3(_00382_),
    .B1(_00389_),
    .X(_00390_));
 sky130_fd_sc_hd__or3_1 _06564_ (.A(_00307_),
    .B(_00308_),
    .C(_00309_),
    .X(_00391_));
 sky130_fd_sc_hd__and2_1 _06565_ (.A(_00310_),
    .B(_00391_),
    .X(_00392_));
 sky130_fd_sc_hd__nand2_1 _06566_ (.A(_00390_),
    .B(_00392_),
    .Y(_00393_));
 sky130_fd_sc_hd__a21o_1 _06567_ (.A1(_00293_),
    .A2(_00295_),
    .B1(_00297_),
    .X(_00394_));
 sky130_fd_sc_hd__nand2_1 _06568_ (.A(_00298_),
    .B(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__or2_1 _06569_ (.A(_00393_),
    .B(_00395_),
    .X(_00396_));
 sky130_fd_sc_hd__nand2_1 _06570_ (.A(_00393_),
    .B(_00395_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _06571_ (.A(_00396_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__and3_1 _06572_ (.A(_00358_),
    .B(_00377_),
    .C(_00398_),
    .X(_00399_));
 sky130_fd_sc_hd__a21o_1 _06573_ (.A1(_00358_),
    .A2(_00377_),
    .B1(_00398_),
    .X(_00400_));
 sky130_fd_sc_hd__and2b_1 _06574_ (.A_N(_00399_),
    .B(_00400_),
    .X(_00401_));
 sky130_fd_sc_hd__nand2_1 _06575_ (.A(_00311_),
    .B(_00300_),
    .Y(_00402_));
 sky130_fd_sc_hd__and2b_1 _06576_ (.A_N(_00312_),
    .B(_00402_),
    .X(_00403_));
 sky130_fd_sc_hd__nand2_1 _06577_ (.A(_00401_),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__or2_1 _06578_ (.A(_00317_),
    .B(_00319_),
    .X(_00405_));
 sky130_fd_sc_hd__nand2_1 _06579_ (.A(_00320_),
    .B(_00405_),
    .Y(_00406_));
 sky130_fd_sc_hd__xnor2_1 _06580_ (.A(_00404_),
    .B(_00406_),
    .Y(_00407_));
 sky130_fd_sc_hd__o21ba_1 _06581_ (.A1(_01120_),
    .A2(_00290_),
    .B1_N(_00289_),
    .X(_00408_));
 sky130_fd_sc_hd__or4bb_1 _06582_ (.A(_00288_),
    .B(_00294_),
    .C_N(_00396_),
    .D_N(_00400_),
    .X(_00409_));
 sky130_fd_sc_hd__a2bb2o_1 _06583_ (.A1_N(_00288_),
    .A2_N(_00294_),
    .B1(_00396_),
    .B2(_00400_),
    .X(_00410_));
 sky130_fd_sc_hd__nand2_1 _06584_ (.A(_00409_),
    .B(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__or2_1 _06585_ (.A(_00408_),
    .B(_00411_),
    .X(_00412_));
 sky130_fd_sc_hd__and2_1 _06586_ (.A(_00411_),
    .B(_00408_),
    .X(_00413_));
 sky130_fd_sc_hd__inv_2 _06587_ (.A(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__nand2_1 _06588_ (.A(_00412_),
    .B(_00414_),
    .Y(_00415_));
 sky130_fd_sc_hd__or3b_1 _06589_ (.A(_00413_),
    .B(_00407_),
    .C_N(_00412_),
    .X(_00416_));
 sky130_fd_sc_hd__o21ai_1 _06590_ (.A1(_00404_),
    .A2(_00406_),
    .B1(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__o21ai_1 _06591_ (.A1(_00328_),
    .A2(_00329_),
    .B1(_00331_),
    .Y(_00418_));
 sky130_fd_sc_hd__and2_1 _06592_ (.A(_00332_),
    .B(_00418_),
    .X(_00419_));
 sky130_fd_sc_hd__xnor2_1 _06593_ (.A(_00417_),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__a21o_1 _06594_ (.A1(_00410_),
    .A2(_00412_),
    .B1(_00420_),
    .X(_00421_));
 sky130_fd_sc_hd__a21bo_1 _06595_ (.A1(_00417_),
    .A2(_00419_),
    .B1_N(_00421_),
    .X(_00422_));
 sky130_fd_sc_hd__xor2_1 _06596_ (.A(_00335_),
    .B(_00337_),
    .X(_00423_));
 sky130_fd_sc_hd__xnor2_1 _06597_ (.A(_00422_),
    .B(_00423_),
    .Y(_00424_));
 sky130_fd_sc_hd__and4_1 _06598_ (.A(net10),
    .B(net9),
    .C(net37),
    .D(net36),
    .X(_00425_));
 sky130_fd_sc_hd__a22oi_1 _06599_ (.A1(net9),
    .A2(net37),
    .B1(net36),
    .B2(net10),
    .Y(_00426_));
 sky130_fd_sc_hd__and4bb_1 _06600_ (.A_N(_00425_),
    .B_N(_00426_),
    .C(net8),
    .D(net38),
    .X(_00427_));
 sky130_fd_sc_hd__nor2_1 _06601_ (.A(_00425_),
    .B(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__o2bb2a_1 _06602_ (.A1_N(net41),
    .A2_N(net6),
    .B1(_00348_),
    .B2(_00349_),
    .X(_00429_));
 sky130_fd_sc_hd__nor2_1 _06603_ (.A(_00351_),
    .B(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__o21a_1 _06604_ (.A1(_00425_),
    .A2(_00427_),
    .B1(_00430_),
    .X(_00431_));
 sky130_fd_sc_hd__and4_1 _06605_ (.A(net40),
    .B(net39),
    .C(net7),
    .D(net6),
    .X(_00432_));
 sky130_fd_sc_hd__a22oi_1 _06606_ (.A1(net39),
    .A2(net7),
    .B1(net6),
    .B2(net40),
    .Y(_00433_));
 sky130_fd_sc_hd__a22o_1 _06607_ (.A1(net39),
    .A2(net7),
    .B1(net6),
    .B2(net40),
    .X(_00434_));
 sky130_fd_sc_hd__and4b_1 _06608_ (.A_N(_00432_),
    .B(_00434_),
    .C(net41),
    .D(net5),
    .X(_00435_));
 sky130_fd_sc_hd__a31o_1 _06609_ (.A1(_00434_),
    .A2(net5),
    .A3(net41),
    .B1(_00432_),
    .X(_00436_));
 sky130_fd_sc_hd__xnor2_1 _06610_ (.A(_00428_),
    .B(_00430_),
    .Y(_00437_));
 sky130_fd_sc_hd__o21a_1 _06611_ (.A1(_00432_),
    .A2(_00435_),
    .B1(_00437_),
    .X(_00438_));
 sky130_fd_sc_hd__a21o_1 _06612_ (.A1(_00437_),
    .A2(_00436_),
    .B1(_00431_),
    .X(_00439_));
 sky130_fd_sc_hd__nor2_1 _06613_ (.A(_00352_),
    .B(_00354_),
    .Y(_00440_));
 sky130_fd_sc_hd__nor2_1 _06614_ (.A(_00355_),
    .B(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__o21a_1 _06615_ (.A1(_00431_),
    .A2(_00438_),
    .B1(_00441_),
    .X(_00442_));
 sky130_fd_sc_hd__and4_1 _06616_ (.A(net43),
    .B(net42),
    .C(net5),
    .D(net4),
    .X(_00443_));
 sky130_fd_sc_hd__nand4_2 _06617_ (.A(net43),
    .B(net42),
    .C(net5),
    .D(net4),
    .Y(_00444_));
 sky130_fd_sc_hd__a22oi_1 _06618_ (.A1(net42),
    .A2(net5),
    .B1(net4),
    .B2(net43),
    .Y(_00445_));
 sky130_fd_sc_hd__and4b_1 _06619_ (.A_N(_00445_),
    .B(net3),
    .C(net45),
    .D(_00444_),
    .X(_00446_));
 sky130_fd_sc_hd__or4_1 _06620_ (.A(_01054_),
    .B(_00445_),
    .C(_01120_),
    .D(_00443_),
    .X(_00447_));
 sky130_fd_sc_hd__o2bb2a_1 _06621_ (.A1_N(net45),
    .A2_N(net4),
    .B1(_00359_),
    .B2(_00361_),
    .X(_00448_));
 sky130_fd_sc_hd__o211a_1 _06622_ (.A1(_00362_),
    .A2(_00448_),
    .B1(_00447_),
    .C1(_00444_),
    .X(_00449_));
 sky130_fd_sc_hd__a211oi_2 _06623_ (.A1(_00444_),
    .A2(_00447_),
    .B1(_00448_),
    .C1(_00362_),
    .Y(_00450_));
 sky130_fd_sc_hd__nor2_1 _06624_ (.A(_00449_),
    .B(_00450_),
    .Y(_00451_));
 sky130_fd_sc_hd__and4_1 _06625_ (.A(net46),
    .B(net47),
    .C(net3),
    .D(net2),
    .X(_00452_));
 sky130_fd_sc_hd__o2bb2a_1 _06626_ (.A1_N(net46),
    .A2_N(net3),
    .B1(_01131_),
    .B2(_01043_),
    .X(_00453_));
 sky130_fd_sc_hd__nor2_1 _06627_ (.A(_00452_),
    .B(_00453_),
    .Y(_00454_));
 sky130_fd_sc_hd__and2_1 _06628_ (.A(net32),
    .B(_00454_),
    .X(_00455_));
 sky130_fd_sc_hd__nor2_1 _06629_ (.A(net32),
    .B(_00454_),
    .Y(_00456_));
 sky130_fd_sc_hd__or2_1 _06630_ (.A(_00455_),
    .B(_00456_),
    .X(_00457_));
 sky130_fd_sc_hd__nor3_1 _06631_ (.A(_00449_),
    .B(_00450_),
    .C(_00457_),
    .Y(_00458_));
 sky130_fd_sc_hd__xor2_1 _06632_ (.A(_00451_),
    .B(_00457_),
    .X(_00459_));
 sky130_fd_sc_hd__nor2_1 _06633_ (.A(_00439_),
    .B(_00441_),
    .Y(_00460_));
 sky130_fd_sc_hd__or2_1 _06634_ (.A(_00442_),
    .B(_00460_),
    .X(_00461_));
 sky130_fd_sc_hd__nor2_1 _06635_ (.A(_00459_),
    .B(_00461_),
    .Y(_00462_));
 sky130_fd_sc_hd__and3_1 _06636_ (.A(net15),
    .B(net63),
    .C(net62),
    .X(_00463_));
 sky130_fd_sc_hd__nor2_1 _06637_ (.A(_00385_),
    .B(_00388_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_1 _06638_ (.A(_00389_),
    .B(_00464_),
    .Y(_00465_));
 sky130_fd_sc_hd__and4_1 _06639_ (.A(net14),
    .B(net13),
    .C(net34),
    .D(net64),
    .X(_00466_));
 sky130_fd_sc_hd__a22oi_1 _06640_ (.A1(net13),
    .A2(net34),
    .B1(net64),
    .B2(net14),
    .Y(_00467_));
 sky130_fd_sc_hd__and4bb_1 _06641_ (.A_N(_00466_),
    .B_N(_00467_),
    .C(net11),
    .D(net35),
    .X(_00468_));
 sky130_fd_sc_hd__o2bb2a_1 _06642_ (.A1_N(net13),
    .A2_N(net35),
    .B1(_00378_),
    .B2(_00379_),
    .X(_00469_));
 sky130_fd_sc_hd__nor2_1 _06643_ (.A(_00380_),
    .B(_00469_),
    .Y(_00470_));
 sky130_fd_sc_hd__o21a_1 _06644_ (.A1(_00466_),
    .A2(_00468_),
    .B1(_00470_),
    .X(_00471_));
 sky130_fd_sc_hd__a2bb2o_1 _06645_ (.A1_N(_00342_),
    .A2_N(_00344_),
    .B1(net9),
    .B2(net38),
    .X(_00472_));
 sky130_fd_sc_hd__nand2_1 _06646_ (.A(_00345_),
    .B(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor3_1 _06647_ (.A(_00466_),
    .B(_00468_),
    .C(_00470_),
    .Y(_00474_));
 sky130_fd_sc_hd__or2_1 _06648_ (.A(_00471_),
    .B(_00474_),
    .X(_00475_));
 sky130_fd_sc_hd__nor2_1 _06649_ (.A(_00473_),
    .B(_00475_),
    .Y(_00476_));
 sky130_fd_sc_hd__xor2_1 _06650_ (.A(_00463_),
    .B(_00465_),
    .X(_00477_));
 sky130_fd_sc_hd__o21a_1 _06651_ (.A1(_00471_),
    .A2(_00476_),
    .B1(_00477_),
    .X(_00478_));
 sky130_fd_sc_hd__a41o_1 _06652_ (.A1(net15),
    .A2(net63),
    .A3(net62),
    .A4(_00465_),
    .B1(_00478_),
    .X(_00479_));
 sky130_fd_sc_hd__nand2_1 _06653_ (.A(_00374_),
    .B(_00376_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_1 _06654_ (.A(_00377_),
    .B(_00480_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2b_1 _06655_ (.A_N(_00481_),
    .B(_00479_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2b_1 _06656_ (.A_N(_00479_),
    .B(_00481_),
    .Y(_00483_));
 sky130_fd_sc_hd__a221o_1 _06657_ (.A1(_00441_),
    .A2(_00439_),
    .B1(_00483_),
    .B2(_00482_),
    .C1(_00462_),
    .X(_00484_));
 sky130_fd_sc_hd__o211ai_1 _06658_ (.A1(_00442_),
    .A2(_00462_),
    .B1(_00482_),
    .C1(_00483_),
    .Y(_00485_));
 sky130_fd_sc_hd__and2_1 _06659_ (.A(_00484_),
    .B(_00485_),
    .X(_00486_));
 sky130_fd_sc_hd__a311o_1 _06660_ (.A1(_00304_),
    .A2(_00381_),
    .A3(_00382_),
    .B1(_00389_),
    .C1(_00392_),
    .X(_00487_));
 sky130_fd_sc_hd__and2_1 _06661_ (.A(_00393_),
    .B(_00487_),
    .X(_00488_));
 sky130_fd_sc_hd__nand2_1 _06662_ (.A(_00486_),
    .B(_00488_),
    .Y(_00489_));
 sky130_fd_sc_hd__xnor2_1 _06663_ (.A(_00401_),
    .B(_00403_),
    .Y(_00490_));
 sky130_fd_sc_hd__or2_1 _06664_ (.A(_00489_),
    .B(_00490_),
    .X(_00491_));
 sky130_fd_sc_hd__nand2_1 _06665_ (.A(_00489_),
    .B(_00490_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _06666_ (.A(_00491_),
    .B(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__and4bb_1 _06667_ (.A_N(_00366_),
    .B_N(_00373_),
    .C(_00482_),
    .D(_00485_),
    .X(_00494_));
 sky130_fd_sc_hd__a2bb2oi_1 _06668_ (.A1_N(_00366_),
    .A2_N(_00373_),
    .B1(_00482_),
    .B2(_00485_),
    .Y(_00495_));
 sky130_fd_sc_hd__nor2_1 _06669_ (.A(_00494_),
    .B(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__o21a_1 _06670_ (.A1(_00368_),
    .A2(_00370_),
    .B1(_00496_),
    .X(_00497_));
 sky130_fd_sc_hd__nor3_1 _06671_ (.A(_00368_),
    .B(_00370_),
    .C(_00496_),
    .Y(_00498_));
 sky130_fd_sc_hd__or3_1 _06672_ (.A(_00497_),
    .B(_00498_),
    .C(_00493_),
    .X(_00499_));
 sky130_fd_sc_hd__xnor2_1 _06673_ (.A(_00407_),
    .B(_00415_),
    .Y(_00500_));
 sky130_fd_sc_hd__a21oi_1 _06674_ (.A1(_00491_),
    .A2(_00499_),
    .B1(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__a21o_1 _06675_ (.A1(_00491_),
    .A2(_00499_),
    .B1(_00500_),
    .X(_00502_));
 sky130_fd_sc_hd__nor2_1 _06676_ (.A(_00495_),
    .B(_00497_),
    .Y(_00503_));
 sky130_fd_sc_hd__o311a_1 _06677_ (.A1(_00493_),
    .A2(_00497_),
    .A3(_00498_),
    .B1(_00500_),
    .C1(_00491_),
    .X(_00504_));
 sky130_fd_sc_hd__nor2_1 _06678_ (.A(_00501_),
    .B(_00504_),
    .Y(_00505_));
 sky130_fd_sc_hd__o21ai_1 _06679_ (.A1(_00503_),
    .A2(_00504_),
    .B1(_00502_),
    .Y(_00506_));
 sky130_fd_sc_hd__o211ai_1 _06680_ (.A1(_00411_),
    .A2(_00408_),
    .B1(_00410_),
    .C1(_00420_),
    .Y(_00507_));
 sky130_fd_sc_hd__and2_1 _06681_ (.A(_00421_),
    .B(_00507_),
    .X(_00508_));
 sky130_fd_sc_hd__xnor2_1 _06682_ (.A(_00506_),
    .B(_00508_),
    .Y(_00509_));
 sky130_fd_sc_hd__nor3_1 _06683_ (.A(_00471_),
    .B(_00476_),
    .C(_00477_),
    .Y(_00510_));
 sky130_fd_sc_hd__or2_1 _06684_ (.A(_00478_),
    .B(_00510_),
    .X(_00511_));
 sky130_fd_sc_hd__a21o_1 _06685_ (.A1(net15),
    .A2(net62),
    .B1(_01142_),
    .X(_00512_));
 sky130_fd_sc_hd__and4_1 _06686_ (.A(net13),
    .B(net11),
    .C(net34),
    .D(net64),
    .X(_00513_));
 sky130_fd_sc_hd__a22oi_1 _06687_ (.A1(net11),
    .A2(net34),
    .B1(net64),
    .B2(net13),
    .Y(_00514_));
 sky130_fd_sc_hd__and4bb_1 _06688_ (.A_N(_00513_),
    .B_N(_00514_),
    .C(net10),
    .D(net35),
    .X(_00515_));
 sky130_fd_sc_hd__a41o_1 _06689_ (.A1(net13),
    .A2(net11),
    .A3(net34),
    .A4(net64),
    .B1(_00515_),
    .X(_00516_));
 sky130_fd_sc_hd__o2bb2a_1 _06690_ (.A1_N(net11),
    .A2_N(net35),
    .B1(_00466_),
    .B2(_00467_),
    .X(_00517_));
 sky130_fd_sc_hd__nor2_1 _06691_ (.A(_00468_),
    .B(_00517_),
    .Y(_00518_));
 sky130_fd_sc_hd__o2bb2a_1 _06692_ (.A1_N(net8),
    .A2_N(net38),
    .B1(_00425_),
    .B2(_00426_),
    .X(_00519_));
 sky130_fd_sc_hd__xnor2_1 _06693_ (.A(_00516_),
    .B(_00518_),
    .Y(_00520_));
 sky130_fd_sc_hd__nor3_1 _06694_ (.A(_00427_),
    .B(_00519_),
    .C(_00520_),
    .Y(_00521_));
 sky130_fd_sc_hd__a21o_1 _06695_ (.A1(_00516_),
    .A2(_00518_),
    .B1(_00521_),
    .X(_00522_));
 sky130_fd_sc_hd__a21oi_1 _06696_ (.A1(net15),
    .A2(net63),
    .B1(net62),
    .Y(_00523_));
 sky130_fd_sc_hd__and3_1 _06697_ (.A(net15),
    .B(net62),
    .C(net61),
    .X(_00524_));
 sky130_fd_sc_hd__or3b_2 _06698_ (.A(_01032_),
    .B(_01164_),
    .C_N(net61),
    .X(_00525_));
 sky130_fd_sc_hd__a21oi_1 _06699_ (.A1(net15),
    .A2(net62),
    .B1(net61),
    .Y(_00526_));
 sky130_fd_sc_hd__or4bb_2 _06700_ (.A(_00524_),
    .B(_00526_),
    .C_N(net14),
    .D_N(net63),
    .X(_00527_));
 sky130_fd_sc_hd__a211oi_2 _06701_ (.A1(_00525_),
    .A2(_00527_),
    .B1(_00463_),
    .C1(_00523_),
    .Y(_00528_));
 sky130_fd_sc_hd__and2_1 _06702_ (.A(_00473_),
    .B(_00475_),
    .X(_00529_));
 sky130_fd_sc_hd__nor2_1 _06703_ (.A(_00476_),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__or3b_1 _06704_ (.A(_00476_),
    .B(_00529_),
    .C_N(_00528_),
    .X(_00531_));
 sky130_fd_sc_hd__xor2_1 _06705_ (.A(_00528_),
    .B(_00530_),
    .X(_00532_));
 sky130_fd_sc_hd__nand2_1 _06706_ (.A(_00532_),
    .B(_00522_),
    .Y(_00533_));
 sky130_fd_sc_hd__a211o_1 _06707_ (.A1(_00516_),
    .A2(_00518_),
    .B1(_00521_),
    .C1(_00532_),
    .X(_00534_));
 sky130_fd_sc_hd__nand2_1 _06708_ (.A(_00533_),
    .B(_00534_),
    .Y(_00535_));
 sky130_fd_sc_hd__or3_2 _06709_ (.A(_00511_),
    .B(_00512_),
    .C(_00535_),
    .X(_00536_));
 sky130_fd_sc_hd__and4_1 _06710_ (.A(net9),
    .B(net8),
    .C(net37),
    .D(net36),
    .X(_00537_));
 sky130_fd_sc_hd__a22oi_1 _06711_ (.A1(net8),
    .A2(net37),
    .B1(net36),
    .B2(net9),
    .Y(_00538_));
 sky130_fd_sc_hd__and4bb_1 _06712_ (.A_N(_00537_),
    .B_N(_00538_),
    .C(net7),
    .D(net38),
    .X(_00539_));
 sky130_fd_sc_hd__nor2_1 _06713_ (.A(_00537_),
    .B(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__o2bb2a_1 _06714_ (.A1_N(net41),
    .A2_N(net5),
    .B1(_00432_),
    .B2(_00433_),
    .X(_00541_));
 sky130_fd_sc_hd__nor2_1 _06715_ (.A(_00435_),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__o21a_1 _06716_ (.A1(_00537_),
    .A2(_00539_),
    .B1(_00542_),
    .X(_00543_));
 sky130_fd_sc_hd__and4_1 _06717_ (.A(net40),
    .B(net39),
    .C(net6),
    .D(net5),
    .X(_00544_));
 sky130_fd_sc_hd__a22oi_1 _06718_ (.A1(net39),
    .A2(net6),
    .B1(net5),
    .B2(net40),
    .Y(_00545_));
 sky130_fd_sc_hd__a22o_1 _06719_ (.A1(net39),
    .A2(net6),
    .B1(net5),
    .B2(net40),
    .X(_00546_));
 sky130_fd_sc_hd__and4b_1 _06720_ (.A_N(_00544_),
    .B(_00546_),
    .C(net41),
    .D(net4),
    .X(_00547_));
 sky130_fd_sc_hd__a31o_1 _06721_ (.A1(_00546_),
    .A2(net4),
    .A3(net41),
    .B1(_00544_),
    .X(_00548_));
 sky130_fd_sc_hd__xnor2_1 _06722_ (.A(_00540_),
    .B(_00542_),
    .Y(_00549_));
 sky130_fd_sc_hd__o21a_1 _06723_ (.A1(_00544_),
    .A2(_00547_),
    .B1(_00549_),
    .X(_00550_));
 sky130_fd_sc_hd__nor2_1 _06724_ (.A(_00436_),
    .B(_00437_),
    .Y(_00551_));
 sky130_fd_sc_hd__nor2_1 _06725_ (.A(_00438_),
    .B(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__o21ai_1 _06726_ (.A1(_00543_),
    .A2(_00550_),
    .B1(_00552_),
    .Y(_00553_));
 sky130_fd_sc_hd__and4_1 _06727_ (.A(net43),
    .B(net42),
    .C(net4),
    .D(net3),
    .X(_00554_));
 sky130_fd_sc_hd__nand4_2 _06728_ (.A(net43),
    .B(net42),
    .C(net4),
    .D(net3),
    .Y(_00555_));
 sky130_fd_sc_hd__o2bb2a_1 _06729_ (.A1_N(net42),
    .A2_N(net4),
    .B1(_01120_),
    .B2(_01065_),
    .X(_00556_));
 sky130_fd_sc_hd__and4b_1 _06730_ (.A_N(_00556_),
    .B(net2),
    .C(net45),
    .D(_00555_),
    .X(_00557_));
 sky130_fd_sc_hd__or4_1 _06731_ (.A(_01054_),
    .B(_01131_),
    .C(_00554_),
    .D(_00556_),
    .X(_00558_));
 sky130_fd_sc_hd__o22a_1 _06732_ (.A1(_01054_),
    .A2(_01120_),
    .B1(_00443_),
    .B2(_00445_),
    .X(_00559_));
 sky130_fd_sc_hd__o211a_1 _06733_ (.A1(_00446_),
    .A2(_00559_),
    .B1(_00558_),
    .C1(_00555_),
    .X(_00560_));
 sky130_fd_sc_hd__a211oi_2 _06734_ (.A1(_00555_),
    .A2(_00558_),
    .B1(_00559_),
    .C1(_00446_),
    .Y(_00561_));
 sky130_fd_sc_hd__nor2_1 _06735_ (.A(_00560_),
    .B(_00561_),
    .Y(_00562_));
 sky130_fd_sc_hd__and4_1 _06736_ (.A(net46),
    .B(net47),
    .C(net2),
    .D(net32),
    .X(_00563_));
 sky130_fd_sc_hd__a22oi_1 _06737_ (.A1(net46),
    .A2(net2),
    .B1(net32),
    .B2(net47),
    .Y(_00564_));
 sky130_fd_sc_hd__nor2_1 _06738_ (.A(_00563_),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__xor2_1 _06739_ (.A(_01153_),
    .B(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__nor3_1 _06740_ (.A(_00560_),
    .B(_00566_),
    .C(_00561_),
    .Y(_00567_));
 sky130_fd_sc_hd__xor2_1 _06741_ (.A(_00562_),
    .B(_00566_),
    .X(_00568_));
 sky130_fd_sc_hd__or3_1 _06742_ (.A(_00543_),
    .B(_00550_),
    .C(_00552_),
    .X(_00569_));
 sky130_fd_sc_hd__nand2_1 _06743_ (.A(_00553_),
    .B(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__o21a_1 _06744_ (.A1(_00568_),
    .A2(_00570_),
    .B1(_00553_),
    .X(_00571_));
 sky130_fd_sc_hd__and2_1 _06745_ (.A(_00459_),
    .B(_00461_),
    .X(_00572_));
 sky130_fd_sc_hd__or2_1 _06746_ (.A(_00462_),
    .B(_00572_),
    .X(_00573_));
 sky130_fd_sc_hd__nand3_1 _06747_ (.A(_00531_),
    .B(_00533_),
    .C(_00573_),
    .Y(_00574_));
 sky130_fd_sc_hd__a21o_1 _06748_ (.A1(_00531_),
    .A2(_00533_),
    .B1(_00573_),
    .X(_00575_));
 sky130_fd_sc_hd__nand2_1 _06749_ (.A(_00574_),
    .B(_00575_),
    .Y(_00576_));
 sky130_fd_sc_hd__or2_1 _06750_ (.A(_00571_),
    .B(_00576_),
    .X(_00577_));
 sky130_fd_sc_hd__nand2_1 _06751_ (.A(_00576_),
    .B(_00571_),
    .Y(_00578_));
 sky130_fd_sc_hd__o21ai_1 _06752_ (.A1(_00512_),
    .A2(_00535_),
    .B1(_00511_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand4_2 _06753_ (.A(_00536_),
    .B(_00577_),
    .C(_00578_),
    .D(_00579_),
    .Y(_00580_));
 sky130_fd_sc_hd__or2_1 _06754_ (.A(_00486_),
    .B(_00488_),
    .X(_00581_));
 sky130_fd_sc_hd__nand2_1 _06755_ (.A(_00489_),
    .B(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__a21oi_2 _06756_ (.A1(_00536_),
    .A2(_00580_),
    .B1(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__inv_2 _06757_ (.A(_00583_),
    .Y(_00584_));
 sky130_fd_sc_hd__o311a_1 _06758_ (.A1(_00511_),
    .A2(_00512_),
    .A3(_00535_),
    .B1(_00580_),
    .C1(_00582_),
    .X(_00585_));
 sky130_fd_sc_hd__and4bb_1 _06759_ (.A_N(_00450_),
    .B_N(_00458_),
    .C(_00575_),
    .D(_00577_),
    .X(_00586_));
 sky130_fd_sc_hd__a2bb2oi_1 _06760_ (.A1_N(_00450_),
    .A2_N(_00458_),
    .B1(_00575_),
    .B2(_00577_),
    .Y(_00587_));
 sky130_fd_sc_hd__nor2_1 _06761_ (.A(_00586_),
    .B(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__o21a_1 _06762_ (.A1(_00452_),
    .A2(_00455_),
    .B1(_00588_),
    .X(_00589_));
 sky130_fd_sc_hd__a211oi_1 _06763_ (.A1(net32),
    .A2(_00454_),
    .B1(_00588_),
    .C1(_00452_),
    .Y(_00590_));
 sky130_fd_sc_hd__or4_1 _06764_ (.A(_00583_),
    .B(_00585_),
    .C(_00589_),
    .D(_00590_),
    .X(_00591_));
 sky130_fd_sc_hd__o21ai_1 _06765_ (.A1(_00497_),
    .A2(_00498_),
    .B1(_00493_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _06766_ (.A(_00499_),
    .B(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__a21oi_1 _06767_ (.A1(_00584_),
    .A2(_00591_),
    .B1(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__o311a_1 _06768_ (.A1(_00585_),
    .A2(_00589_),
    .A3(_00590_),
    .B1(_00593_),
    .C1(_00584_),
    .X(_00595_));
 sky130_fd_sc_hd__nor2_1 _06769_ (.A(_00594_),
    .B(_00595_),
    .Y(_00596_));
 sky130_fd_sc_hd__o21a_1 _06770_ (.A1(_00587_),
    .A2(_00589_),
    .B1(_00596_),
    .X(_00597_));
 sky130_fd_sc_hd__xnor2_1 _06771_ (.A(_00503_),
    .B(_00505_),
    .Y(_00598_));
 sky130_fd_sc_hd__o21ai_1 _06772_ (.A1(_00594_),
    .A2(_00597_),
    .B1(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__or3_1 _06773_ (.A(_00594_),
    .B(_00597_),
    .C(_00598_),
    .X(_00600_));
 sky130_fd_sc_hd__and2_1 _06774_ (.A(_00599_),
    .B(_00600_),
    .X(_00601_));
 sky130_fd_sc_hd__o211a_1 _06775_ (.A1(_00463_),
    .A2(_00523_),
    .B1(_00525_),
    .C1(_00527_),
    .X(_00602_));
 sky130_fd_sc_hd__and4_1 _06776_ (.A(net11),
    .B(net10),
    .C(net34),
    .D(net64),
    .X(_00603_));
 sky130_fd_sc_hd__a22oi_1 _06777_ (.A1(net10),
    .A2(net34),
    .B1(net64),
    .B2(net11),
    .Y(_00604_));
 sky130_fd_sc_hd__nor4_1 _06778_ (.A(_01076_),
    .B(_00604_),
    .C(_01109_),
    .D(_00603_),
    .Y(_00605_));
 sky130_fd_sc_hd__nor2_1 _06779_ (.A(_00603_),
    .B(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__o2bb2a_1 _06780_ (.A1_N(net10),
    .A2_N(net35),
    .B1(_00513_),
    .B2(_00514_),
    .X(_00607_));
 sky130_fd_sc_hd__nor2_1 _06781_ (.A(_00515_),
    .B(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__or3_1 _06782_ (.A(_00515_),
    .B(_00606_),
    .C(_00607_),
    .X(_00609_));
 sky130_fd_sc_hd__o2bb2a_1 _06783_ (.A1_N(net7),
    .A2_N(net38),
    .B1(_00537_),
    .B2(_00538_),
    .X(_00610_));
 sky130_fd_sc_hd__xor2_1 _06784_ (.A(_00606_),
    .B(_00608_),
    .X(_00611_));
 sky130_fd_sc_hd__or3_1 _06785_ (.A(_00539_),
    .B(_00610_),
    .C(_00611_),
    .X(_00612_));
 sky130_fd_sc_hd__and4_1 _06786_ (.A(net15),
    .B(net14),
    .C(net62),
    .D(net61),
    .X(_00613_));
 sky130_fd_sc_hd__a22oi_1 _06787_ (.A1(net14),
    .A2(net62),
    .B1(net61),
    .B2(net15),
    .Y(_00614_));
 sky130_fd_sc_hd__and4bb_1 _06788_ (.A_N(_00613_),
    .B_N(_00614_),
    .C(net13),
    .D(net63),
    .X(_00615_));
 sky130_fd_sc_hd__a2bb2o_1 _06789_ (.A1_N(_00524_),
    .A2_N(_00526_),
    .B1(net14),
    .B2(net63),
    .X(_00616_));
 sky130_fd_sc_hd__o211ai_2 _06790_ (.A1(_00613_),
    .A2(_00615_),
    .B1(_00616_),
    .C1(_00527_),
    .Y(_00617_));
 sky130_fd_sc_hd__o21a_1 _06791_ (.A1(_00427_),
    .A2(_00519_),
    .B1(_00520_),
    .X(_00618_));
 sky130_fd_sc_hd__o21a_1 _06792_ (.A1(_00521_),
    .A2(_00618_),
    .B1(_00617_),
    .X(_00619_));
 sky130_fd_sc_hd__nor3_1 _06793_ (.A(_00617_),
    .B(_00618_),
    .C(_00521_),
    .Y(_00620_));
 sky130_fd_sc_hd__a211oi_2 _06794_ (.A1(_00609_),
    .A2(_00612_),
    .B1(_00619_),
    .C1(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hd__o211ai_1 _06795_ (.A1(_00619_),
    .A2(_00620_),
    .B1(_00609_),
    .C1(_00612_),
    .Y(_00622_));
 sky130_fd_sc_hd__inv_2 _06796_ (.A(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__or4_1 _06797_ (.A(_00528_),
    .B(_00602_),
    .C(_00621_),
    .D(_00623_),
    .X(_00624_));
 sky130_fd_sc_hd__inv_2 _06798_ (.A(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__xor2_1 _06799_ (.A(_00512_),
    .B(_00535_),
    .X(_00626_));
 sky130_fd_sc_hd__xor2_1 _06800_ (.A(_00624_),
    .B(_00626_),
    .X(_00627_));
 sky130_fd_sc_hd__and4_1 _06801_ (.A(net8),
    .B(net7),
    .C(net37),
    .D(net36),
    .X(_00628_));
 sky130_fd_sc_hd__a22oi_1 _06802_ (.A1(net7),
    .A2(net37),
    .B1(net36),
    .B2(net8),
    .Y(_00629_));
 sky130_fd_sc_hd__and4bb_1 _06803_ (.A_N(_00628_),
    .B_N(_00629_),
    .C(net38),
    .D(net6),
    .X(_00630_));
 sky130_fd_sc_hd__nor2_1 _06804_ (.A(_00628_),
    .B(_00630_),
    .Y(_00631_));
 sky130_fd_sc_hd__o2bb2a_1 _06805_ (.A1_N(net41),
    .A2_N(net4),
    .B1(_00544_),
    .B2(_00545_),
    .X(_00632_));
 sky130_fd_sc_hd__nor2_1 _06806_ (.A(_00547_),
    .B(_00632_),
    .Y(_00633_));
 sky130_fd_sc_hd__o21a_1 _06807_ (.A1(_00628_),
    .A2(_00630_),
    .B1(_00633_),
    .X(_00634_));
 sky130_fd_sc_hd__and4_1 _06808_ (.A(net40),
    .B(net39),
    .C(net5),
    .D(net4),
    .X(_00635_));
 sky130_fd_sc_hd__a22oi_1 _06809_ (.A1(net39),
    .A2(net5),
    .B1(net4),
    .B2(net40),
    .Y(_00636_));
 sky130_fd_sc_hd__a22o_1 _06810_ (.A1(net39),
    .A2(net5),
    .B1(net4),
    .B2(net40),
    .X(_00637_));
 sky130_fd_sc_hd__and4b_1 _06811_ (.A_N(_00635_),
    .B(_00637_),
    .C(net41),
    .D(net3),
    .X(_00638_));
 sky130_fd_sc_hd__a31o_1 _06812_ (.A1(_00637_),
    .A2(net3),
    .A3(net41),
    .B1(_00635_),
    .X(_00639_));
 sky130_fd_sc_hd__xnor2_1 _06813_ (.A(_00631_),
    .B(_00633_),
    .Y(_00640_));
 sky130_fd_sc_hd__o21a_1 _06814_ (.A1(_00635_),
    .A2(_00638_),
    .B1(_00640_),
    .X(_00641_));
 sky130_fd_sc_hd__nor2_1 _06815_ (.A(_00548_),
    .B(_00549_),
    .Y(_00642_));
 sky130_fd_sc_hd__nor2_1 _06816_ (.A(_00550_),
    .B(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hd__o21ai_1 _06817_ (.A1(_00634_),
    .A2(_00641_),
    .B1(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__and4_1 _06818_ (.A(net43),
    .B(net42),
    .C(net3),
    .D(net2),
    .X(_00645_));
 sky130_fd_sc_hd__nand4_2 _06819_ (.A(net43),
    .B(net42),
    .C(net3),
    .D(net2),
    .Y(_00646_));
 sky130_fd_sc_hd__o2bb2a_1 _06820_ (.A1_N(net42),
    .A2_N(net3),
    .B1(_01131_),
    .B2(_01065_),
    .X(_00647_));
 sky130_fd_sc_hd__and4b_1 _06821_ (.A_N(_00647_),
    .B(net32),
    .C(net45),
    .D(_00646_),
    .X(_00648_));
 sky130_fd_sc_hd__or4b_1 _06822_ (.A(_01054_),
    .B(_00645_),
    .C(_00647_),
    .D_N(net32),
    .X(_00649_));
 sky130_fd_sc_hd__o22a_1 _06823_ (.A1(_01054_),
    .A2(_01131_),
    .B1(_00554_),
    .B2(_00556_),
    .X(_00650_));
 sky130_fd_sc_hd__o211a_1 _06824_ (.A1(_00557_),
    .A2(_00650_),
    .B1(_00649_),
    .C1(_00646_),
    .X(_00651_));
 sky130_fd_sc_hd__a211oi_2 _06825_ (.A1(_00646_),
    .A2(_00649_),
    .B1(_00650_),
    .C1(_00557_),
    .Y(_00652_));
 sky130_fd_sc_hd__nor2_1 _06826_ (.A(_00651_),
    .B(_00652_),
    .Y(_00653_));
 sky130_fd_sc_hd__and4_1 _06827_ (.A(net46),
    .B(net47),
    .C(net32),
    .D(net31),
    .X(_00654_));
 sky130_fd_sc_hd__o2bb2a_1 _06828_ (.A1_N(net46),
    .A2_N(net32),
    .B1(_01153_),
    .B2(_01043_),
    .X(_00655_));
 sky130_fd_sc_hd__nor3_1 _06829_ (.A(_01175_),
    .B(_00654_),
    .C(_00655_),
    .Y(_00656_));
 sky130_fd_sc_hd__o21ai_1 _06830_ (.A1(_00654_),
    .A2(_00655_),
    .B1(_01175_),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2b_1 _06831_ (.A_N(_00656_),
    .B(_00657_),
    .Y(_00658_));
 sky130_fd_sc_hd__nor3_1 _06832_ (.A(_00651_),
    .B(_00658_),
    .C(_00652_),
    .Y(_00659_));
 sky130_fd_sc_hd__xor2_1 _06833_ (.A(_00653_),
    .B(_00658_),
    .X(_00660_));
 sky130_fd_sc_hd__or3_1 _06834_ (.A(_00634_),
    .B(_00641_),
    .C(_00643_),
    .X(_00661_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_00644_),
    .B(_00661_),
    .Y(_00662_));
 sky130_fd_sc_hd__o21a_1 _06836_ (.A1(_00660_),
    .A2(_00662_),
    .B1(_00644_),
    .X(_00663_));
 sky130_fd_sc_hd__xor2_1 _06837_ (.A(_00568_),
    .B(_00570_),
    .X(_00664_));
 sky130_fd_sc_hd__or3_1 _06838_ (.A(_00620_),
    .B(_00621_),
    .C(_00664_),
    .X(_00665_));
 sky130_fd_sc_hd__o21ai_1 _06839_ (.A1(_00620_),
    .A2(_00621_),
    .B1(_00664_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(_00665_),
    .B(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__or2_1 _06841_ (.A(_00663_),
    .B(_00667_),
    .X(_00668_));
 sky130_fd_sc_hd__nand2_1 _06842_ (.A(_00667_),
    .B(_00663_),
    .Y(_00669_));
 sky130_fd_sc_hd__and2_1 _06843_ (.A(_00668_),
    .B(_00669_),
    .X(_00670_));
 sky130_fd_sc_hd__and2b_1 _06844_ (.A_N(_00627_),
    .B(_00670_),
    .X(_00671_));
 sky130_fd_sc_hd__a21oi_1 _06845_ (.A1(_00625_),
    .A2(_00626_),
    .B1(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__a22o_1 _06846_ (.A1(_00577_),
    .A2(_00578_),
    .B1(_00579_),
    .B2(_00536_),
    .X(_00673_));
 sky130_fd_sc_hd__nand2_1 _06847_ (.A(_00580_),
    .B(_00673_),
    .Y(_00674_));
 sky130_fd_sc_hd__nor2_1 _06848_ (.A(_00674_),
    .B(_00672_),
    .Y(_00675_));
 sky130_fd_sc_hd__xnor2_1 _06849_ (.A(_00672_),
    .B(_00674_),
    .Y(_00676_));
 sky130_fd_sc_hd__a21o_1 _06850_ (.A1(net31),
    .A2(_00565_),
    .B1(_00563_),
    .X(_00677_));
 sky130_fd_sc_hd__and4bb_1 _06851_ (.A_N(_00561_),
    .B_N(_00567_),
    .C(_00666_),
    .D(_00668_),
    .X(_00678_));
 sky130_fd_sc_hd__a2bb2oi_1 _06852_ (.A1_N(_00561_),
    .A2_N(_00567_),
    .B1(_00666_),
    .B2(_00668_),
    .Y(_00679_));
 sky130_fd_sc_hd__nor2_1 _06853_ (.A(_00678_),
    .B(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__xnor2_1 _06854_ (.A(_00677_),
    .B(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__nor2_1 _06855_ (.A(_00676_),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__o22ai_1 _06856_ (.A1(_00583_),
    .A2(_00585_),
    .B1(_00589_),
    .B2(_00590_),
    .Y(_00683_));
 sky130_fd_sc_hd__o211a_1 _06857_ (.A1(_00675_),
    .A2(_00682_),
    .B1(_00683_),
    .C1(_00591_),
    .X(_00684_));
 sky130_fd_sc_hd__a21oi_1 _06858_ (.A1(_00680_),
    .A2(_00677_),
    .B1(_00679_),
    .Y(_00685_));
 sky130_fd_sc_hd__a211oi_1 _06859_ (.A1(_00591_),
    .A2(_00683_),
    .B1(_00682_),
    .C1(_00675_),
    .Y(_00686_));
 sky130_fd_sc_hd__nor3_1 _06860_ (.A(_00684_),
    .B(_00685_),
    .C(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__nor3_1 _06861_ (.A(_00587_),
    .B(_00589_),
    .C(_00596_),
    .Y(_00688_));
 sky130_fd_sc_hd__or2_1 _06862_ (.A(_00597_),
    .B(_00688_),
    .X(_00689_));
 sky130_fd_sc_hd__o21bai_1 _06863_ (.A1(_00684_),
    .A2(_00687_),
    .B1_N(_00689_),
    .Y(_00690_));
 sky130_fd_sc_hd__or3b_1 _06864_ (.A(_00684_),
    .B(_00687_),
    .C_N(_00689_),
    .X(_00691_));
 sky130_fd_sc_hd__nand2_1 _06865_ (.A(_00690_),
    .B(_00691_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(_00676_),
    .B(_00681_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2b_1 _06867_ (.A_N(_00682_),
    .B(_00693_),
    .Y(_00694_));
 sky130_fd_sc_hd__a211o_1 _06868_ (.A1(_00527_),
    .A2(_00616_),
    .B1(_00615_),
    .C1(_00613_),
    .X(_00695_));
 sky130_fd_sc_hd__nand2_1 _06869_ (.A(_00617_),
    .B(_00695_),
    .Y(_00696_));
 sky130_fd_sc_hd__and4_1 _06870_ (.A(net14),
    .B(net13),
    .C(net62),
    .D(net61),
    .X(_00697_));
 sky130_fd_sc_hd__a22oi_1 _06871_ (.A1(net13),
    .A2(net62),
    .B1(net61),
    .B2(net14),
    .Y(_00698_));
 sky130_fd_sc_hd__and4bb_1 _06872_ (.A_N(_00697_),
    .B_N(_00698_),
    .C(net11),
    .D(net63),
    .X(_00699_));
 sky130_fd_sc_hd__and3_1 _06873_ (.A(net15),
    .B(net60),
    .C(net59),
    .X(_00700_));
 sky130_fd_sc_hd__o2bb2a_1 _06874_ (.A1_N(net13),
    .A2_N(net63),
    .B1(_00613_),
    .B2(_00614_),
    .X(_00701_));
 sky130_fd_sc_hd__or3b_1 _06875_ (.A(_00615_),
    .B(_00701_),
    .C_N(_00700_),
    .X(_00702_));
 sky130_fd_sc_hd__o21bai_1 _06876_ (.A1(_00615_),
    .A2(_00701_),
    .B1_N(_00700_),
    .Y(_00703_));
 sky130_fd_sc_hd__and2_1 _06877_ (.A(_00702_),
    .B(_00703_),
    .X(_00704_));
 sky130_fd_sc_hd__o21ai_1 _06878_ (.A1(_00697_),
    .A2(_00699_),
    .B1(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__or3_1 _06879_ (.A(_00697_),
    .B(_00699_),
    .C(_00704_),
    .X(_00706_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(_00705_),
    .B(_00706_),
    .Y(_00707_));
 sky130_fd_sc_hd__or2_1 _06881_ (.A(_01197_),
    .B(_00707_),
    .X(_00708_));
 sky130_fd_sc_hd__or3_1 _06882_ (.A(_01197_),
    .B(_00696_),
    .C(_00707_),
    .X(_00709_));
 sky130_fd_sc_hd__and4_1 _06883_ (.A(net10),
    .B(net9),
    .C(net34),
    .D(net64),
    .X(_00710_));
 sky130_fd_sc_hd__a22oi_1 _06884_ (.A1(net9),
    .A2(net34),
    .B1(net64),
    .B2(net10),
    .Y(_00711_));
 sky130_fd_sc_hd__and4bb_1 _06885_ (.A_N(_00710_),
    .B_N(_00711_),
    .C(net8),
    .D(net35),
    .X(_00712_));
 sky130_fd_sc_hd__a41o_1 _06886_ (.A1(net10),
    .A2(net9),
    .A3(net34),
    .A4(net64),
    .B1(_00712_),
    .X(_00713_));
 sky130_fd_sc_hd__o22a_1 _06887_ (.A1(_01076_),
    .A2(_01109_),
    .B1(_00603_),
    .B2(_00604_),
    .X(_00714_));
 sky130_fd_sc_hd__nor2_1 _06888_ (.A(_00605_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__o2bb2a_1 _06889_ (.A1_N(net38),
    .A2_N(net6),
    .B1(_00628_),
    .B2(_00629_),
    .X(_00716_));
 sky130_fd_sc_hd__xnor2_1 _06890_ (.A(_00713_),
    .B(_00715_),
    .Y(_00717_));
 sky130_fd_sc_hd__nor3_1 _06891_ (.A(_00630_),
    .B(_00716_),
    .C(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__a21o_1 _06892_ (.A1(_00713_),
    .A2(_00715_),
    .B1(_00718_),
    .X(_00719_));
 sky130_fd_sc_hd__o21ai_1 _06893_ (.A1(_00539_),
    .A2(_00610_),
    .B1(_00611_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand2_1 _06894_ (.A(_00612_),
    .B(_00720_),
    .Y(_00721_));
 sky130_fd_sc_hd__and3_1 _06895_ (.A(_00702_),
    .B(_00705_),
    .C(_00721_),
    .X(_00722_));
 sky130_fd_sc_hd__a21o_1 _06896_ (.A1(_00702_),
    .A2(_00705_),
    .B1(_00721_),
    .X(_00723_));
 sky130_fd_sc_hd__and2b_1 _06897_ (.A_N(_00722_),
    .B(_00723_),
    .X(_00724_));
 sky130_fd_sc_hd__nand2_1 _06898_ (.A(_00724_),
    .B(_00719_),
    .Y(_00725_));
 sky130_fd_sc_hd__a211o_1 _06899_ (.A1(_00713_),
    .A2(_00715_),
    .B1(_00718_),
    .C1(_00724_),
    .X(_00726_));
 sky130_fd_sc_hd__nand2_1 _06900_ (.A(_00725_),
    .B(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__a2bb2o_1 _06901_ (.A1_N(_01197_),
    .A2_N(_00707_),
    .B1(_00695_),
    .B2(_00617_),
    .X(_00728_));
 sky130_fd_sc_hd__nand2_1 _06902_ (.A(_00709_),
    .B(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__or2_1 _06903_ (.A(_00727_),
    .B(_00729_),
    .X(_00730_));
 sky130_fd_sc_hd__o22a_1 _06904_ (.A1(_00528_),
    .A2(_00602_),
    .B1(_00621_),
    .B2(_00623_),
    .X(_00731_));
 sky130_fd_sc_hd__a211oi_1 _06905_ (.A1(_00709_),
    .A2(_00730_),
    .B1(_00731_),
    .C1(_00625_),
    .Y(_00732_));
 sky130_fd_sc_hd__and4_1 _06906_ (.A(net7),
    .B(net6),
    .C(net37),
    .D(net36),
    .X(_00733_));
 sky130_fd_sc_hd__nand4_1 _06907_ (.A(net7),
    .B(net6),
    .C(net37),
    .D(net36),
    .Y(_00734_));
 sky130_fd_sc_hd__a22oi_1 _06908_ (.A1(net6),
    .A2(net37),
    .B1(net36),
    .B2(net7),
    .Y(_00735_));
 sky130_fd_sc_hd__or4_1 _06909_ (.A(_01087_),
    .B(_00735_),
    .C(_01098_),
    .D(_00733_),
    .X(_00736_));
 sky130_fd_sc_hd__o2bb2a_1 _06910_ (.A1_N(net41),
    .A2_N(net3),
    .B1(_00635_),
    .B2(_00636_),
    .X(_00737_));
 sky130_fd_sc_hd__a211oi_1 _06911_ (.A1(_00734_),
    .A2(_00736_),
    .B1(_00737_),
    .C1(_00638_),
    .Y(_00738_));
 sky130_fd_sc_hd__and4_1 _06912_ (.A(net40),
    .B(net39),
    .C(net4),
    .D(net3),
    .X(_00739_));
 sky130_fd_sc_hd__a22oi_1 _06913_ (.A1(net39),
    .A2(net4),
    .B1(net3),
    .B2(net40),
    .Y(_00740_));
 sky130_fd_sc_hd__a22o_1 _06914_ (.A1(net39),
    .A2(net4),
    .B1(net3),
    .B2(net40),
    .X(_00741_));
 sky130_fd_sc_hd__and4b_1 _06915_ (.A_N(_00739_),
    .B(_00741_),
    .C(net41),
    .D(net2),
    .X(_00742_));
 sky130_fd_sc_hd__a31o_1 _06916_ (.A1(_00741_),
    .A2(net2),
    .A3(net41),
    .B1(_00739_),
    .X(_00743_));
 sky130_fd_sc_hd__o211a_1 _06917_ (.A1(_00638_),
    .A2(_00737_),
    .B1(_00736_),
    .C1(_00734_),
    .X(_00744_));
 sky130_fd_sc_hd__nor2_1 _06918_ (.A(_00738_),
    .B(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__o21a_1 _06919_ (.A1(_00739_),
    .A2(_00742_),
    .B1(_00745_),
    .X(_00746_));
 sky130_fd_sc_hd__nor2_1 _06920_ (.A(_00639_),
    .B(_00640_),
    .Y(_00747_));
 sky130_fd_sc_hd__nor2_1 _06921_ (.A(_00641_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__o21ai_1 _06922_ (.A1(_00738_),
    .A2(_00746_),
    .B1(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__and4_1 _06923_ (.A(net43),
    .B(net42),
    .C(net2),
    .D(net32),
    .X(_00750_));
 sky130_fd_sc_hd__nand4_2 _06924_ (.A(net43),
    .B(net42),
    .C(net2),
    .D(net32),
    .Y(_00751_));
 sky130_fd_sc_hd__a22oi_1 _06925_ (.A1(net42),
    .A2(net2),
    .B1(net32),
    .B2(net43),
    .Y(_00752_));
 sky130_fd_sc_hd__and4b_1 _06926_ (.A_N(_00752_),
    .B(net31),
    .C(net45),
    .D(_00751_),
    .X(_00753_));
 sky130_fd_sc_hd__or4_1 _06927_ (.A(_01054_),
    .B(_00752_),
    .C(_01153_),
    .D(_00750_),
    .X(_00754_));
 sky130_fd_sc_hd__o2bb2a_1 _06928_ (.A1_N(net45),
    .A2_N(net32),
    .B1(_00645_),
    .B2(_00647_),
    .X(_00755_));
 sky130_fd_sc_hd__o211a_1 _06929_ (.A1(_00648_),
    .A2(_00755_),
    .B1(_00754_),
    .C1(_00751_),
    .X(_00756_));
 sky130_fd_sc_hd__a211oi_2 _06930_ (.A1(_00751_),
    .A2(_00754_),
    .B1(_00755_),
    .C1(_00648_),
    .Y(_00757_));
 sky130_fd_sc_hd__nor2_1 _06931_ (.A(_00756_),
    .B(_00757_),
    .Y(_00758_));
 sky130_fd_sc_hd__and4_1 _06932_ (.A(net46),
    .B(net47),
    .C(net31),
    .D(net30),
    .X(_00759_));
 sky130_fd_sc_hd__o2bb2a_1 _06933_ (.A1_N(net46),
    .A2_N(net31),
    .B1(_01175_),
    .B2(_01043_),
    .X(_00760_));
 sky130_fd_sc_hd__nor2_1 _06934_ (.A(_00759_),
    .B(_00760_),
    .Y(_00761_));
 sky130_fd_sc_hd__xor2_1 _06935_ (.A(_01186_),
    .B(_00761_),
    .X(_00762_));
 sky130_fd_sc_hd__nor3_1 _06936_ (.A(_00762_),
    .B(_00757_),
    .C(_00756_),
    .Y(_00763_));
 sky130_fd_sc_hd__xor2_1 _06937_ (.A(_00758_),
    .B(_00762_),
    .X(_00764_));
 sky130_fd_sc_hd__or3_1 _06938_ (.A(_00738_),
    .B(_00746_),
    .C(_00748_),
    .X(_00765_));
 sky130_fd_sc_hd__nand2_1 _06939_ (.A(_00749_),
    .B(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hd__o21a_1 _06940_ (.A1(_00764_),
    .A2(_00766_),
    .B1(_00749_),
    .X(_00767_));
 sky130_fd_sc_hd__xnor2_1 _06941_ (.A(_00660_),
    .B(_00662_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand3_1 _06942_ (.A(_00723_),
    .B(_00725_),
    .C(_00768_),
    .Y(_00769_));
 sky130_fd_sc_hd__a21o_1 _06943_ (.A1(_00723_),
    .A2(_00725_),
    .B1(_00768_),
    .X(_00770_));
 sky130_fd_sc_hd__nand2_1 _06944_ (.A(_00769_),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__or2_1 _06945_ (.A(_00767_),
    .B(_00771_),
    .X(_00772_));
 sky130_fd_sc_hd__nand2_1 _06946_ (.A(_00771_),
    .B(_00767_),
    .Y(_00773_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(_00772_),
    .B(_00773_),
    .Y(_00774_));
 sky130_fd_sc_hd__o221a_1 _06948_ (.A1(_00696_),
    .A2(_00708_),
    .B1(_00731_),
    .B2(_00625_),
    .C1(_00730_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _06949_ (.A(_00732_),
    .B(_00775_),
    .X(_00776_));
 sky130_fd_sc_hd__nor2_1 _06950_ (.A(_00774_),
    .B(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__xnor2_1 _06951_ (.A(_00627_),
    .B(_00670_),
    .Y(_00778_));
 sky130_fd_sc_hd__o21ai_1 _06952_ (.A1(_00732_),
    .A2(_00777_),
    .B1(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hd__or3_1 _06953_ (.A(_00732_),
    .B(_00777_),
    .C(_00778_),
    .X(_00780_));
 sky130_fd_sc_hd__nand2_1 _06954_ (.A(_00779_),
    .B(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hd__and4bb_1 _06955_ (.A_N(_00652_),
    .B_N(_00659_),
    .C(_00770_),
    .D(_00772_),
    .X(_00782_));
 sky130_fd_sc_hd__a2bb2oi_1 _06956_ (.A1_N(_00652_),
    .A2_N(_00659_),
    .B1(_00770_),
    .B2(_00772_),
    .Y(_00783_));
 sky130_fd_sc_hd__nor2_1 _06957_ (.A(_00782_),
    .B(_00783_),
    .Y(_00784_));
 sky130_fd_sc_hd__o21a_1 _06958_ (.A1(_00654_),
    .A2(_00656_),
    .B1(_00784_),
    .X(_00785_));
 sky130_fd_sc_hd__nor3_1 _06959_ (.A(_00654_),
    .B(_00656_),
    .C(_00784_),
    .Y(_00786_));
 sky130_fd_sc_hd__or3_1 _06960_ (.A(_00785_),
    .B(_00786_),
    .C(_00781_),
    .X(_00787_));
 sky130_fd_sc_hd__a21oi_1 _06961_ (.A1(_00779_),
    .A2(_00787_),
    .B1(_00694_),
    .Y(_00788_));
 sky130_fd_sc_hd__or2_1 _06962_ (.A(_00783_),
    .B(_00785_),
    .X(_00789_));
 sky130_fd_sc_hd__o311a_1 _06963_ (.A1(_00781_),
    .A2(_00785_),
    .A3(_00786_),
    .B1(_00779_),
    .C1(_00694_),
    .X(_00790_));
 sky130_fd_sc_hd__nor2_1 _06964_ (.A(_00788_),
    .B(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__a21o_1 _06965_ (.A1(_00791_),
    .A2(_00789_),
    .B1(_00788_),
    .X(_00792_));
 sky130_fd_sc_hd__o21a_1 _06966_ (.A1(_00684_),
    .A2(_00686_),
    .B1(_00685_),
    .X(_00793_));
 sky130_fd_sc_hd__nor2_1 _06967_ (.A(_00687_),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__o21ai_1 _06968_ (.A1(_00785_),
    .A2(_00786_),
    .B1(_00781_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand2_1 _06969_ (.A(_00787_),
    .B(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand2_1 _06970_ (.A(_00727_),
    .B(_00729_),
    .Y(_00797_));
 sky130_fd_sc_hd__and2_1 _06971_ (.A(_00730_),
    .B(_00797_),
    .X(_00798_));
 sky130_fd_sc_hd__and4_1 _06972_ (.A(net13),
    .B(net11),
    .C(net62),
    .D(net61),
    .X(_00799_));
 sky130_fd_sc_hd__a22oi_1 _06973_ (.A1(net11),
    .A2(net62),
    .B1(net61),
    .B2(net13),
    .Y(_00800_));
 sky130_fd_sc_hd__and4bb_1 _06974_ (.A_N(_00799_),
    .B_N(_00800_),
    .C(net10),
    .D(net63),
    .X(_00801_));
 sky130_fd_sc_hd__nand3_1 _06975_ (.A(net15),
    .B(net59),
    .C(net58),
    .Y(_00802_));
 sky130_fd_sc_hd__a21o_1 _06976_ (.A1(net15),
    .A2(net59),
    .B1(net58),
    .X(_00803_));
 sky130_fd_sc_hd__nand4_1 _06977_ (.A(_00803_),
    .B(net60),
    .C(net14),
    .D(_00802_),
    .Y(_00804_));
 sky130_fd_sc_hd__o2bb2a_1 _06978_ (.A1_N(net11),
    .A2_N(net63),
    .B1(_00697_),
    .B2(_00698_),
    .X(_00805_));
 sky130_fd_sc_hd__a211o_1 _06979_ (.A1(_00802_),
    .A2(_00804_),
    .B1(_00805_),
    .C1(_00699_),
    .X(_00806_));
 sky130_fd_sc_hd__o211ai_1 _06980_ (.A1(_00699_),
    .A2(_00805_),
    .B1(_00804_),
    .C1(_00802_),
    .Y(_00807_));
 sky130_fd_sc_hd__and2_1 _06981_ (.A(_00806_),
    .B(_00807_),
    .X(_00808_));
 sky130_fd_sc_hd__o21ai_1 _06982_ (.A1(_00799_),
    .A2(_00801_),
    .B1(_00808_),
    .Y(_00809_));
 sky130_fd_sc_hd__or3_1 _06983_ (.A(_00799_),
    .B(_00801_),
    .C(_00808_),
    .X(_00810_));
 sky130_fd_sc_hd__nand2_1 _06984_ (.A(_00809_),
    .B(_00810_),
    .Y(_00811_));
 sky130_fd_sc_hd__a21oi_1 _06985_ (.A1(net15),
    .A2(net60),
    .B1(net59),
    .Y(_00812_));
 sky130_fd_sc_hd__or3_1 _06986_ (.A(_00700_),
    .B(_00812_),
    .C(_00811_),
    .X(_00813_));
 sky130_fd_sc_hd__nand2_1 _06987_ (.A(_01197_),
    .B(_00707_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _06988_ (.A(_00708_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__nor2_1 _06989_ (.A(_00813_),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__and4_1 _06990_ (.A(net9),
    .B(net8),
    .C(net34),
    .D(net64),
    .X(_00817_));
 sky130_fd_sc_hd__a22oi_1 _06991_ (.A1(net8),
    .A2(net34),
    .B1(net64),
    .B2(net9),
    .Y(_00818_));
 sky130_fd_sc_hd__a22o_1 _06992_ (.A1(net8),
    .A2(net34),
    .B1(net64),
    .B2(net9),
    .X(_00819_));
 sky130_fd_sc_hd__and4b_1 _06993_ (.A_N(_00817_),
    .B(_00819_),
    .C(net7),
    .D(net35),
    .X(_00820_));
 sky130_fd_sc_hd__a31o_1 _06994_ (.A1(_00819_),
    .A2(net35),
    .A3(net7),
    .B1(_00817_),
    .X(_00821_));
 sky130_fd_sc_hd__o2bb2a_1 _06995_ (.A1_N(net8),
    .A2_N(net35),
    .B1(_00710_),
    .B2(_00711_),
    .X(_00822_));
 sky130_fd_sc_hd__nor2_1 _06996_ (.A(_00712_),
    .B(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__a2bb2o_1 _06997_ (.A1_N(_00733_),
    .A2_N(_00735_),
    .B1(net38),
    .B2(net5),
    .X(_00824_));
 sky130_fd_sc_hd__nand2_1 _06998_ (.A(_00736_),
    .B(_00824_),
    .Y(_00825_));
 sky130_fd_sc_hd__xnor2_1 _06999_ (.A(_00821_),
    .B(_00823_),
    .Y(_00826_));
 sky130_fd_sc_hd__nor2_1 _07000_ (.A(_00825_),
    .B(_00826_),
    .Y(_00827_));
 sky130_fd_sc_hd__a21o_1 _07001_ (.A1(_00821_),
    .A2(_00823_),
    .B1(_00827_),
    .X(_00828_));
 sky130_fd_sc_hd__o21a_1 _07002_ (.A1(_00630_),
    .A2(_00716_),
    .B1(_00717_),
    .X(_00829_));
 sky130_fd_sc_hd__o211a_1 _07003_ (.A1(_00718_),
    .A2(_00829_),
    .B1(_00809_),
    .C1(_00806_),
    .X(_00830_));
 sky130_fd_sc_hd__a211oi_1 _07004_ (.A1(_00806_),
    .A2(_00809_),
    .B1(_00829_),
    .C1(_00718_),
    .Y(_00831_));
 sky130_fd_sc_hd__nor2_1 _07005_ (.A(_00830_),
    .B(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__xor2_1 _07006_ (.A(_00828_),
    .B(_00832_),
    .X(_00833_));
 sky130_fd_sc_hd__o31a_1 _07007_ (.A1(_00700_),
    .A2(_00811_),
    .A3(_00812_),
    .B1(_00815_),
    .X(_00834_));
 sky130_fd_sc_hd__nor2_1 _07008_ (.A(_00816_),
    .B(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__and2_1 _07009_ (.A(_00833_),
    .B(_00835_),
    .X(_00836_));
 sky130_fd_sc_hd__o21a_1 _07010_ (.A1(_00816_),
    .A2(_00836_),
    .B1(_00798_),
    .X(_00837_));
 sky130_fd_sc_hd__and4_1 _07011_ (.A(net6),
    .B(net37),
    .C(net5),
    .D(net36),
    .X(_00838_));
 sky130_fd_sc_hd__nand4_1 _07012_ (.A(net6),
    .B(net37),
    .C(net5),
    .D(net36),
    .Y(_00839_));
 sky130_fd_sc_hd__a22oi_1 _07013_ (.A1(net37),
    .A2(net5),
    .B1(net36),
    .B2(net6),
    .Y(_00840_));
 sky130_fd_sc_hd__or4b_1 _07014_ (.A(_00840_),
    .B(_01087_),
    .C(_00838_),
    .D_N(net4),
    .X(_00841_));
 sky130_fd_sc_hd__o2bb2a_1 _07015_ (.A1_N(net41),
    .A2_N(net2),
    .B1(_00739_),
    .B2(_00740_),
    .X(_00842_));
 sky130_fd_sc_hd__a211oi_1 _07016_ (.A1(_00839_),
    .A2(_00841_),
    .B1(_00842_),
    .C1(_00742_),
    .Y(_00843_));
 sky130_fd_sc_hd__and4_1 _07017_ (.A(net40),
    .B(net39),
    .C(net3),
    .D(net2),
    .X(_00844_));
 sky130_fd_sc_hd__a22oi_1 _07018_ (.A1(net39),
    .A2(net3),
    .B1(net2),
    .B2(net40),
    .Y(_00845_));
 sky130_fd_sc_hd__a22o_1 _07019_ (.A1(net39),
    .A2(net3),
    .B1(net2),
    .B2(net40),
    .X(_00846_));
 sky130_fd_sc_hd__and4b_1 _07020_ (.A_N(_00844_),
    .B(_00846_),
    .C(net41),
    .D(net32),
    .X(_00847_));
 sky130_fd_sc_hd__a31o_1 _07021_ (.A1(_00846_),
    .A2(net32),
    .A3(net41),
    .B1(_00844_),
    .X(_00848_));
 sky130_fd_sc_hd__o211a_1 _07022_ (.A1(_00742_),
    .A2(_00842_),
    .B1(_00841_),
    .C1(_00839_),
    .X(_00849_));
 sky130_fd_sc_hd__nor2_1 _07023_ (.A(_00843_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__o21a_1 _07024_ (.A1(_00844_),
    .A2(_00847_),
    .B1(_00850_),
    .X(_00851_));
 sky130_fd_sc_hd__nor2_1 _07025_ (.A(_00743_),
    .B(_00745_),
    .Y(_00852_));
 sky130_fd_sc_hd__nor2_1 _07026_ (.A(_00746_),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__o21ai_1 _07027_ (.A1(_00843_),
    .A2(_00851_),
    .B1(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__and4_1 _07028_ (.A(net43),
    .B(net42),
    .C(net32),
    .D(net31),
    .X(_00855_));
 sky130_fd_sc_hd__nand4_2 _07029_ (.A(net43),
    .B(net42),
    .C(net32),
    .D(net31),
    .Y(_00856_));
 sky130_fd_sc_hd__o2bb2a_1 _07030_ (.A1_N(net42),
    .A2_N(net32),
    .B1(_01153_),
    .B2(_01065_),
    .X(_00857_));
 sky130_fd_sc_hd__and4b_1 _07031_ (.A_N(_00857_),
    .B(net30),
    .C(net45),
    .D(_00856_),
    .X(_00858_));
 sky130_fd_sc_hd__or4_1 _07032_ (.A(_01054_),
    .B(_01175_),
    .C(_00855_),
    .D(_00857_),
    .X(_00859_));
 sky130_fd_sc_hd__o22a_1 _07033_ (.A1(_01054_),
    .A2(_01153_),
    .B1(_00750_),
    .B2(_00752_),
    .X(_00860_));
 sky130_fd_sc_hd__o211a_1 _07034_ (.A1(_00753_),
    .A2(_00860_),
    .B1(_00859_),
    .C1(_00856_),
    .X(_00861_));
 sky130_fd_sc_hd__a211oi_2 _07035_ (.A1(_00856_),
    .A2(_00859_),
    .B1(_00860_),
    .C1(_00753_),
    .Y(_00862_));
 sky130_fd_sc_hd__nor2_1 _07036_ (.A(_00861_),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__and4_1 _07037_ (.A(net46),
    .B(net47),
    .C(net30),
    .D(net29),
    .X(_00864_));
 sky130_fd_sc_hd__o2bb2a_1 _07038_ (.A1_N(net46),
    .A2_N(net30),
    .B1(_01186_),
    .B2(_01043_),
    .X(_00865_));
 sky130_fd_sc_hd__nor2_1 _07039_ (.A(_00864_),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__and2_1 _07040_ (.A(net28),
    .B(_00866_),
    .X(_00867_));
 sky130_fd_sc_hd__nor2_1 _07041_ (.A(net28),
    .B(_00866_),
    .Y(_00868_));
 sky130_fd_sc_hd__or2_1 _07042_ (.A(_00867_),
    .B(_00868_),
    .X(_00869_));
 sky130_fd_sc_hd__nor3_1 _07043_ (.A(_00861_),
    .B(_00869_),
    .C(_00862_),
    .Y(_00870_));
 sky130_fd_sc_hd__xor2_1 _07044_ (.A(_00863_),
    .B(_00869_),
    .X(_00871_));
 sky130_fd_sc_hd__or3_1 _07045_ (.A(_00843_),
    .B(_00851_),
    .C(_00853_),
    .X(_00872_));
 sky130_fd_sc_hd__nand2_1 _07046_ (.A(_00854_),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__or2_1 _07047_ (.A(_00871_),
    .B(_00873_),
    .X(_00874_));
 sky130_fd_sc_hd__a21oi_1 _07048_ (.A1(_00832_),
    .A2(_00828_),
    .B1(_00831_),
    .Y(_00875_));
 sky130_fd_sc_hd__xnor2_1 _07049_ (.A(_00764_),
    .B(_00766_),
    .Y(_00876_));
 sky130_fd_sc_hd__or2_1 _07050_ (.A(_00875_),
    .B(_00876_),
    .X(_00877_));
 sky130_fd_sc_hd__xnor2_1 _07051_ (.A(_00875_),
    .B(_00876_),
    .Y(_00878_));
 sky130_fd_sc_hd__a21o_1 _07052_ (.A1(_00854_),
    .A2(_00874_),
    .B1(_00878_),
    .X(_00879_));
 sky130_fd_sc_hd__o211ai_1 _07053_ (.A1(_00871_),
    .A2(_00873_),
    .B1(_00878_),
    .C1(_00854_),
    .Y(_00880_));
 sky130_fd_sc_hd__and2_1 _07054_ (.A(_00879_),
    .B(_00880_),
    .X(_00881_));
 sky130_fd_sc_hd__a211oi_1 _07055_ (.A1(_00833_),
    .A2(_00835_),
    .B1(_00798_),
    .C1(_00816_),
    .Y(_00882_));
 sky130_fd_sc_hd__nor2_1 _07056_ (.A(_00837_),
    .B(_00882_),
    .Y(_00883_));
 sky130_fd_sc_hd__and2_1 _07057_ (.A(_00881_),
    .B(_00883_),
    .X(_00884_));
 sky130_fd_sc_hd__a21o_1 _07058_ (.A1(_00881_),
    .A2(_00883_),
    .B1(_00837_),
    .X(_00885_));
 sky130_fd_sc_hd__and2_1 _07059_ (.A(_00774_),
    .B(_00776_),
    .X(_00886_));
 sky130_fd_sc_hd__nor2_1 _07060_ (.A(_00777_),
    .B(_00886_),
    .Y(_00887_));
 sky130_fd_sc_hd__xnor2_1 _07061_ (.A(_00885_),
    .B(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__a21o_1 _07062_ (.A1(net29),
    .A2(_00761_),
    .B1(_00759_),
    .X(_00889_));
 sky130_fd_sc_hd__and4bb_1 _07063_ (.A_N(_00757_),
    .B_N(_00763_),
    .C(_00877_),
    .D(_00879_),
    .X(_00890_));
 sky130_fd_sc_hd__a2bb2oi_1 _07064_ (.A1_N(_00757_),
    .A2_N(_00763_),
    .B1(_00877_),
    .B2(_00879_),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2_1 _07065_ (.A(_00890_),
    .B(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__xnor2_1 _07066_ (.A(_00889_),
    .B(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__nor2_1 _07067_ (.A(_00888_),
    .B(_00893_),
    .Y(_00894_));
 sky130_fd_sc_hd__a21o_1 _07068_ (.A1(_00885_),
    .A2(_00887_),
    .B1(_00894_),
    .X(_00895_));
 sky130_fd_sc_hd__nand2b_1 _07069_ (.A_N(_00796_),
    .B(_00895_),
    .Y(_00896_));
 sky130_fd_sc_hd__xnor2_1 _07070_ (.A(_00796_),
    .B(_00895_),
    .Y(_00897_));
 sky130_fd_sc_hd__a21oi_1 _07071_ (.A1(_00892_),
    .A2(_00889_),
    .B1(_00891_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand2b_1 _07072_ (.A_N(_00898_),
    .B(_00897_),
    .Y(_00899_));
 sky130_fd_sc_hd__xnor2_1 _07073_ (.A(_00789_),
    .B(_00791_),
    .Y(_00900_));
 sky130_fd_sc_hd__a21oi_1 _07074_ (.A1(_00896_),
    .A2(_00899_),
    .B1(_00900_),
    .Y(_00901_));
 sky130_fd_sc_hd__and3_1 _07075_ (.A(_00896_),
    .B(_00899_),
    .C(_00900_),
    .X(_00902_));
 sky130_fd_sc_hd__nor2_1 _07076_ (.A(_00901_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__xnor2_1 _07077_ (.A(_00897_),
    .B(_00898_),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_1 _07078_ (.A(_00888_),
    .B(_00893_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2b_1 _07079_ (.A_N(_00894_),
    .B(_00905_),
    .Y(_00906_));
 sky130_fd_sc_hd__a22o_1 _07080_ (.A1(net14),
    .A2(net60),
    .B1(_00802_),
    .B2(_00803_),
    .X(_00907_));
 sky130_fd_sc_hd__and2_1 _07081_ (.A(_00804_),
    .B(_00907_),
    .X(_00908_));
 sky130_fd_sc_hd__nand2_2 _07082_ (.A(net15),
    .B(net44),
    .Y(_00909_));
 sky130_fd_sc_hd__nand4_2 _07083_ (.A(net15),
    .B(net14),
    .C(net59),
    .D(net58),
    .Y(_00910_));
 sky130_fd_sc_hd__a22o_1 _07084_ (.A1(net14),
    .A2(net59),
    .B1(net58),
    .B2(net15),
    .X(_00911_));
 sky130_fd_sc_hd__and4_1 _07085_ (.A(_00911_),
    .B(net60),
    .C(net13),
    .D(_00910_),
    .X(_00912_));
 sky130_fd_sc_hd__nand4_1 _07086_ (.A(_00911_),
    .B(net60),
    .C(net13),
    .D(_00910_),
    .Y(_00913_));
 sky130_fd_sc_hd__a22oi_1 _07087_ (.A1(net13),
    .A2(net60),
    .B1(_00910_),
    .B2(_00911_),
    .Y(_00914_));
 sky130_fd_sc_hd__a2111o_1 _07088_ (.A1(net15),
    .A2(net44),
    .B1(_01230_),
    .C1(_00914_),
    .D1(_00912_),
    .X(_00915_));
 sky130_fd_sc_hd__inv_2 _07089_ (.A(_00915_),
    .Y(_00916_));
 sky130_fd_sc_hd__a31o_1 _07090_ (.A1(net15),
    .A2(net55),
    .A3(net44),
    .B1(_00916_),
    .X(_00917_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(_00917_),
    .B(_00908_),
    .Y(_00918_));
 sky130_fd_sc_hd__and4_2 _07092_ (.A(net11),
    .B(net10),
    .C(net62),
    .D(net61),
    .X(_00919_));
 sky130_fd_sc_hd__a22oi_1 _07093_ (.A1(net10),
    .A2(net62),
    .B1(net61),
    .B2(net11),
    .Y(_00920_));
 sky130_fd_sc_hd__a22o_1 _07094_ (.A1(net10),
    .A2(net62),
    .B1(net61),
    .B2(net11),
    .X(_00921_));
 sky130_fd_sc_hd__and4b_1 _07095_ (.A_N(_00919_),
    .B(_00921_),
    .C(net9),
    .D(net63),
    .X(_00922_));
 sky130_fd_sc_hd__o2bb2a_1 _07096_ (.A1_N(net10),
    .A2_N(net63),
    .B1(_00799_),
    .B2(_00800_),
    .X(_00923_));
 sky130_fd_sc_hd__o211a_1 _07097_ (.A1(_00801_),
    .A2(_00923_),
    .B1(_00913_),
    .C1(_00910_),
    .X(_00924_));
 sky130_fd_sc_hd__a211o_1 _07098_ (.A1(_00910_),
    .A2(_00913_),
    .B1(_00923_),
    .C1(_00801_),
    .X(_00925_));
 sky130_fd_sc_hd__and2b_1 _07099_ (.A_N(_00924_),
    .B(_00925_),
    .X(_00926_));
 sky130_fd_sc_hd__o21ai_4 _07100_ (.A1(_00919_),
    .A2(_00922_),
    .B1(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__a311o_1 _07101_ (.A1(net9),
    .A2(_00921_),
    .A3(net63),
    .B1(_00919_),
    .C1(_00926_),
    .X(_00928_));
 sky130_fd_sc_hd__a311o_1 _07102_ (.A1(net15),
    .A2(net55),
    .A3(net44),
    .B1(_00908_),
    .C1(_00916_),
    .X(_00929_));
 sky130_fd_sc_hd__nand4_2 _07103_ (.A(_00918_),
    .B(_00927_),
    .C(_00928_),
    .D(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__o21ai_1 _07104_ (.A1(_00700_),
    .A2(_00812_),
    .B1(_00811_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _07105_ (.A(_00813_),
    .B(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__a21o_1 _07106_ (.A1(_00918_),
    .A2(_00930_),
    .B1(_00932_),
    .X(_00933_));
 sky130_fd_sc_hd__and4_1 _07107_ (.A(net8),
    .B(net7),
    .C(net34),
    .D(net64),
    .X(_00934_));
 sky130_fd_sc_hd__a22oi_1 _07108_ (.A1(net7),
    .A2(net34),
    .B1(net64),
    .B2(net8),
    .Y(_00935_));
 sky130_fd_sc_hd__a22o_1 _07109_ (.A1(net7),
    .A2(net34),
    .B1(net64),
    .B2(net8),
    .X(_00936_));
 sky130_fd_sc_hd__and4b_1 _07110_ (.A_N(_00934_),
    .B(_00936_),
    .C(net6),
    .D(net35),
    .X(_00937_));
 sky130_fd_sc_hd__o2bb2a_1 _07111_ (.A1_N(net7),
    .A2_N(net35),
    .B1(_00817_),
    .B2(_00818_),
    .X(_00938_));
 sky130_fd_sc_hd__nor2_1 _07112_ (.A(_00820_),
    .B(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__o21ai_1 _07113_ (.A1(_00934_),
    .A2(_00937_),
    .B1(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__a2bb2o_1 _07114_ (.A1_N(_00838_),
    .A2_N(_00840_),
    .B1(net38),
    .B2(net4),
    .X(_00941_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(_00841_),
    .B(_00941_),
    .Y(_00942_));
 sky130_fd_sc_hd__a311o_1 _07116_ (.A1(net6),
    .A2(_00936_),
    .A3(net35),
    .B1(_00934_),
    .C1(_00939_),
    .X(_00943_));
 sky130_fd_sc_hd__nand2_1 _07117_ (.A(_00940_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__nor2_1 _07118_ (.A(_00942_),
    .B(_00944_),
    .Y(_00945_));
 sky130_fd_sc_hd__or2_1 _07119_ (.A(_00942_),
    .B(_00944_),
    .X(_00946_));
 sky130_fd_sc_hd__and2_1 _07120_ (.A(_00825_),
    .B(_00826_),
    .X(_00947_));
 sky130_fd_sc_hd__o211a_1 _07121_ (.A1(_00827_),
    .A2(_00947_),
    .B1(_00927_),
    .C1(_00925_),
    .X(_00948_));
 sky130_fd_sc_hd__a211oi_4 _07122_ (.A1(_00925_),
    .A2(_00927_),
    .B1(_00947_),
    .C1(_00827_),
    .Y(_00949_));
 sky130_fd_sc_hd__a211oi_2 _07123_ (.A1(_00940_),
    .A2(_00946_),
    .B1(_00948_),
    .C1(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__o221a_1 _07124_ (.A1(_00942_),
    .A2(_00944_),
    .B1(_00948_),
    .B2(_00949_),
    .C1(_00940_),
    .X(_00951_));
 sky130_fd_sc_hd__nor2_1 _07125_ (.A(_00950_),
    .B(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand3_1 _07126_ (.A(_00918_),
    .B(_00930_),
    .C(_00932_),
    .Y(_00953_));
 sky130_fd_sc_hd__and2_1 _07127_ (.A(_00933_),
    .B(_00953_),
    .X(_00954_));
 sky130_fd_sc_hd__nand2_2 _07128_ (.A(_00952_),
    .B(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__nor2_1 _07129_ (.A(_00833_),
    .B(_00835_),
    .Y(_00956_));
 sky130_fd_sc_hd__a211o_1 _07130_ (.A1(_00933_),
    .A2(_00955_),
    .B1(_00956_),
    .C1(_00836_),
    .X(_00957_));
 sky130_fd_sc_hd__and4_1 _07131_ (.A(net37),
    .B(net5),
    .C(net36),
    .D(net4),
    .X(_00958_));
 sky130_fd_sc_hd__nand4_1 _07132_ (.A(net37),
    .B(net5),
    .C(net36),
    .D(net4),
    .Y(_00959_));
 sky130_fd_sc_hd__a22oi_1 _07133_ (.A1(net5),
    .A2(net36),
    .B1(net4),
    .B2(net37),
    .Y(_00960_));
 sky130_fd_sc_hd__or4_2 _07134_ (.A(_01087_),
    .B(_00960_),
    .C(_01120_),
    .D(_00958_),
    .X(_00961_));
 sky130_fd_sc_hd__o2bb2a_1 _07135_ (.A1_N(net41),
    .A2_N(net32),
    .B1(_00844_),
    .B2(_00845_),
    .X(_00962_));
 sky130_fd_sc_hd__a211oi_2 _07136_ (.A1(_00959_),
    .A2(_00961_),
    .B1(_00962_),
    .C1(_00847_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand4_1 _07137_ (.A(net40),
    .B(net39),
    .C(net2),
    .D(net32),
    .Y(_00964_));
 sky130_fd_sc_hd__a22o_1 _07138_ (.A1(net39),
    .A2(net2),
    .B1(net32),
    .B2(net40),
    .X(_00965_));
 sky130_fd_sc_hd__and4_1 _07139_ (.A(_00965_),
    .B(net31),
    .C(net41),
    .D(_00964_),
    .X(_00967_));
 sky130_fd_sc_hd__a41o_1 _07140_ (.A1(net40),
    .A2(net39),
    .A3(net2),
    .A4(net32),
    .B1(_00967_),
    .X(_00968_));
 sky130_fd_sc_hd__o211a_1 _07141_ (.A1(_00847_),
    .A2(_00962_),
    .B1(_00961_),
    .C1(_00959_),
    .X(_00969_));
 sky130_fd_sc_hd__nor2_1 _07142_ (.A(_00963_),
    .B(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__and2_1 _07143_ (.A(_00970_),
    .B(_00968_),
    .X(_00971_));
 sky130_fd_sc_hd__nor2_1 _07144_ (.A(_00848_),
    .B(_00850_),
    .Y(_00972_));
 sky130_fd_sc_hd__nor2_1 _07145_ (.A(_00851_),
    .B(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__o21a_1 _07146_ (.A1(_00963_),
    .A2(_00971_),
    .B1(_00973_),
    .X(_00974_));
 sky130_fd_sc_hd__o21ai_2 _07147_ (.A1(_00963_),
    .A2(_00971_),
    .B1(_00973_),
    .Y(_00975_));
 sky130_fd_sc_hd__and4_1 _07148_ (.A(net43),
    .B(net42),
    .C(net31),
    .D(net30),
    .X(_00976_));
 sky130_fd_sc_hd__nand4_2 _07149_ (.A(net43),
    .B(net42),
    .C(net31),
    .D(net30),
    .Y(_00978_));
 sky130_fd_sc_hd__o2bb2a_1 _07150_ (.A1_N(net42),
    .A2_N(net31),
    .B1(_01175_),
    .B2(_01065_),
    .X(_00979_));
 sky130_fd_sc_hd__and4b_1 _07151_ (.A_N(_00979_),
    .B(net29),
    .C(net45),
    .D(_00978_),
    .X(_00980_));
 sky130_fd_sc_hd__or4_1 _07152_ (.A(_01054_),
    .B(_01186_),
    .C(_00976_),
    .D(_00979_),
    .X(_00981_));
 sky130_fd_sc_hd__o22a_1 _07153_ (.A1(_01054_),
    .A2(_01175_),
    .B1(_00855_),
    .B2(_00857_),
    .X(_00982_));
 sky130_fd_sc_hd__o211a_1 _07154_ (.A1(_00858_),
    .A2(_00982_),
    .B1(_00981_),
    .C1(_00978_),
    .X(_00983_));
 sky130_fd_sc_hd__a211oi_2 _07155_ (.A1(_00978_),
    .A2(_00981_),
    .B1(_00982_),
    .C1(_00858_),
    .Y(_00984_));
 sky130_fd_sc_hd__and4_1 _07156_ (.A(net46),
    .B(net47),
    .C(net29),
    .D(net28),
    .X(_00985_));
 sky130_fd_sc_hd__a22oi_1 _07157_ (.A1(net46),
    .A2(net29),
    .B1(net28),
    .B2(net47),
    .Y(_00986_));
 sky130_fd_sc_hd__nor3_1 _07158_ (.A(_00986_),
    .B(_01208_),
    .C(_00985_),
    .Y(_00987_));
 sky130_fd_sc_hd__o21ai_1 _07159_ (.A1(_00985_),
    .A2(_00986_),
    .B1(_01208_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2b_1 _07160_ (.A_N(_00987_),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__o21a_1 _07161_ (.A1(_00983_),
    .A2(_00984_),
    .B1(_00990_),
    .X(_00991_));
 sky130_fd_sc_hd__nor3_1 _07162_ (.A(_00983_),
    .B(_00990_),
    .C(_00984_),
    .Y(_00992_));
 sky130_fd_sc_hd__or2_1 _07163_ (.A(_00991_),
    .B(_00992_),
    .X(_00993_));
 sky130_fd_sc_hd__a211oi_1 _07164_ (.A1(_00970_),
    .A2(_00968_),
    .B1(_00963_),
    .C1(_00973_),
    .Y(_00994_));
 sky130_fd_sc_hd__or2_1 _07165_ (.A(_00974_),
    .B(_00994_),
    .X(_00995_));
 sky130_fd_sc_hd__or3_1 _07166_ (.A(_00991_),
    .B(_00992_),
    .C(_00995_),
    .X(_00996_));
 sky130_fd_sc_hd__nand2_1 _07167_ (.A(_00871_),
    .B(_00873_),
    .Y(_00997_));
 sky130_fd_sc_hd__a211oi_2 _07168_ (.A1(_00874_),
    .A2(_00997_),
    .B1(_00950_),
    .C1(_00949_),
    .Y(_00998_));
 sky130_fd_sc_hd__o211a_1 _07169_ (.A1(_00949_),
    .A2(_00950_),
    .B1(_00997_),
    .C1(_00874_),
    .X(_01000_));
 sky130_fd_sc_hd__o211ai_1 _07170_ (.A1(_00949_),
    .A2(_00950_),
    .B1(_00997_),
    .C1(_00874_),
    .Y(_01001_));
 sky130_fd_sc_hd__a211o_1 _07171_ (.A1(_00975_),
    .A2(_00996_),
    .B1(_00998_),
    .C1(_01000_),
    .X(_01002_));
 sky130_fd_sc_hd__o221ai_4 _07172_ (.A1(_00993_),
    .A2(_00995_),
    .B1(_00998_),
    .B2(_01000_),
    .C1(_00975_),
    .Y(_01003_));
 sky130_fd_sc_hd__o211ai_2 _07173_ (.A1(_00836_),
    .A2(_00956_),
    .B1(_00955_),
    .C1(_00933_),
    .Y(_01004_));
 sky130_fd_sc_hd__nand4_2 _07174_ (.A(_00957_),
    .B(_01002_),
    .C(_01003_),
    .D(_01004_),
    .Y(_01005_));
 sky130_fd_sc_hd__nor2_1 _07175_ (.A(_00881_),
    .B(_00883_),
    .Y(_01006_));
 sky130_fd_sc_hd__a211oi_2 _07176_ (.A1(_00957_),
    .A2(_01005_),
    .B1(_01006_),
    .C1(_00884_),
    .Y(_01007_));
 sky130_fd_sc_hd__inv_2 _07177_ (.A(_01007_),
    .Y(_01008_));
 sky130_fd_sc_hd__o211a_1 _07178_ (.A1(_00884_),
    .A2(_01006_),
    .B1(_01005_),
    .C1(_00957_),
    .X(_01009_));
 sky130_fd_sc_hd__and4bb_1 _07179_ (.A_N(_00862_),
    .B_N(_00870_),
    .C(_01001_),
    .D(_01002_),
    .X(_01011_));
 sky130_fd_sc_hd__a2bb2oi_1 _07180_ (.A1_N(_00862_),
    .A2_N(_00870_),
    .B1(_01001_),
    .B2(_01002_),
    .Y(_01012_));
 sky130_fd_sc_hd__nor2_1 _07181_ (.A(_01011_),
    .B(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__o21a_1 _07182_ (.A1(_00864_),
    .A2(_00867_),
    .B1(_01013_),
    .X(_01014_));
 sky130_fd_sc_hd__a211oi_1 _07183_ (.A1(net28),
    .A2(_00866_),
    .B1(_01013_),
    .C1(_00864_),
    .Y(_01015_));
 sky130_fd_sc_hd__or4_1 _07184_ (.A(_01007_),
    .B(_01009_),
    .C(_01014_),
    .D(_01015_),
    .X(_01016_));
 sky130_fd_sc_hd__o311a_1 _07185_ (.A1(_01009_),
    .A2(_01014_),
    .A3(_01015_),
    .B1(_01008_),
    .C1(_00906_),
    .X(_01017_));
 sky130_fd_sc_hd__a21o_1 _07186_ (.A1(_01008_),
    .A2(_01016_),
    .B1(_00906_),
    .X(_01018_));
 sky130_fd_sc_hd__nor2_1 _07187_ (.A(_01012_),
    .B(_01014_),
    .Y(_01019_));
 sky130_fd_sc_hd__o21ai_1 _07188_ (.A1(_01017_),
    .A2(_01019_),
    .B1(_01018_),
    .Y(_01020_));
 sky130_fd_sc_hd__and2_1 _07189_ (.A(_00904_),
    .B(_01020_),
    .X(_01022_));
 sky130_fd_sc_hd__xor2_1 _07190_ (.A(_00904_),
    .B(_01020_),
    .X(_01023_));
 sky130_fd_sc_hd__a22o_1 _07191_ (.A1(_00927_),
    .A2(_00928_),
    .B1(_00929_),
    .B2(_00918_),
    .X(_01024_));
 sky130_fd_sc_hd__nand2_1 _07192_ (.A(_00930_),
    .B(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__a2bb2o_1 _07193_ (.A1_N(_00912_),
    .A2_N(_00914_),
    .B1(net55),
    .B2(_00909_),
    .X(_01026_));
 sky130_fd_sc_hd__a21o_1 _07194_ (.A1(net15),
    .A2(net55),
    .B1(net44),
    .X(_01027_));
 sky130_fd_sc_hd__o21ai_1 _07195_ (.A1(_01230_),
    .A2(_00909_),
    .B1(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand3_2 _07196_ (.A(net15),
    .B(net44),
    .C(net33),
    .Y(_01029_));
 sky130_fd_sc_hd__a21o_1 _07197_ (.A1(net15),
    .A2(net44),
    .B1(net33),
    .X(_01030_));
 sky130_fd_sc_hd__nand4_2 _07198_ (.A(_01030_),
    .B(net55),
    .C(net14),
    .D(_01029_),
    .Y(_01031_));
 sky130_fd_sc_hd__a21o_1 _07199_ (.A1(_01029_),
    .A2(_01031_),
    .B1(_01028_),
    .X(_01033_));
 sky130_fd_sc_hd__a22o_1 _07200_ (.A1(net13),
    .A2(net59),
    .B1(net58),
    .B2(net14),
    .X(_01034_));
 sky130_fd_sc_hd__nand4_2 _07201_ (.A(net14),
    .B(net13),
    .C(net59),
    .D(net58),
    .Y(_01035_));
 sky130_fd_sc_hd__nand4_2 _07202_ (.A(_01034_),
    .B(_01035_),
    .C(net11),
    .D(net60),
    .Y(_01036_));
 sky130_fd_sc_hd__a22o_1 _07203_ (.A1(net11),
    .A2(net60),
    .B1(_01034_),
    .B2(_01035_),
    .X(_01037_));
 sky130_fd_sc_hd__nand3_1 _07204_ (.A(_01028_),
    .B(_01029_),
    .C(_01031_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand4_1 _07205_ (.A(_01033_),
    .B(_01036_),
    .C(_01037_),
    .D(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__nand2_1 _07206_ (.A(_01033_),
    .B(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__and3_1 _07207_ (.A(_00915_),
    .B(_01026_),
    .C(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__nand4_2 _07208_ (.A(net10),
    .B(net9),
    .C(net62),
    .D(net61),
    .Y(_01042_));
 sky130_fd_sc_hd__a22o_1 _07209_ (.A1(net9),
    .A2(net62),
    .B1(net61),
    .B2(net10),
    .X(_01044_));
 sky130_fd_sc_hd__nand4_2 _07210_ (.A(_01044_),
    .B(net63),
    .C(net8),
    .D(_01042_),
    .Y(_01045_));
 sky130_fd_sc_hd__o22a_1 _07211_ (.A1(_01076_),
    .A2(_01142_),
    .B1(_00919_),
    .B2(_00920_),
    .X(_01046_));
 sky130_fd_sc_hd__o211a_1 _07212_ (.A1(_00922_),
    .A2(_01046_),
    .B1(_01036_),
    .C1(_01035_),
    .X(_01047_));
 sky130_fd_sc_hd__a211o_1 _07213_ (.A1(_01035_),
    .A2(_01036_),
    .B1(_01046_),
    .C1(_00922_),
    .X(_01048_));
 sky130_fd_sc_hd__inv_2 _07214_ (.A(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__a211o_1 _07215_ (.A1(_01042_),
    .A2(_01045_),
    .B1(_01047_),
    .C1(_01049_),
    .X(_01050_));
 sky130_fd_sc_hd__o211ai_2 _07216_ (.A1(_01047_),
    .A2(_01049_),
    .B1(_01042_),
    .C1(_01045_),
    .Y(_01051_));
 sky130_fd_sc_hd__a21o_1 _07217_ (.A1(_00915_),
    .A2(_01026_),
    .B1(_01040_),
    .X(_01052_));
 sky130_fd_sc_hd__and2b_1 _07218_ (.A_N(_01041_),
    .B(_01052_),
    .X(_01053_));
 sky130_fd_sc_hd__nand3_1 _07219_ (.A(_01053_),
    .B(_01051_),
    .C(_01050_),
    .Y(_01055_));
 sky130_fd_sc_hd__a31o_1 _07220_ (.A1(_01050_),
    .A2(_01051_),
    .A3(_01052_),
    .B1(_01041_),
    .X(_01056_));
 sky130_fd_sc_hd__and3_1 _07221_ (.A(_00930_),
    .B(_01024_),
    .C(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__nand2_1 _07222_ (.A(net6),
    .B(net34),
    .Y(_01058_));
 sky130_fd_sc_hd__nand4_2 _07223_ (.A(net7),
    .B(net6),
    .C(net34),
    .D(net64),
    .Y(_01059_));
 sky130_fd_sc_hd__a22o_1 _07224_ (.A1(net6),
    .A2(net34),
    .B1(net64),
    .B2(net7),
    .X(_01060_));
 sky130_fd_sc_hd__nand4_2 _07225_ (.A(_01060_),
    .B(net35),
    .C(net5),
    .D(_01059_),
    .Y(_01061_));
 sky130_fd_sc_hd__o2bb2a_1 _07226_ (.A1_N(net6),
    .A2_N(net35),
    .B1(_00934_),
    .B2(_00935_),
    .X(_01062_));
 sky130_fd_sc_hd__a211oi_1 _07227_ (.A1(_01059_),
    .A2(_01061_),
    .B1(_01062_),
    .C1(_00937_),
    .Y(_01063_));
 sky130_fd_sc_hd__a2bb2o_1 _07228_ (.A1_N(_00958_),
    .A2_N(_00960_),
    .B1(net38),
    .B2(net3),
    .X(_01064_));
 sky130_fd_sc_hd__nand2_1 _07229_ (.A(_00961_),
    .B(_01064_),
    .Y(_01066_));
 sky130_fd_sc_hd__o211a_1 _07230_ (.A1(_00937_),
    .A2(_01062_),
    .B1(_01061_),
    .C1(_01059_),
    .X(_01067_));
 sky130_fd_sc_hd__nor3_1 _07231_ (.A(_01063_),
    .B(_01066_),
    .C(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__nor2_1 _07232_ (.A(_01063_),
    .B(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__and2_1 _07233_ (.A(_00942_),
    .B(_00944_),
    .X(_01070_));
 sky130_fd_sc_hd__o211a_1 _07234_ (.A1(_00945_),
    .A2(_01070_),
    .B1(_01050_),
    .C1(_01048_),
    .X(_01071_));
 sky130_fd_sc_hd__a211oi_2 _07235_ (.A1(_01048_),
    .A2(_01050_),
    .B1(_01070_),
    .C1(_00945_),
    .Y(_01072_));
 sky130_fd_sc_hd__nor3_1 _07236_ (.A(_01069_),
    .B(_01071_),
    .C(_01072_),
    .Y(_01073_));
 sky130_fd_sc_hd__o21a_1 _07237_ (.A1(_01071_),
    .A2(_01072_),
    .B1(_01069_),
    .X(_01074_));
 sky130_fd_sc_hd__nor2_1 _07238_ (.A(_01073_),
    .B(_01074_),
    .Y(_01075_));
 sky130_fd_sc_hd__xnor2_1 _07239_ (.A(_01025_),
    .B(_01056_),
    .Y(_01077_));
 sky130_fd_sc_hd__and2_1 _07240_ (.A(_01075_),
    .B(_01077_),
    .X(_01078_));
 sky130_fd_sc_hd__or2_1 _07241_ (.A(_00952_),
    .B(_00954_),
    .X(_01079_));
 sky130_fd_sc_hd__o211a_1 _07242_ (.A1(_01057_),
    .A2(_01078_),
    .B1(_01079_),
    .C1(_00955_),
    .X(_01080_));
 sky130_fd_sc_hd__nand4_2 _07243_ (.A(net37),
    .B(net36),
    .C(net4),
    .D(net3),
    .Y(_01081_));
 sky130_fd_sc_hd__a22o_1 _07244_ (.A1(net36),
    .A2(net4),
    .B1(net3),
    .B2(net37),
    .X(_01082_));
 sky130_fd_sc_hd__nand4_2 _07245_ (.A(_01082_),
    .B(net2),
    .C(net38),
    .D(_01081_),
    .Y(_01083_));
 sky130_fd_sc_hd__a22oi_1 _07246_ (.A1(net41),
    .A2(net31),
    .B1(_00964_),
    .B2(_00965_),
    .Y(_01084_));
 sky130_fd_sc_hd__a211oi_1 _07247_ (.A1(_01081_),
    .A2(_01083_),
    .B1(_01084_),
    .C1(_00967_),
    .Y(_01085_));
 sky130_fd_sc_hd__and4_1 _07248_ (.A(net40),
    .B(net39),
    .C(net32),
    .D(net31),
    .X(_01086_));
 sky130_fd_sc_hd__nand4_1 _07249_ (.A(net40),
    .B(net39),
    .C(net32),
    .D(net31),
    .Y(_01088_));
 sky130_fd_sc_hd__a22o_1 _07250_ (.A1(net39),
    .A2(net32),
    .B1(net31),
    .B2(net40),
    .X(_01089_));
 sky130_fd_sc_hd__and4_1 _07251_ (.A(_01089_),
    .B(net30),
    .C(net41),
    .D(_01088_),
    .X(_01090_));
 sky130_fd_sc_hd__a31o_1 _07252_ (.A1(_01089_),
    .A2(net30),
    .A3(net41),
    .B1(_01086_),
    .X(_01091_));
 sky130_fd_sc_hd__o211a_1 _07253_ (.A1(_00967_),
    .A2(_01084_),
    .B1(_01083_),
    .C1(_01081_),
    .X(_01092_));
 sky130_fd_sc_hd__nor2_1 _07254_ (.A(_01085_),
    .B(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__o21a_1 _07255_ (.A1(_01086_),
    .A2(_01090_),
    .B1(_01093_),
    .X(_01094_));
 sky130_fd_sc_hd__a21oi_1 _07256_ (.A1(_01093_),
    .A2(_01091_),
    .B1(_01085_),
    .Y(_01095_));
 sky130_fd_sc_hd__nor2_1 _07257_ (.A(_00968_),
    .B(_00970_),
    .Y(_01096_));
 sky130_fd_sc_hd__nor2_1 _07258_ (.A(_00971_),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__o21ai_1 _07259_ (.A1(_01085_),
    .A2(_01094_),
    .B1(_01097_),
    .Y(_01099_));
 sky130_fd_sc_hd__and4_1 _07260_ (.A(net43),
    .B(net42),
    .C(net30),
    .D(net29),
    .X(_01100_));
 sky130_fd_sc_hd__nand4_1 _07261_ (.A(net43),
    .B(net42),
    .C(net30),
    .D(net29),
    .Y(_01101_));
 sky130_fd_sc_hd__o2bb2a_1 _07262_ (.A1_N(net42),
    .A2_N(net30),
    .B1(_01186_),
    .B2(_01065_),
    .X(_01102_));
 sky130_fd_sc_hd__and4b_1 _07263_ (.A_N(_01102_),
    .B(net28),
    .C(net45),
    .D(_01101_),
    .X(_01103_));
 sky130_fd_sc_hd__or4b_1 _07264_ (.A(_01054_),
    .B(_01100_),
    .C(_01102_),
    .D_N(net28),
    .X(_01104_));
 sky130_fd_sc_hd__o22a_1 _07265_ (.A1(_01054_),
    .A2(_01186_),
    .B1(_00976_),
    .B2(_00979_),
    .X(_01105_));
 sky130_fd_sc_hd__o211a_1 _07266_ (.A1(_00980_),
    .A2(_01105_),
    .B1(_01104_),
    .C1(_01101_),
    .X(_01106_));
 sky130_fd_sc_hd__a211oi_1 _07267_ (.A1(_01101_),
    .A2(_01104_),
    .B1(_01105_),
    .C1(_00980_),
    .Y(_01107_));
 sky130_fd_sc_hd__nor2_1 _07268_ (.A(_01106_),
    .B(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__and4_1 _07269_ (.A(net46),
    .B(net47),
    .C(net28),
    .D(net27),
    .X(_01110_));
 sky130_fd_sc_hd__o2bb2a_1 _07270_ (.A1_N(net46),
    .A2_N(net28),
    .B1(_01208_),
    .B2(_01043_),
    .X(_01111_));
 sky130_fd_sc_hd__or3_1 _07271_ (.A(_01219_),
    .B(_01110_),
    .C(_01111_),
    .X(_01112_));
 sky130_fd_sc_hd__o21ai_1 _07272_ (.A1(_01110_),
    .A2(_01111_),
    .B1(_01219_),
    .Y(_01113_));
 sky130_fd_sc_hd__a21oi_1 _07273_ (.A1(_01112_),
    .A2(_01113_),
    .B1(_01108_),
    .Y(_01114_));
 sky130_fd_sc_hd__and3_1 _07274_ (.A(_01108_),
    .B(_01112_),
    .C(_01113_),
    .X(_01115_));
 sky130_fd_sc_hd__or2_1 _07275_ (.A(_01114_),
    .B(_01115_),
    .X(_01116_));
 sky130_fd_sc_hd__xor2_1 _07276_ (.A(_01095_),
    .B(_01097_),
    .X(_01117_));
 sky130_fd_sc_hd__o21ai_1 _07277_ (.A1(_01116_),
    .A2(_01117_),
    .B1(_01099_),
    .Y(_01118_));
 sky130_fd_sc_hd__o21ai_1 _07278_ (.A1(_00991_),
    .A2(_00992_),
    .B1(_00995_),
    .Y(_01119_));
 sky130_fd_sc_hd__a211oi_1 _07279_ (.A1(_00996_),
    .A2(_01119_),
    .B1(_01073_),
    .C1(_01072_),
    .Y(_01121_));
 sky130_fd_sc_hd__o211a_1 _07280_ (.A1(_01072_),
    .A2(_01073_),
    .B1(_01119_),
    .C1(_00996_),
    .X(_01122_));
 sky130_fd_sc_hd__nor2_1 _07281_ (.A(_01121_),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__and2_1 _07282_ (.A(_01123_),
    .B(_01118_),
    .X(_01124_));
 sky130_fd_sc_hd__nor2_1 _07283_ (.A(_01118_),
    .B(_01123_),
    .Y(_01125_));
 sky130_fd_sc_hd__or2_1 _07284_ (.A(_01124_),
    .B(_01125_),
    .X(_01126_));
 sky130_fd_sc_hd__a221oi_2 _07285_ (.A1(_01075_),
    .A2(_01077_),
    .B1(_01079_),
    .B2(_00955_),
    .C1(_01057_),
    .Y(_01127_));
 sky130_fd_sc_hd__or3_1 _07286_ (.A(_01080_),
    .B(_01127_),
    .C(_01126_),
    .X(_01128_));
 sky130_fd_sc_hd__o21bai_1 _07287_ (.A1(_01127_),
    .A2(_01126_),
    .B1_N(_01080_),
    .Y(_01129_));
 sky130_fd_sc_hd__a22o_1 _07288_ (.A1(_01002_),
    .A2(_01003_),
    .B1(_01004_),
    .B2(_00957_),
    .X(_01130_));
 sky130_fd_sc_hd__and3_1 _07289_ (.A(_01005_),
    .B(_01129_),
    .C(_01130_),
    .X(_01132_));
 sky130_fd_sc_hd__a21oi_1 _07290_ (.A1(_01005_),
    .A2(_01130_),
    .B1(_01129_),
    .Y(_01133_));
 sky130_fd_sc_hd__or2_1 _07291_ (.A(_01132_),
    .B(_01133_),
    .X(_01134_));
 sky130_fd_sc_hd__a41o_1 _07292_ (.A1(net46),
    .A2(net47),
    .A3(net29),
    .A4(net28),
    .B1(_00987_),
    .X(_01135_));
 sky130_fd_sc_hd__nor4_1 _07293_ (.A(_00984_),
    .B(_00992_),
    .C(_01122_),
    .D(_01124_),
    .Y(_01136_));
 sky130_fd_sc_hd__o22a_1 _07294_ (.A1(_00984_),
    .A2(_00992_),
    .B1(_01122_),
    .B2(_01124_),
    .X(_01137_));
 sky130_fd_sc_hd__nor2_1 _07295_ (.A(_01136_),
    .B(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__o21a_1 _07296_ (.A1(_00985_),
    .A2(_00987_),
    .B1(_01138_),
    .X(_01139_));
 sky130_fd_sc_hd__nor2_1 _07297_ (.A(_01135_),
    .B(_01138_),
    .Y(_01140_));
 sky130_fd_sc_hd__or2_1 _07298_ (.A(_01139_),
    .B(_01140_),
    .X(_01141_));
 sky130_fd_sc_hd__nor2_1 _07299_ (.A(_01134_),
    .B(_01141_),
    .Y(_01143_));
 sky130_fd_sc_hd__o22ai_1 _07300_ (.A1(_01007_),
    .A2(_01009_),
    .B1(_01014_),
    .B2(_01015_),
    .Y(_01144_));
 sky130_fd_sc_hd__and2_1 _07301_ (.A(_01016_),
    .B(_01144_),
    .X(_01145_));
 sky130_fd_sc_hd__o211a_1 _07302_ (.A1(_01132_),
    .A2(_01143_),
    .B1(_01144_),
    .C1(_01016_),
    .X(_01146_));
 sky130_fd_sc_hd__a311oi_1 _07303_ (.A1(_01005_),
    .A2(_01129_),
    .A3(_01130_),
    .B1(_01143_),
    .C1(_01145_),
    .Y(_01147_));
 sky130_fd_sc_hd__nor2_1 _07304_ (.A(_01146_),
    .B(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__o21a_1 _07305_ (.A1(_01137_),
    .A2(_01139_),
    .B1(_01148_),
    .X(_01149_));
 sky130_fd_sc_hd__or2_1 _07306_ (.A(_01146_),
    .B(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__nand2b_1 _07307_ (.A_N(_01017_),
    .B(_01018_),
    .Y(_01151_));
 sky130_fd_sc_hd__xor2_1 _07308_ (.A(_01019_),
    .B(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__o21a_1 _07309_ (.A1(_01146_),
    .A2(_01149_),
    .B1(_01152_),
    .X(_01154_));
 sky130_fd_sc_hd__nor2_1 _07310_ (.A(_01150_),
    .B(_01152_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _07311_ (.A(_01154_),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__o21ai_1 _07312_ (.A1(_01080_),
    .A2(_01127_),
    .B1(_01126_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand2_1 _07313_ (.A(_01128_),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__a21o_1 _07314_ (.A1(_01050_),
    .A2(_01051_),
    .B1(_01053_),
    .X(_01159_));
 sky130_fd_sc_hd__a22o_1 _07315_ (.A1(_01036_),
    .A2(_01037_),
    .B1(_01038_),
    .B2(_01033_),
    .X(_01160_));
 sky130_fd_sc_hd__nand2_1 _07316_ (.A(net14),
    .B(net33),
    .Y(_01161_));
 sky130_fd_sc_hd__nand4_1 _07317_ (.A(net15),
    .B(net14),
    .C(net44),
    .D(net33),
    .Y(_01162_));
 sky130_fd_sc_hd__a22o_1 _07318_ (.A1(net14),
    .A2(net44),
    .B1(net33),
    .B2(net15),
    .X(_01163_));
 sky130_fd_sc_hd__o2111ai_4 _07319_ (.A1(_00909_),
    .A2(_01161_),
    .B1(net13),
    .C1(net55),
    .D1(_01163_),
    .Y(_01165_));
 sky130_fd_sc_hd__o21ai_1 _07320_ (.A1(_00909_),
    .A2(_01161_),
    .B1(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__a22o_1 _07321_ (.A1(net14),
    .A2(net55),
    .B1(_01029_),
    .B2(_01030_),
    .X(_01167_));
 sky130_fd_sc_hd__and3_1 _07322_ (.A(_01031_),
    .B(_01166_),
    .C(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__nand3_1 _07323_ (.A(_01031_),
    .B(_01166_),
    .C(_01167_),
    .Y(_01169_));
 sky130_fd_sc_hd__a21o_1 _07324_ (.A1(_01031_),
    .A2(_01167_),
    .B1(_01166_),
    .X(_01170_));
 sky130_fd_sc_hd__a22oi_2 _07325_ (.A1(net11),
    .A2(net59),
    .B1(net58),
    .B2(net13),
    .Y(_01171_));
 sky130_fd_sc_hd__a22o_1 _07326_ (.A1(net11),
    .A2(net59),
    .B1(net58),
    .B2(net13),
    .X(_01172_));
 sky130_fd_sc_hd__and4_1 _07327_ (.A(net13),
    .B(net11),
    .C(net59),
    .D(net58),
    .X(_01173_));
 sky130_fd_sc_hd__a211oi_2 _07328_ (.A1(net10),
    .A2(net60),
    .B1(_01171_),
    .C1(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__o211a_1 _07329_ (.A1(_01171_),
    .A2(_01173_),
    .B1(net10),
    .C1(net60),
    .X(_01176_));
 sky130_fd_sc_hd__o211a_1 _07330_ (.A1(_01174_),
    .A2(_01176_),
    .B1(_01169_),
    .C1(_01170_),
    .X(_01177_));
 sky130_fd_sc_hd__o211ai_2 _07331_ (.A1(_01174_),
    .A2(_01176_),
    .B1(_01169_),
    .C1(_01170_),
    .Y(_01178_));
 sky130_fd_sc_hd__o211a_1 _07332_ (.A1(_01168_),
    .A2(_01177_),
    .B1(_01039_),
    .C1(_01160_),
    .X(_01179_));
 sky130_fd_sc_hd__and4_1 _07333_ (.A(net9),
    .B(net8),
    .C(net62),
    .D(net61),
    .X(_01180_));
 sky130_fd_sc_hd__nand4_1 _07334_ (.A(net9),
    .B(net8),
    .C(net62),
    .D(net61),
    .Y(_01181_));
 sky130_fd_sc_hd__a22o_1 _07335_ (.A1(net8),
    .A2(net62),
    .B1(net61),
    .B2(net9),
    .X(_01182_));
 sky130_fd_sc_hd__and4_1 _07336_ (.A(_01182_),
    .B(net63),
    .C(net7),
    .D(_01181_),
    .X(_01183_));
 sky130_fd_sc_hd__nand4_1 _07337_ (.A(_01182_),
    .B(net63),
    .C(net7),
    .D(_01181_),
    .Y(_01184_));
 sky130_fd_sc_hd__a31o_1 _07338_ (.A1(_01172_),
    .A2(net60),
    .A3(net10),
    .B1(_01173_),
    .X(_01185_));
 sky130_fd_sc_hd__a22o_1 _07339_ (.A1(net8),
    .A2(net63),
    .B1(_01042_),
    .B2(_01044_),
    .X(_01187_));
 sky130_fd_sc_hd__a21o_1 _07340_ (.A1(_01045_),
    .A2(_01187_),
    .B1(_01185_),
    .X(_01188_));
 sky130_fd_sc_hd__nand3_2 _07341_ (.A(_01045_),
    .B(_01185_),
    .C(_01187_),
    .Y(_01189_));
 sky130_fd_sc_hd__o211ai_4 _07342_ (.A1(_01180_),
    .A2(_01183_),
    .B1(_01188_),
    .C1(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__a211o_1 _07343_ (.A1(_01188_),
    .A2(_01189_),
    .B1(_01180_),
    .C1(_01183_),
    .X(_01191_));
 sky130_fd_sc_hd__and2_1 _07344_ (.A(_01190_),
    .B(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__a211oi_1 _07345_ (.A1(_01039_),
    .A2(_01160_),
    .B1(_01168_),
    .C1(_01177_),
    .Y(_01193_));
 sky130_fd_sc_hd__nor2_1 _07346_ (.A(_01179_),
    .B(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__and3_1 _07347_ (.A(_01194_),
    .B(_01191_),
    .C(_01190_),
    .X(_01195_));
 sky130_fd_sc_hd__or3b_1 _07348_ (.A(_01179_),
    .B(_01193_),
    .C_N(_01192_),
    .X(_01196_));
 sky130_fd_sc_hd__o211a_1 _07349_ (.A1(_01179_),
    .A2(_01195_),
    .B1(_01055_),
    .C1(_01159_),
    .X(_01198_));
 sky130_fd_sc_hd__o211ai_1 _07350_ (.A1(_01179_),
    .A2(_01195_),
    .B1(_01055_),
    .C1(_01159_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _07351_ (.A(net5),
    .B(net64),
    .Y(_01200_));
 sky130_fd_sc_hd__or2_1 _07352_ (.A(_01058_),
    .B(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__a22o_1 _07353_ (.A1(net5),
    .A2(net34),
    .B1(net64),
    .B2(net6),
    .X(_01202_));
 sky130_fd_sc_hd__o2111ai_2 _07354_ (.A1(_01058_),
    .A2(_01200_),
    .B1(net4),
    .C1(net35),
    .D1(_01202_),
    .Y(_01203_));
 sky130_fd_sc_hd__o21ai_1 _07355_ (.A1(_01058_),
    .A2(_01200_),
    .B1(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__a22o_1 _07356_ (.A1(net5),
    .A2(net35),
    .B1(_01059_),
    .B2(_01060_),
    .X(_01205_));
 sky130_fd_sc_hd__nand3_2 _07357_ (.A(_01061_),
    .B(_01204_),
    .C(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__a22o_1 _07358_ (.A1(net38),
    .A2(net2),
    .B1(_01081_),
    .B2(_01082_),
    .X(_01207_));
 sky130_fd_sc_hd__a21o_1 _07359_ (.A1(_01061_),
    .A2(_01205_),
    .B1(_01204_),
    .X(_01209_));
 sky130_fd_sc_hd__nand4_2 _07360_ (.A(_01083_),
    .B(_01206_),
    .C(_01207_),
    .D(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__o2bb2a_1 _07361_ (.A1_N(_00961_),
    .A2_N(_01064_),
    .B1(_01067_),
    .B2(_01063_),
    .X(_01211_));
 sky130_fd_sc_hd__a211oi_2 _07362_ (.A1(_01189_),
    .A2(_01190_),
    .B1(_01211_),
    .C1(_01068_),
    .Y(_01212_));
 sky130_fd_sc_hd__o211a_1 _07363_ (.A1(_01068_),
    .A2(_01211_),
    .B1(_01190_),
    .C1(_01189_),
    .X(_01213_));
 sky130_fd_sc_hd__a211o_1 _07364_ (.A1(_01206_),
    .A2(_01210_),
    .B1(_01212_),
    .C1(_01213_),
    .X(_01214_));
 sky130_fd_sc_hd__o211ai_2 _07365_ (.A1(_01212_),
    .A2(_01213_),
    .B1(_01206_),
    .C1(_01210_),
    .Y(_01215_));
 sky130_fd_sc_hd__a221o_1 _07366_ (.A1(_01192_),
    .A2(_01194_),
    .B1(_01055_),
    .B2(_01159_),
    .C1(_01179_),
    .X(_01216_));
 sky130_fd_sc_hd__and4_1 _07367_ (.A(_01199_),
    .B(_01214_),
    .C(_01215_),
    .D(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__nor2_1 _07368_ (.A(_01075_),
    .B(_01077_),
    .Y(_01218_));
 sky130_fd_sc_hd__nor2_1 _07369_ (.A(_01078_),
    .B(_01218_),
    .Y(_01220_));
 sky130_fd_sc_hd__o21a_1 _07370_ (.A1(_01198_),
    .A2(_01217_),
    .B1(_01220_),
    .X(_01221_));
 sky130_fd_sc_hd__o21ai_1 _07371_ (.A1(_01198_),
    .A2(_01217_),
    .B1(_01220_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand4_2 _07372_ (.A(net37),
    .B(net36),
    .C(net3),
    .D(net2),
    .Y(_01223_));
 sky130_fd_sc_hd__a22o_1 _07373_ (.A1(net36),
    .A2(net3),
    .B1(net2),
    .B2(net37),
    .X(_01224_));
 sky130_fd_sc_hd__nand4_2 _07374_ (.A(_01224_),
    .B(net32),
    .C(net38),
    .D(_01223_),
    .Y(_01225_));
 sky130_fd_sc_hd__a22oi_1 _07375_ (.A1(net41),
    .A2(net30),
    .B1(_01088_),
    .B2(_01089_),
    .Y(_01226_));
 sky130_fd_sc_hd__a211o_1 _07376_ (.A1(_01223_),
    .A2(_01225_),
    .B1(_01226_),
    .C1(_01090_),
    .X(_01227_));
 sky130_fd_sc_hd__and4_1 _07377_ (.A(net40),
    .B(net39),
    .C(net31),
    .D(net30),
    .X(_01228_));
 sky130_fd_sc_hd__nand4_1 _07378_ (.A(net40),
    .B(net39),
    .C(net31),
    .D(net30),
    .Y(_01229_));
 sky130_fd_sc_hd__a22o_1 _07379_ (.A1(net39),
    .A2(net31),
    .B1(net30),
    .B2(net40),
    .X(_01231_));
 sky130_fd_sc_hd__nand4_1 _07380_ (.A(_01231_),
    .B(net29),
    .C(net41),
    .D(_01229_),
    .Y(_01232_));
 sky130_fd_sc_hd__o211ai_1 _07381_ (.A1(_01090_),
    .A2(_01226_),
    .B1(_01225_),
    .C1(_01223_),
    .Y(_01233_));
 sky130_fd_sc_hd__and2_1 _07382_ (.A(_01227_),
    .B(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__a21bo_1 _07383_ (.A1(_01229_),
    .A2(_01232_),
    .B1_N(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__nand2_1 _07384_ (.A(_01227_),
    .B(_01235_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_1 _07385_ (.A(_01091_),
    .B(_01093_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(_01094_),
    .B(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__and2_1 _07387_ (.A(_01236_),
    .B(_01238_),
    .X(_01239_));
 sky130_fd_sc_hd__nand4_2 _07388_ (.A(net43),
    .B(net42),
    .C(net29),
    .D(net28),
    .Y(_01240_));
 sky130_fd_sc_hd__a22o_1 _07389_ (.A1(net42),
    .A2(net29),
    .B1(net28),
    .B2(net43),
    .X(_01242_));
 sky130_fd_sc_hd__nand4_2 _07390_ (.A(_01242_),
    .B(net27),
    .C(net45),
    .D(_01240_),
    .Y(_01243_));
 sky130_fd_sc_hd__o2bb2a_1 _07391_ (.A1_N(net45),
    .A2_N(net28),
    .B1(_01100_),
    .B2(_01102_),
    .X(_01244_));
 sky130_fd_sc_hd__o211a_1 _07392_ (.A1(_01103_),
    .A2(_01244_),
    .B1(_01243_),
    .C1(_01240_),
    .X(_01245_));
 sky130_fd_sc_hd__a211oi_1 _07393_ (.A1(_01240_),
    .A2(_01243_),
    .B1(_01244_),
    .C1(_01103_),
    .Y(_01246_));
 sky130_fd_sc_hd__nand2_1 _07394_ (.A(net46),
    .B(net26),
    .Y(_01247_));
 sky130_fd_sc_hd__a22o_1 _07395_ (.A1(net46),
    .A2(net27),
    .B1(net26),
    .B2(net47),
    .X(_01248_));
 sky130_fd_sc_hd__o31a_1 _07396_ (.A1(_01043_),
    .A2(_01208_),
    .A3(_01247_),
    .B1(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__and2_1 _07397_ (.A(net23),
    .B(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__nor2_1 _07398_ (.A(net23),
    .B(_01249_),
    .Y(_01251_));
 sky130_fd_sc_hd__or2_1 _07399_ (.A(_01250_),
    .B(_01251_),
    .X(_01253_));
 sky130_fd_sc_hd__o21a_1 _07400_ (.A1(_01245_),
    .A2(_01246_),
    .B1(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__nor3_1 _07401_ (.A(_01245_),
    .B(_01246_),
    .C(_01253_),
    .Y(_01255_));
 sky130_fd_sc_hd__xnor2_1 _07402_ (.A(_01236_),
    .B(_01238_),
    .Y(_01256_));
 sky130_fd_sc_hd__nor3_2 _07403_ (.A(_01254_),
    .B(_01255_),
    .C(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__and2b_1 _07404_ (.A_N(_01212_),
    .B(_01214_),
    .X(_01258_));
 sky130_fd_sc_hd__xnor2_1 _07405_ (.A(_01116_),
    .B(_01117_),
    .Y(_01259_));
 sky130_fd_sc_hd__nor2_1 _07406_ (.A(_01258_),
    .B(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__and3b_1 _07407_ (.A_N(_01212_),
    .B(_01214_),
    .C(_01259_),
    .X(_01261_));
 sky130_fd_sc_hd__nor2_1 _07408_ (.A(_01260_),
    .B(_01261_),
    .Y(_01262_));
 sky130_fd_sc_hd__o21a_1 _07409_ (.A1(_01239_),
    .A2(_01257_),
    .B1(_01262_),
    .X(_01264_));
 sky130_fd_sc_hd__a211oi_1 _07410_ (.A1(_01236_),
    .A2(_01238_),
    .B1(_01257_),
    .C1(_01262_),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _07411_ (.A(_01264_),
    .B(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__inv_2 _07412_ (.A(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__a311o_1 _07413_ (.A1(_01214_),
    .A2(_01215_),
    .A3(_01216_),
    .B1(_01220_),
    .C1(_01198_),
    .X(_01268_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(_01222_),
    .B(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_1 _07415_ (.A(_01267_),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__o21bai_1 _07416_ (.A1(_01221_),
    .A2(_01270_),
    .B1_N(_01158_),
    .Y(_01271_));
 sky130_fd_sc_hd__o211ai_1 _07417_ (.A1(_01267_),
    .A2(_01269_),
    .B1(_01158_),
    .C1(_01222_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _07418_ (.A(_01271_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__o21bai_1 _07419_ (.A1(_01219_),
    .A2(_01111_),
    .B1_N(_01110_),
    .Y(_01275_));
 sky130_fd_sc_hd__o22a_1 _07420_ (.A1(_01107_),
    .A2(_01115_),
    .B1(_01260_),
    .B2(_01264_),
    .X(_01276_));
 sky130_fd_sc_hd__nor4_1 _07421_ (.A(_01107_),
    .B(_01115_),
    .C(_01260_),
    .D(_01264_),
    .Y(_01277_));
 sky130_fd_sc_hd__nor2_1 _07422_ (.A(_01276_),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__xnor2_1 _07423_ (.A(_01275_),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__or2_1 _07424_ (.A(_01273_),
    .B(_01279_),
    .X(_01280_));
 sky130_fd_sc_hd__and2_1 _07425_ (.A(_01134_),
    .B(_01141_),
    .X(_01281_));
 sky130_fd_sc_hd__or2_1 _07426_ (.A(_01143_),
    .B(_01281_),
    .X(_01282_));
 sky130_fd_sc_hd__a21o_1 _07427_ (.A1(_01271_),
    .A2(_01280_),
    .B1(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__a21oi_1 _07428_ (.A1(_01278_),
    .A2(_01275_),
    .B1(_01276_),
    .Y(_01284_));
 sky130_fd_sc_hd__o211ai_1 _07429_ (.A1(_01273_),
    .A2(_01279_),
    .B1(_01282_),
    .C1(_01271_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _07430_ (.A(_01283_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__or2_1 _07431_ (.A(_01284_),
    .B(_01287_),
    .X(_01288_));
 sky130_fd_sc_hd__a211oi_1 _07432_ (.A1(_01138_),
    .A2(_01135_),
    .B1(_01137_),
    .C1(_01148_),
    .Y(_01289_));
 sky130_fd_sc_hd__or2_1 _07433_ (.A(_01149_),
    .B(_01289_),
    .X(_01290_));
 sky130_fd_sc_hd__a21oi_1 _07434_ (.A1(_01283_),
    .A2(_01288_),
    .B1(_01290_),
    .Y(_01291_));
 sky130_fd_sc_hd__and3_1 _07435_ (.A(_01283_),
    .B(_01288_),
    .C(_01290_),
    .X(_01292_));
 sky130_fd_sc_hd__nor2_1 _07436_ (.A(_01291_),
    .B(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__a22oi_1 _07437_ (.A1(_01214_),
    .A2(_01215_),
    .B1(_01216_),
    .B2(_01199_),
    .Y(_01294_));
 sky130_fd_sc_hd__or2_1 _07438_ (.A(_01217_),
    .B(_01294_),
    .X(_01295_));
 sky130_fd_sc_hd__nand2_2 _07439_ (.A(net13),
    .B(net44),
    .Y(_01297_));
 sky130_fd_sc_hd__nand4_1 _07440_ (.A(net14),
    .B(net13),
    .C(net44),
    .D(net33),
    .Y(_01298_));
 sky130_fd_sc_hd__a22o_1 _07441_ (.A1(net13),
    .A2(net44),
    .B1(net33),
    .B2(net14),
    .X(_01299_));
 sky130_fd_sc_hd__nand4_2 _07442_ (.A(_01299_),
    .B(net55),
    .C(net11),
    .D(_01298_),
    .Y(_01300_));
 sky130_fd_sc_hd__o21ai_1 _07443_ (.A1(_01161_),
    .A2(_01297_),
    .B1(_01300_),
    .Y(_01301_));
 sky130_fd_sc_hd__a22o_1 _07444_ (.A1(net13),
    .A2(net55),
    .B1(_01162_),
    .B2(_01163_),
    .X(_01302_));
 sky130_fd_sc_hd__and3_1 _07445_ (.A(_01165_),
    .B(_01301_),
    .C(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__nand3_1 _07446_ (.A(_01165_),
    .B(_01301_),
    .C(_01302_),
    .Y(_01304_));
 sky130_fd_sc_hd__a22o_1 _07447_ (.A1(net10),
    .A2(net59),
    .B1(net58),
    .B2(net11),
    .X(_01305_));
 sky130_fd_sc_hd__nand4_1 _07448_ (.A(net11),
    .B(net10),
    .C(net59),
    .D(net58),
    .Y(_01306_));
 sky130_fd_sc_hd__nand4_1 _07449_ (.A(_01305_),
    .B(_01306_),
    .C(net9),
    .D(net60),
    .Y(_01308_));
 sky130_fd_sc_hd__a22o_1 _07450_ (.A1(net9),
    .A2(net60),
    .B1(_01305_),
    .B2(_01306_),
    .X(_01309_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__a21o_1 _07452_ (.A1(_01165_),
    .A2(_01302_),
    .B1(_01301_),
    .X(_01311_));
 sky130_fd_sc_hd__a31o_1 _07453_ (.A1(_01308_),
    .A2(_01309_),
    .A3(_01311_),
    .B1(_01303_),
    .X(_01312_));
 sky130_fd_sc_hd__a211o_1 _07454_ (.A1(_01169_),
    .A2(_01170_),
    .B1(_01174_),
    .C1(_01176_),
    .X(_01313_));
 sky130_fd_sc_hd__nand3_1 _07455_ (.A(_01178_),
    .B(_01312_),
    .C(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__a21o_1 _07456_ (.A1(_01178_),
    .A2(_01313_),
    .B1(_01312_),
    .X(_01315_));
 sky130_fd_sc_hd__nand4_2 _07457_ (.A(net8),
    .B(net7),
    .C(net62),
    .D(net61),
    .Y(_01316_));
 sky130_fd_sc_hd__a22o_1 _07458_ (.A1(net7),
    .A2(net62),
    .B1(net61),
    .B2(net8),
    .X(_01317_));
 sky130_fd_sc_hd__nand4_2 _07459_ (.A(_01317_),
    .B(net63),
    .C(net6),
    .D(_01316_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand2_1 _07460_ (.A(_01316_),
    .B(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand2_1 _07461_ (.A(_01306_),
    .B(_01308_),
    .Y(_01321_));
 sky130_fd_sc_hd__a22o_1 _07462_ (.A1(net7),
    .A2(net63),
    .B1(_01181_),
    .B2(_01182_),
    .X(_01322_));
 sky130_fd_sc_hd__a21o_1 _07463_ (.A1(_01184_),
    .A2(_01322_),
    .B1(_01321_),
    .X(_01323_));
 sky130_fd_sc_hd__nand3_1 _07464_ (.A(_01184_),
    .B(_01321_),
    .C(_01322_),
    .Y(_01324_));
 sky130_fd_sc_hd__a22oi_1 _07465_ (.A1(_01316_),
    .A2(_01319_),
    .B1(_01323_),
    .B2(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__and3b_1 _07466_ (.A_N(_01320_),
    .B(_01323_),
    .C(_01324_),
    .X(_01326_));
 sky130_fd_sc_hd__o211a_1 _07467_ (.A1(_01325_),
    .A2(_01326_),
    .B1(_01314_),
    .C1(_01315_),
    .X(_01327_));
 sky130_fd_sc_hd__a31o_1 _07468_ (.A1(_01178_),
    .A2(_01312_),
    .A3(_01313_),
    .B1(_01327_),
    .X(_01328_));
 sky130_fd_sc_hd__a21o_1 _07469_ (.A1(_01190_),
    .A2(_01191_),
    .B1(_01194_),
    .X(_01330_));
 sky130_fd_sc_hd__and3_1 _07470_ (.A(_01196_),
    .B(_01328_),
    .C(_01330_),
    .X(_01331_));
 sky130_fd_sc_hd__nand2_2 _07471_ (.A(net4),
    .B(net34),
    .Y(_01332_));
 sky130_fd_sc_hd__or2_1 _07472_ (.A(_01200_),
    .B(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__a22o_1 _07473_ (.A1(net4),
    .A2(net34),
    .B1(net64),
    .B2(net5),
    .X(_01334_));
 sky130_fd_sc_hd__nand4_1 _07474_ (.A(_01333_),
    .B(_01334_),
    .C(net35),
    .D(net3),
    .Y(_01335_));
 sky130_fd_sc_hd__o21ai_1 _07475_ (.A1(_01200_),
    .A2(_01332_),
    .B1(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__a22o_1 _07476_ (.A1(net4),
    .A2(net35),
    .B1(_01201_),
    .B2(_01202_),
    .X(_01337_));
 sky130_fd_sc_hd__and3_1 _07477_ (.A(_01203_),
    .B(_01336_),
    .C(_01337_),
    .X(_01338_));
 sky130_fd_sc_hd__nand3_1 _07478_ (.A(_01203_),
    .B(_01336_),
    .C(_01337_),
    .Y(_01339_));
 sky130_fd_sc_hd__a22o_1 _07479_ (.A1(net38),
    .A2(net32),
    .B1(_01223_),
    .B2(_01224_),
    .X(_01341_));
 sky130_fd_sc_hd__a21o_1 _07480_ (.A1(_01203_),
    .A2(_01337_),
    .B1(_01336_),
    .X(_01342_));
 sky130_fd_sc_hd__a31o_1 _07481_ (.A1(_01225_),
    .A2(_01341_),
    .A3(_01342_),
    .B1(_01338_),
    .X(_01343_));
 sky130_fd_sc_hd__a21bo_1 _07482_ (.A1(_01320_),
    .A2(_01323_),
    .B1_N(_01324_),
    .X(_01344_));
 sky130_fd_sc_hd__a22o_1 _07483_ (.A1(_01083_),
    .A2(_01207_),
    .B1(_01209_),
    .B2(_01206_),
    .X(_01345_));
 sky130_fd_sc_hd__a21oi_1 _07484_ (.A1(_01210_),
    .A2(_01345_),
    .B1(_01344_),
    .Y(_01346_));
 sky130_fd_sc_hd__and3_1 _07485_ (.A(_01210_),
    .B(_01344_),
    .C(_01345_),
    .X(_01347_));
 sky130_fd_sc_hd__nor2_1 _07486_ (.A(_01346_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__xnor2_1 _07487_ (.A(_01343_),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__a21oi_1 _07488_ (.A1(_01196_),
    .A2(_01330_),
    .B1(_01328_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor3_1 _07489_ (.A(_01349_),
    .B(_01350_),
    .C(_01331_),
    .Y(_01352_));
 sky130_fd_sc_hd__a31o_1 _07490_ (.A1(_01196_),
    .A2(_01328_),
    .A3(_01330_),
    .B1(_01352_),
    .X(_01353_));
 sky130_fd_sc_hd__or3b_1 _07491_ (.A(_01217_),
    .B(_01294_),
    .C_N(_01353_),
    .X(_01354_));
 sky130_fd_sc_hd__nand4_2 _07492_ (.A(net37),
    .B(net36),
    .C(net2),
    .D(net32),
    .Y(_01355_));
 sky130_fd_sc_hd__a22o_1 _07493_ (.A1(net36),
    .A2(net2),
    .B1(net32),
    .B2(net37),
    .X(_01356_));
 sky130_fd_sc_hd__nand4_2 _07494_ (.A(_01356_),
    .B(net31),
    .C(net38),
    .D(_01355_),
    .Y(_01357_));
 sky130_fd_sc_hd__nand2_1 _07495_ (.A(_01355_),
    .B(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__a22o_1 _07496_ (.A1(net41),
    .A2(net29),
    .B1(_01229_),
    .B2(_01231_),
    .X(_01359_));
 sky130_fd_sc_hd__nand3_1 _07497_ (.A(_01232_),
    .B(_01358_),
    .C(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand4_1 _07498_ (.A(net40),
    .B(net39),
    .C(net30),
    .D(net29),
    .Y(_01361_));
 sky130_fd_sc_hd__a22o_1 _07499_ (.A1(net39),
    .A2(net30),
    .B1(net29),
    .B2(net40),
    .X(_01363_));
 sky130_fd_sc_hd__nand4_1 _07500_ (.A(_01363_),
    .B(net28),
    .C(net41),
    .D(_01361_),
    .Y(_01364_));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(_01361_),
    .B(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__a21o_1 _07502_ (.A1(_01232_),
    .A2(_01359_),
    .B1(_01358_),
    .X(_01366_));
 sky130_fd_sc_hd__nand3_1 _07503_ (.A(_01360_),
    .B(_01365_),
    .C(_01366_),
    .Y(_01367_));
 sky130_fd_sc_hd__a311o_1 _07504_ (.A1(net41),
    .A2(_01231_),
    .A3(net29),
    .B1(_01228_),
    .C1(_01234_),
    .X(_01368_));
 sky130_fd_sc_hd__nand2_1 _07505_ (.A(_01235_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__a21oi_1 _07506_ (.A1(_01360_),
    .A2(_01367_),
    .B1(_01369_),
    .Y(_01370_));
 sky130_fd_sc_hd__nand4_1 _07507_ (.A(net43),
    .B(net42),
    .C(net28),
    .D(net27),
    .Y(_01371_));
 sky130_fd_sc_hd__a22o_1 _07508_ (.A1(net42),
    .A2(net28),
    .B1(net27),
    .B2(net43),
    .X(_01372_));
 sky130_fd_sc_hd__nand4_1 _07509_ (.A(_01372_),
    .B(net26),
    .C(net45),
    .D(_01371_),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _07510_ (.A(_01371_),
    .B(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__a22o_1 _07511_ (.A1(net45),
    .A2(net27),
    .B1(_01240_),
    .B2(_01242_),
    .X(_01376_));
 sky130_fd_sc_hd__a21oi_1 _07512_ (.A1(_01243_),
    .A2(_01376_),
    .B1(_01375_),
    .Y(_01377_));
 sky130_fd_sc_hd__and3_1 _07513_ (.A(_01243_),
    .B(_01375_),
    .C(_01376_),
    .X(_01378_));
 sky130_fd_sc_hd__nor2_1 _07514_ (.A(_01377_),
    .B(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__and4_1 _07515_ (.A(net46),
    .B(net47),
    .C(net26),
    .D(net23),
    .X(_01380_));
 sky130_fd_sc_hd__a22oi_1 _07516_ (.A1(net46),
    .A2(net26),
    .B1(net23),
    .B2(net47),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _07517_ (.A(_01380_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__xor2_1 _07518_ (.A(_01241_),
    .B(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__xor2_1 _07519_ (.A(_01379_),
    .B(_01383_),
    .X(_01385_));
 sky130_fd_sc_hd__and3_1 _07520_ (.A(_01360_),
    .B(_01367_),
    .C(_01369_),
    .X(_01386_));
 sky130_fd_sc_hd__nor3_1 _07521_ (.A(_01370_),
    .B(_01385_),
    .C(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_1 _07522_ (.A(_01370_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__a21oi_2 _07523_ (.A1(_01348_),
    .A2(_01343_),
    .B1(_01347_),
    .Y(_01389_));
 sky130_fd_sc_hd__o21a_1 _07524_ (.A1(_01254_),
    .A2(_01255_),
    .B1(_01256_),
    .X(_01390_));
 sky130_fd_sc_hd__nor2_1 _07525_ (.A(_01257_),
    .B(_01390_),
    .Y(_01391_));
 sky130_fd_sc_hd__xnor2_1 _07526_ (.A(_01389_),
    .B(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__o21ai_1 _07527_ (.A1(_01370_),
    .A2(_01387_),
    .B1(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__xnor2_2 _07528_ (.A(_01388_),
    .B(_01392_),
    .Y(_01394_));
 sky130_fd_sc_hd__xnor2_2 _07529_ (.A(_01295_),
    .B(_01353_),
    .Y(_01396_));
 sky130_fd_sc_hd__a21boi_1 _07530_ (.A1(_01394_),
    .A2(_01396_),
    .B1_N(_01354_),
    .Y(_01397_));
 sky130_fd_sc_hd__and2_1 _07531_ (.A(_01267_),
    .B(_01269_),
    .X(_01398_));
 sky130_fd_sc_hd__or2_1 _07532_ (.A(_01270_),
    .B(_01398_),
    .X(_01399_));
 sky130_fd_sc_hd__xor2_1 _07533_ (.A(_01397_),
    .B(_01399_),
    .X(_01400_));
 sky130_fd_sc_hd__a41o_1 _07534_ (.A1(net46),
    .A2(net47),
    .A3(net27),
    .A4(net26),
    .B1(_01250_),
    .X(_01401_));
 sky130_fd_sc_hd__or2_1 _07535_ (.A(_01246_),
    .B(_01255_),
    .X(_01402_));
 sky130_fd_sc_hd__o31ai_2 _07536_ (.A1(_01257_),
    .A2(_01389_),
    .A3(_01390_),
    .B1(_01393_),
    .Y(_01403_));
 sky130_fd_sc_hd__xor2_1 _07537_ (.A(_01402_),
    .B(_01403_),
    .X(_01404_));
 sky130_fd_sc_hd__xnor2_1 _07538_ (.A(_01401_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__inv_2 _07539_ (.A(_01405_),
    .Y(_01407_));
 sky130_fd_sc_hd__o2bb2a_1 _07540_ (.A1_N(_01400_),
    .A2_N(_01407_),
    .B1(_01397_),
    .B2(_01399_),
    .X(_01408_));
 sky130_fd_sc_hd__xnor2_1 _07541_ (.A(_01273_),
    .B(_01279_),
    .Y(_01409_));
 sky130_fd_sc_hd__or2_1 _07542_ (.A(_01408_),
    .B(_01409_),
    .X(_01410_));
 sky130_fd_sc_hd__a22oi_2 _07543_ (.A1(_01402_),
    .A2(_01403_),
    .B1(_01404_),
    .B2(_01401_),
    .Y(_01411_));
 sky130_fd_sc_hd__nand2_1 _07544_ (.A(_01409_),
    .B(_01408_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _07545_ (.A(_01410_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__o21ai_1 _07546_ (.A1(_01411_),
    .A2(_01413_),
    .B1(_01410_),
    .Y(_01414_));
 sky130_fd_sc_hd__nand2_1 _07547_ (.A(_01287_),
    .B(_01284_),
    .Y(_01415_));
 sky130_fd_sc_hd__and2_1 _07548_ (.A(_01288_),
    .B(_01415_),
    .X(_01416_));
 sky130_fd_sc_hd__and2_1 _07549_ (.A(_01416_),
    .B(_01414_),
    .X(_01418_));
 sky130_fd_sc_hd__xnor2_1 _07550_ (.A(_01414_),
    .B(_01416_),
    .Y(_01419_));
 sky130_fd_sc_hd__xnor2_1 _07551_ (.A(_01400_),
    .B(_01405_),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _07552_ (.A(net11),
    .B(net33),
    .Y(_01421_));
 sky130_fd_sc_hd__or2_1 _07553_ (.A(_01297_),
    .B(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__a22o_1 _07554_ (.A1(net11),
    .A2(net44),
    .B1(net33),
    .B2(net13),
    .X(_01423_));
 sky130_fd_sc_hd__o2111ai_4 _07555_ (.A1(_01297_),
    .A2(_01421_),
    .B1(net10),
    .C1(net55),
    .D1(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__o21ai_1 _07556_ (.A1(_01297_),
    .A2(_01421_),
    .B1(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__a22o_1 _07557_ (.A1(net11),
    .A2(net55),
    .B1(_01298_),
    .B2(_01299_),
    .X(_01426_));
 sky130_fd_sc_hd__nand3_2 _07558_ (.A(_01300_),
    .B(_01425_),
    .C(_01426_),
    .Y(_01427_));
 sky130_fd_sc_hd__a22o_1 _07559_ (.A1(net9),
    .A2(net59),
    .B1(net58),
    .B2(net10),
    .X(_01429_));
 sky130_fd_sc_hd__nand4_1 _07560_ (.A(net10),
    .B(net9),
    .C(net59),
    .D(net58),
    .Y(_01430_));
 sky130_fd_sc_hd__nand4_1 _07561_ (.A(_01429_),
    .B(_01430_),
    .C(net8),
    .D(net60),
    .Y(_01431_));
 sky130_fd_sc_hd__a22o_1 _07562_ (.A1(net8),
    .A2(net60),
    .B1(_01429_),
    .B2(_01430_),
    .X(_01432_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(_01431_),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__a21o_1 _07564_ (.A1(_01300_),
    .A2(_01426_),
    .B1(_01425_),
    .X(_01434_));
 sky130_fd_sc_hd__nand4_1 _07565_ (.A(_01427_),
    .B(_01431_),
    .C(_01432_),
    .D(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__a21o_1 _07566_ (.A1(_01304_),
    .A2(_01311_),
    .B1(_01310_),
    .X(_01436_));
 sky130_fd_sc_hd__nand3_1 _07567_ (.A(_01304_),
    .B(_01310_),
    .C(_01311_),
    .Y(_01437_));
 sky130_fd_sc_hd__a22o_1 _07568_ (.A1(_01427_),
    .A2(_01435_),
    .B1(_01436_),
    .B2(_01437_),
    .X(_01438_));
 sky130_fd_sc_hd__nand4_2 _07569_ (.A(net7),
    .B(net6),
    .C(net62),
    .D(net61),
    .Y(_01440_));
 sky130_fd_sc_hd__a22o_1 _07570_ (.A1(net6),
    .A2(net62),
    .B1(net61),
    .B2(net7),
    .X(_01441_));
 sky130_fd_sc_hd__nand4_2 _07571_ (.A(_01441_),
    .B(net63),
    .C(net5),
    .D(_01440_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _07572_ (.A(_01440_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _07573_ (.A(_01430_),
    .B(_01431_),
    .Y(_01444_));
 sky130_fd_sc_hd__a22o_1 _07574_ (.A1(net6),
    .A2(net63),
    .B1(_01316_),
    .B2(_01317_),
    .X(_01445_));
 sky130_fd_sc_hd__a21o_1 _07575_ (.A1(_01319_),
    .A2(_01445_),
    .B1(_01444_),
    .X(_01446_));
 sky130_fd_sc_hd__nand3_1 _07576_ (.A(_01319_),
    .B(_01444_),
    .C(_01445_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand3_1 _07577_ (.A(_01443_),
    .B(_01446_),
    .C(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__a21o_1 _07578_ (.A1(_01446_),
    .A2(_01447_),
    .B1(_01443_),
    .X(_01449_));
 sky130_fd_sc_hd__nand2_1 _07579_ (.A(_01448_),
    .B(_01449_),
    .Y(_01451_));
 sky130_fd_sc_hd__nand4_1 _07580_ (.A(_01427_),
    .B(_01435_),
    .C(_01436_),
    .D(_01437_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand4_1 _07581_ (.A(_01438_),
    .B(_01448_),
    .C(_01449_),
    .D(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__a211o_1 _07582_ (.A1(_01314_),
    .A2(_01315_),
    .B1(_01325_),
    .C1(_01326_),
    .X(_01454_));
 sky130_fd_sc_hd__nand2b_1 _07583_ (.A_N(_01327_),
    .B(_01454_),
    .Y(_01455_));
 sky130_fd_sc_hd__a21o_1 _07584_ (.A1(_01438_),
    .A2(_01453_),
    .B1(_01455_),
    .X(_01456_));
 sky130_fd_sc_hd__nand3_1 _07585_ (.A(_01438_),
    .B(_01453_),
    .C(_01455_),
    .Y(_01457_));
 sky130_fd_sc_hd__nand2_1 _07586_ (.A(net3),
    .B(net64),
    .Y(_01458_));
 sky130_fd_sc_hd__or2_1 _07587_ (.A(_01332_),
    .B(_01458_),
    .X(_01459_));
 sky130_fd_sc_hd__a22o_1 _07588_ (.A1(net3),
    .A2(net34),
    .B1(net64),
    .B2(net4),
    .X(_01460_));
 sky130_fd_sc_hd__o2111ai_4 _07589_ (.A1(_01332_),
    .A2(_01458_),
    .B1(net35),
    .C1(net2),
    .D1(_01460_),
    .Y(_01462_));
 sky130_fd_sc_hd__o21ai_1 _07590_ (.A1(_01332_),
    .A2(_01458_),
    .B1(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__a22o_1 _07591_ (.A1(net35),
    .A2(net3),
    .B1(_01333_),
    .B2(_01334_),
    .X(_01464_));
 sky130_fd_sc_hd__nand3_1 _07592_ (.A(_01335_),
    .B(_01463_),
    .C(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__a22o_1 _07593_ (.A1(net38),
    .A2(net31),
    .B1(_01355_),
    .B2(_01356_),
    .X(_01466_));
 sky130_fd_sc_hd__a21o_1 _07594_ (.A1(_01335_),
    .A2(_01464_),
    .B1(_01463_),
    .X(_01467_));
 sky130_fd_sc_hd__nand4_2 _07595_ (.A(_01357_),
    .B(_01465_),
    .C(_01466_),
    .D(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _07596_ (.A(_01465_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__and2_1 _07597_ (.A(_01447_),
    .B(_01448_),
    .X(_01470_));
 sky130_fd_sc_hd__a22oi_1 _07598_ (.A1(_01225_),
    .A2(_01341_),
    .B1(_01342_),
    .B2(_01339_),
    .Y(_01471_));
 sky130_fd_sc_hd__a41o_1 _07599_ (.A1(_01225_),
    .A2(_01339_),
    .A3(_01341_),
    .A4(_01342_),
    .B1(_01471_),
    .X(_01473_));
 sky130_fd_sc_hd__xor2_1 _07600_ (.A(_01470_),
    .B(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__nand2_1 _07601_ (.A(_01474_),
    .B(_01469_),
    .Y(_01475_));
 sky130_fd_sc_hd__or2_1 _07602_ (.A(_01469_),
    .B(_01474_),
    .X(_01476_));
 sky130_fd_sc_hd__nand4_2 _07603_ (.A(_01456_),
    .B(_01457_),
    .C(_01475_),
    .D(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__o21a_1 _07604_ (.A1(_01331_),
    .A2(_01350_),
    .B1(_01349_),
    .X(_01478_));
 sky130_fd_sc_hd__or2_1 _07605_ (.A(_01352_),
    .B(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__a21oi_1 _07606_ (.A1(_01456_),
    .A2(_01477_),
    .B1(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nand4_2 _07607_ (.A(net37),
    .B(net36),
    .C(net32),
    .D(net31),
    .Y(_01481_));
 sky130_fd_sc_hd__a22o_1 _07608_ (.A1(net36),
    .A2(net32),
    .B1(net31),
    .B2(net37),
    .X(_01482_));
 sky130_fd_sc_hd__nand4_2 _07609_ (.A(_01482_),
    .B(net30),
    .C(net38),
    .D(_01481_),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(_01481_),
    .B(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__a22o_1 _07611_ (.A1(net41),
    .A2(net28),
    .B1(_01361_),
    .B2(_01363_),
    .X(_01486_));
 sky130_fd_sc_hd__nand3_1 _07612_ (.A(_01364_),
    .B(_01485_),
    .C(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand4_1 _07613_ (.A(net40),
    .B(net39),
    .C(net29),
    .D(net28),
    .Y(_01488_));
 sky130_fd_sc_hd__a22o_1 _07614_ (.A1(net39),
    .A2(net29),
    .B1(net28),
    .B2(net40),
    .X(_01489_));
 sky130_fd_sc_hd__nand4_1 _07615_ (.A(_01489_),
    .B(net27),
    .C(net41),
    .D(_01488_),
    .Y(_01490_));
 sky130_fd_sc_hd__nand2_1 _07616_ (.A(_01488_),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__a21o_1 _07617_ (.A1(_01364_),
    .A2(_01486_),
    .B1(_01485_),
    .X(_01492_));
 sky130_fd_sc_hd__nand3_1 _07618_ (.A(_01487_),
    .B(_01491_),
    .C(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand2_1 _07619_ (.A(_01487_),
    .B(_01493_),
    .Y(_01495_));
 sky130_fd_sc_hd__a21o_1 _07620_ (.A1(_01360_),
    .A2(_01366_),
    .B1(_01365_),
    .X(_01496_));
 sky130_fd_sc_hd__nand3_1 _07621_ (.A(_01367_),
    .B(_01495_),
    .C(_01496_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand4_2 _07622_ (.A(net43),
    .B(net42),
    .C(net27),
    .D(net26),
    .Y(_01498_));
 sky130_fd_sc_hd__a22o_1 _07623_ (.A1(net42),
    .A2(net27),
    .B1(net26),
    .B2(net43),
    .X(_01499_));
 sky130_fd_sc_hd__nand4_2 _07624_ (.A(_01499_),
    .B(net23),
    .C(net45),
    .D(_01498_),
    .Y(_01500_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(_01498_),
    .B(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__a22o_1 _07626_ (.A1(net45),
    .A2(net26),
    .B1(_01371_),
    .B2(_01372_),
    .X(_01502_));
 sky130_fd_sc_hd__a21o_1 _07627_ (.A1(_01374_),
    .A2(_01502_),
    .B1(_01501_),
    .X(_01503_));
 sky130_fd_sc_hd__nand3_1 _07628_ (.A(_01374_),
    .B(_01501_),
    .C(_01502_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _07629_ (.A(_01503_),
    .B(_01504_),
    .Y(_01506_));
 sky130_fd_sc_hd__and4_1 _07630_ (.A(net46),
    .B(net47),
    .C(net23),
    .D(net12),
    .X(_01507_));
 sky130_fd_sc_hd__o2bb2a_1 _07631_ (.A1_N(net46),
    .A2_N(net23),
    .B1(_01241_),
    .B2(_01043_),
    .X(_01508_));
 sky130_fd_sc_hd__nor3_1 _07632_ (.A(_01263_),
    .B(_01507_),
    .C(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__o21a_1 _07633_ (.A1(_01507_),
    .A2(_01508_),
    .B1(_01263_),
    .X(_01510_));
 sky130_fd_sc_hd__nor2_1 _07634_ (.A(_01509_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__xor2_1 _07635_ (.A(_01506_),
    .B(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__a21o_1 _07636_ (.A1(_01367_),
    .A2(_01496_),
    .B1(_01495_),
    .X(_01513_));
 sky130_fd_sc_hd__nand2_1 _07637_ (.A(_01497_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__o21ai_1 _07638_ (.A1(_01512_),
    .A2(_01514_),
    .B1(_01497_),
    .Y(_01515_));
 sky130_fd_sc_hd__o21ai_1 _07639_ (.A1(_01470_),
    .A2(_01473_),
    .B1(_01475_),
    .Y(_01517_));
 sky130_fd_sc_hd__o21a_1 _07640_ (.A1(_01370_),
    .A2(_01386_),
    .B1(_01385_),
    .X(_01518_));
 sky130_fd_sc_hd__or2_1 _07641_ (.A(_01387_),
    .B(_01518_),
    .X(_01519_));
 sky130_fd_sc_hd__and2b_1 _07642_ (.A_N(_01519_),
    .B(_01517_),
    .X(_01520_));
 sky130_fd_sc_hd__xnor2_1 _07643_ (.A(_01517_),
    .B(_01519_),
    .Y(_01521_));
 sky130_fd_sc_hd__xnor2_1 _07644_ (.A(_01515_),
    .B(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__and3_1 _07645_ (.A(_01456_),
    .B(_01477_),
    .C(_01479_),
    .X(_01523_));
 sky130_fd_sc_hd__nor2_1 _07646_ (.A(_01480_),
    .B(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__and2b_1 _07647_ (.A_N(_01522_),
    .B(_01524_),
    .X(_01525_));
 sky130_fd_sc_hd__nor2_1 _07648_ (.A(_01480_),
    .B(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__xnor2_2 _07649_ (.A(_01394_),
    .B(_01396_),
    .Y(_01528_));
 sky130_fd_sc_hd__xnor2_1 _07650_ (.A(_01526_),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__a21o_1 _07651_ (.A1(net12),
    .A2(_01382_),
    .B1(_01380_),
    .X(_01530_));
 sky130_fd_sc_hd__o21ba_1 _07652_ (.A1(_01377_),
    .A2(_01383_),
    .B1_N(_01378_),
    .X(_01531_));
 sky130_fd_sc_hd__a21oi_1 _07653_ (.A1(_01521_),
    .A2(_01515_),
    .B1(_01520_),
    .Y(_01532_));
 sky130_fd_sc_hd__xor2_1 _07654_ (.A(_01531_),
    .B(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__xnor2_1 _07655_ (.A(_01530_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__o22ai_2 _07656_ (.A1(_01528_),
    .A2(_01526_),
    .B1(_01534_),
    .B2(_01529_),
    .Y(_01535_));
 sky130_fd_sc_hd__o2bb2a_1 _07657_ (.A1_N(_01530_),
    .A2_N(_01533_),
    .B1(_01532_),
    .B2(_01531_),
    .X(_01536_));
 sky130_fd_sc_hd__xor2_1 _07658_ (.A(_01420_),
    .B(_01535_),
    .X(_01537_));
 sky130_fd_sc_hd__and2b_1 _07659_ (.A_N(_01536_),
    .B(_01537_),
    .X(_01539_));
 sky130_fd_sc_hd__a21o_1 _07660_ (.A1(_01420_),
    .A2(_01535_),
    .B1(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__xnor2_1 _07661_ (.A(_01411_),
    .B(_01413_),
    .Y(_01541_));
 sky130_fd_sc_hd__and2b_1 _07662_ (.A_N(_01541_),
    .B(_01540_),
    .X(_01542_));
 sky130_fd_sc_hd__and4_1 _07663_ (.A(net11),
    .B(net10),
    .C(net44),
    .D(net33),
    .X(_01543_));
 sky130_fd_sc_hd__nand4_1 _07664_ (.A(net11),
    .B(net10),
    .C(net44),
    .D(net33),
    .Y(_01544_));
 sky130_fd_sc_hd__a22o_1 _07665_ (.A1(net10),
    .A2(net44),
    .B1(net33),
    .B2(net11),
    .X(_01545_));
 sky130_fd_sc_hd__nand4_1 _07666_ (.A(_01545_),
    .B(net55),
    .C(net9),
    .D(_01544_),
    .Y(_01546_));
 sky130_fd_sc_hd__a31o_1 _07667_ (.A1(_01545_),
    .A2(net55),
    .A3(net9),
    .B1(_01543_),
    .X(_01547_));
 sky130_fd_sc_hd__a22o_1 _07668_ (.A1(net10),
    .A2(net55),
    .B1(_01422_),
    .B2(_01423_),
    .X(_01548_));
 sky130_fd_sc_hd__nand3_2 _07669_ (.A(_01424_),
    .B(_01547_),
    .C(_01548_),
    .Y(_01550_));
 sky130_fd_sc_hd__a22o_1 _07670_ (.A1(net8),
    .A2(net59),
    .B1(net58),
    .B2(net9),
    .X(_01551_));
 sky130_fd_sc_hd__nand4_2 _07671_ (.A(net9),
    .B(net8),
    .C(net59),
    .D(net58),
    .Y(_01552_));
 sky130_fd_sc_hd__nand4_2 _07672_ (.A(_01551_),
    .B(_01552_),
    .C(net7),
    .D(net60),
    .Y(_01553_));
 sky130_fd_sc_hd__a22o_1 _07673_ (.A1(net7),
    .A2(net60),
    .B1(_01551_),
    .B2(_01552_),
    .X(_01554_));
 sky130_fd_sc_hd__a21o_1 _07674_ (.A1(_01424_),
    .A2(_01548_),
    .B1(_01547_),
    .X(_01555_));
 sky130_fd_sc_hd__nand4_2 _07675_ (.A(_01550_),
    .B(_01553_),
    .C(_01554_),
    .D(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__a21o_1 _07676_ (.A1(_01427_),
    .A2(_01434_),
    .B1(_01433_),
    .X(_01557_));
 sky130_fd_sc_hd__nand3_1 _07677_ (.A(_01427_),
    .B(_01433_),
    .C(_01434_),
    .Y(_01558_));
 sky130_fd_sc_hd__a22o_1 _07678_ (.A1(_01550_),
    .A2(_01556_),
    .B1(_01557_),
    .B2(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__nand4_2 _07679_ (.A(net6),
    .B(net5),
    .C(net62),
    .D(net61),
    .Y(_01561_));
 sky130_fd_sc_hd__a22o_1 _07680_ (.A1(net5),
    .A2(net62),
    .B1(net61),
    .B2(net6),
    .X(_01562_));
 sky130_fd_sc_hd__nand4_2 _07681_ (.A(_01562_),
    .B(net63),
    .C(net4),
    .D(_01561_),
    .Y(_01563_));
 sky130_fd_sc_hd__nand2_1 _07682_ (.A(_01561_),
    .B(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__nand2_1 _07683_ (.A(_01552_),
    .B(_01553_),
    .Y(_01565_));
 sky130_fd_sc_hd__a22o_1 _07684_ (.A1(net5),
    .A2(net63),
    .B1(_01440_),
    .B2(_01441_),
    .X(_01566_));
 sky130_fd_sc_hd__a21o_1 _07685_ (.A1(_01442_),
    .A2(_01566_),
    .B1(_01565_),
    .X(_01567_));
 sky130_fd_sc_hd__nand3_1 _07686_ (.A(_01442_),
    .B(_01565_),
    .C(_01566_),
    .Y(_01568_));
 sky130_fd_sc_hd__and3_1 _07687_ (.A(_01564_),
    .B(_01567_),
    .C(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__a21oi_1 _07688_ (.A1(_01567_),
    .A2(_01568_),
    .B1(_01564_),
    .Y(_01570_));
 sky130_fd_sc_hd__nor2_1 _07689_ (.A(_01569_),
    .B(_01570_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand4_1 _07690_ (.A(_01550_),
    .B(_01556_),
    .C(_01557_),
    .D(_01558_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand3_1 _07691_ (.A(_01559_),
    .B(_01572_),
    .C(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__a21o_1 _07692_ (.A1(_01438_),
    .A2(_01452_),
    .B1(_01451_),
    .X(_01575_));
 sky130_fd_sc_hd__nand3_1 _07693_ (.A(_01438_),
    .B(_01451_),
    .C(_01452_),
    .Y(_01576_));
 sky130_fd_sc_hd__a22oi_2 _07694_ (.A1(_01559_),
    .A2(_01574_),
    .B1(_01575_),
    .B2(_01576_),
    .Y(_01577_));
 sky130_fd_sc_hd__and4_1 _07695_ (.A(net3),
    .B(net34),
    .C(net2),
    .D(net64),
    .X(_01578_));
 sky130_fd_sc_hd__nand4_1 _07696_ (.A(net3),
    .B(net34),
    .C(net2),
    .D(net64),
    .Y(_01579_));
 sky130_fd_sc_hd__a22o_1 _07697_ (.A1(net34),
    .A2(net2),
    .B1(net64),
    .B2(net3),
    .X(_01580_));
 sky130_fd_sc_hd__and4_2 _07698_ (.A(_01580_),
    .B(net32),
    .C(net35),
    .D(_01579_),
    .X(_01581_));
 sky130_fd_sc_hd__a22o_1 _07699_ (.A1(net35),
    .A2(net2),
    .B1(_01459_),
    .B2(_01460_),
    .X(_01583_));
 sky130_fd_sc_hd__o211ai_4 _07700_ (.A1(_01578_),
    .A2(_01581_),
    .B1(_01583_),
    .C1(_01462_),
    .Y(_01584_));
 sky130_fd_sc_hd__a22o_1 _07701_ (.A1(net38),
    .A2(net30),
    .B1(_01481_),
    .B2(_01482_),
    .X(_01585_));
 sky130_fd_sc_hd__a211o_1 _07702_ (.A1(_01462_),
    .A2(_01583_),
    .B1(_01581_),
    .C1(_01578_),
    .X(_01586_));
 sky130_fd_sc_hd__nand4_2 _07703_ (.A(_01484_),
    .B(_01584_),
    .C(_01585_),
    .D(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__a31o_1 _07704_ (.A1(_01442_),
    .A2(_01565_),
    .A3(_01566_),
    .B1(_01569_),
    .X(_01588_));
 sky130_fd_sc_hd__a22o_1 _07705_ (.A1(_01357_),
    .A2(_01466_),
    .B1(_01467_),
    .B2(_01465_),
    .X(_01589_));
 sky130_fd_sc_hd__a21oi_1 _07706_ (.A1(_01468_),
    .A2(_01589_),
    .B1(_01588_),
    .Y(_01590_));
 sky130_fd_sc_hd__and3_1 _07707_ (.A(_01468_),
    .B(_01588_),
    .C(_01589_),
    .X(_01591_));
 sky130_fd_sc_hd__a211oi_2 _07708_ (.A1(_01584_),
    .A2(_01587_),
    .B1(_01590_),
    .C1(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__o211a_1 _07709_ (.A1(_01590_),
    .A2(_01591_),
    .B1(_01584_),
    .C1(_01587_),
    .X(_01594_));
 sky130_fd_sc_hd__nor2_1 _07710_ (.A(_01592_),
    .B(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__and4_1 _07711_ (.A(_01559_),
    .B(_01574_),
    .C(_01575_),
    .D(_01576_),
    .X(_01596_));
 sky130_fd_sc_hd__nor2_1 _07712_ (.A(_01577_),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__a21o_1 _07713_ (.A1(_01595_),
    .A2(_01597_),
    .B1(_01577_),
    .X(_01598_));
 sky130_fd_sc_hd__a22o_1 _07714_ (.A1(_01456_),
    .A2(_01457_),
    .B1(_01475_),
    .B2(_01476_),
    .X(_01599_));
 sky130_fd_sc_hd__nand2_1 _07715_ (.A(_01477_),
    .B(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__nand3_1 _07716_ (.A(_01477_),
    .B(_01598_),
    .C(_01599_),
    .Y(_01601_));
 sky130_fd_sc_hd__xnor2_1 _07717_ (.A(_01598_),
    .B(_01600_),
    .Y(_01602_));
 sky130_fd_sc_hd__and4_1 _07718_ (.A(net37),
    .B(net36),
    .C(net31),
    .D(net30),
    .X(_01603_));
 sky130_fd_sc_hd__nand4_1 _07719_ (.A(net37),
    .B(net36),
    .C(net31),
    .D(net30),
    .Y(_01605_));
 sky130_fd_sc_hd__a22o_1 _07720_ (.A1(net36),
    .A2(net31),
    .B1(net30),
    .B2(net37),
    .X(_01606_));
 sky130_fd_sc_hd__or4b_1 _07721_ (.A(_01087_),
    .B(_01186_),
    .C(_01603_),
    .D_N(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__a31o_1 _07722_ (.A1(_01606_),
    .A2(net29),
    .A3(net38),
    .B1(_01603_),
    .X(_01608_));
 sky130_fd_sc_hd__a22o_1 _07723_ (.A1(net41),
    .A2(net27),
    .B1(_01488_),
    .B2(_01489_),
    .X(_01609_));
 sky130_fd_sc_hd__nand3_1 _07724_ (.A(_01490_),
    .B(_01608_),
    .C(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__nand4_2 _07725_ (.A(net40),
    .B(net39),
    .C(net28),
    .D(net27),
    .Y(_01611_));
 sky130_fd_sc_hd__a22o_1 _07726_ (.A1(net39),
    .A2(net28),
    .B1(net27),
    .B2(net40),
    .X(_01612_));
 sky130_fd_sc_hd__nand4_2 _07727_ (.A(_01612_),
    .B(net26),
    .C(net41),
    .D(_01611_),
    .Y(_01613_));
 sky130_fd_sc_hd__nand2_1 _07728_ (.A(_01611_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__a21o_1 _07729_ (.A1(_01490_),
    .A2(_01609_),
    .B1(_01608_),
    .X(_01616_));
 sky130_fd_sc_hd__nand3_1 _07730_ (.A(_01610_),
    .B(_01614_),
    .C(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand2_1 _07731_ (.A(_01610_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__a21o_1 _07732_ (.A1(_01487_),
    .A2(_01492_),
    .B1(_01491_),
    .X(_01619_));
 sky130_fd_sc_hd__nand3_1 _07733_ (.A(_01493_),
    .B(_01618_),
    .C(_01619_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand4_1 _07734_ (.A(net43),
    .B(net42),
    .C(net26),
    .D(net23),
    .Y(_01621_));
 sky130_fd_sc_hd__a22o_1 _07735_ (.A1(net42),
    .A2(net26),
    .B1(net23),
    .B2(net43),
    .X(_01622_));
 sky130_fd_sc_hd__nand4_1 _07736_ (.A(_01622_),
    .B(net12),
    .C(net45),
    .D(_01621_),
    .Y(_01623_));
 sky130_fd_sc_hd__nand2_1 _07737_ (.A(_01621_),
    .B(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__a22o_1 _07738_ (.A1(net45),
    .A2(net23),
    .B1(_01498_),
    .B2(_01499_),
    .X(_01625_));
 sky130_fd_sc_hd__a21oi_1 _07739_ (.A1(_01500_),
    .A2(_01625_),
    .B1(_01624_),
    .Y(_01627_));
 sky130_fd_sc_hd__and3_1 _07740_ (.A(_01500_),
    .B(_01624_),
    .C(_01625_),
    .X(_01628_));
 sky130_fd_sc_hd__and4_1 _07741_ (.A(net46),
    .B(net47),
    .C(net12),
    .D(net1),
    .X(_01629_));
 sky130_fd_sc_hd__o2bb2a_1 _07742_ (.A1_N(net46),
    .A2_N(net12),
    .B1(_01263_),
    .B2(_01043_),
    .X(_01630_));
 sky130_fd_sc_hd__o22a_1 _07743_ (.A1(_01627_),
    .A2(_01628_),
    .B1(_01629_),
    .B2(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__nor4_1 _07744_ (.A(_01627_),
    .B(_01628_),
    .C(_01629_),
    .D(_01630_),
    .Y(_01632_));
 sky130_fd_sc_hd__or2_1 _07745_ (.A(_01631_),
    .B(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__a21o_1 _07746_ (.A1(_01493_),
    .A2(_01619_),
    .B1(_01618_),
    .X(_01634_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_01620_),
    .B(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__o21a_1 _07748_ (.A1(_01633_),
    .A2(_01635_),
    .B1(_01620_),
    .X(_01636_));
 sky130_fd_sc_hd__xor2_1 _07749_ (.A(_01512_),
    .B(_01514_),
    .X(_01638_));
 sky130_fd_sc_hd__a311o_1 _07750_ (.A1(_01468_),
    .A2(_01588_),
    .A3(_01589_),
    .B1(_01592_),
    .C1(_01638_),
    .X(_01639_));
 sky130_fd_sc_hd__o21ai_1 _07751_ (.A1(_01591_),
    .A2(_01592_),
    .B1(_01638_),
    .Y(_01640_));
 sky130_fd_sc_hd__nand2_1 _07752_ (.A(_01639_),
    .B(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hd__xor2_1 _07753_ (.A(_01636_),
    .B(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__nand2_1 _07754_ (.A(_01602_),
    .B(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__xor2_1 _07755_ (.A(_01522_),
    .B(_01524_),
    .X(_01644_));
 sky130_fd_sc_hd__a21oi_1 _07756_ (.A1(_01601_),
    .A2(_01643_),
    .B1(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__a41o_1 _07757_ (.A1(net46),
    .A2(net47),
    .A3(net23),
    .A4(net12),
    .B1(_01509_),
    .X(_01646_));
 sky130_fd_sc_hd__o31a_1 _07758_ (.A1(_01509_),
    .A2(_01510_),
    .A3(_01506_),
    .B1(_01504_),
    .X(_01647_));
 sky130_fd_sc_hd__o21ai_1 _07759_ (.A1(_01636_),
    .A2(_01641_),
    .B1(_01640_),
    .Y(_01649_));
 sky130_fd_sc_hd__and2b_1 _07760_ (.A_N(_01647_),
    .B(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__xnor2_1 _07761_ (.A(_01647_),
    .B(_01649_),
    .Y(_01651_));
 sky130_fd_sc_hd__o21a_1 _07762_ (.A1(_01507_),
    .A2(_01509_),
    .B1(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__nor2_1 _07763_ (.A(_01646_),
    .B(_01651_),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _07764_ (.A(_01652_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__nand3_1 _07765_ (.A(_01601_),
    .B(_01643_),
    .C(_01644_),
    .Y(_01655_));
 sky130_fd_sc_hd__and2b_1 _07766_ (.A_N(_01645_),
    .B(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__and2_1 _07767_ (.A(_01654_),
    .B(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__xor2_1 _07768_ (.A(_01529_),
    .B(_01534_),
    .X(_01658_));
 sky130_fd_sc_hd__o21ai_1 _07769_ (.A1(_01645_),
    .A2(_01657_),
    .B1(_01658_),
    .Y(_01660_));
 sky130_fd_sc_hd__or3_1 _07770_ (.A(_01645_),
    .B(_01657_),
    .C(_01658_),
    .X(_01661_));
 sky130_fd_sc_hd__and2_1 _07771_ (.A(_01660_),
    .B(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__o21ai_1 _07772_ (.A1(_01650_),
    .A2(_01652_),
    .B1(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__xor2_1 _07773_ (.A(_01536_),
    .B(_01537_),
    .X(_01664_));
 sky130_fd_sc_hd__a21o_1 _07774_ (.A1(_01660_),
    .A2(_01663_),
    .B1(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__nand3_1 _07775_ (.A(_01660_),
    .B(_01663_),
    .C(_01664_),
    .Y(_01666_));
 sky130_fd_sc_hd__and2_1 _07776_ (.A(_01665_),
    .B(_01666_),
    .X(_01667_));
 sky130_fd_sc_hd__nand4_2 _07777_ (.A(net10),
    .B(net9),
    .C(net44),
    .D(net33),
    .Y(_01668_));
 sky130_fd_sc_hd__a22o_1 _07778_ (.A1(net9),
    .A2(net44),
    .B1(net33),
    .B2(net10),
    .X(_01669_));
 sky130_fd_sc_hd__nand4_2 _07779_ (.A(_01669_),
    .B(net55),
    .C(net8),
    .D(_01668_),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _07780_ (.A(_01668_),
    .B(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__a22o_1 _07781_ (.A1(net9),
    .A2(net55),
    .B1(_01544_),
    .B2(_01545_),
    .X(_01673_));
 sky130_fd_sc_hd__and3_1 _07782_ (.A(_01546_),
    .B(_01672_),
    .C(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__nand3_1 _07783_ (.A(_01546_),
    .B(_01672_),
    .C(_01673_),
    .Y(_01675_));
 sky130_fd_sc_hd__a22o_1 _07784_ (.A1(net7),
    .A2(net59),
    .B1(net58),
    .B2(net8),
    .X(_01676_));
 sky130_fd_sc_hd__nand4_1 _07785_ (.A(net8),
    .B(net7),
    .C(net59),
    .D(net58),
    .Y(_01677_));
 sky130_fd_sc_hd__nand4_1 _07786_ (.A(_01676_),
    .B(_01677_),
    .C(net6),
    .D(net60),
    .Y(_01678_));
 sky130_fd_sc_hd__a22o_1 _07787_ (.A1(net6),
    .A2(net60),
    .B1(_01676_),
    .B2(_01677_),
    .X(_01679_));
 sky130_fd_sc_hd__nand2_1 _07788_ (.A(_01678_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__a21o_1 _07789_ (.A1(_01546_),
    .A2(_01673_),
    .B1(_01672_),
    .X(_01682_));
 sky130_fd_sc_hd__a31o_1 _07790_ (.A1(_01678_),
    .A2(_01679_),
    .A3(_01682_),
    .B1(_01674_),
    .X(_01683_));
 sky130_fd_sc_hd__a22o_1 _07791_ (.A1(_01553_),
    .A2(_01554_),
    .B1(_01555_),
    .B2(_01550_),
    .X(_01684_));
 sky130_fd_sc_hd__nand3_1 _07792_ (.A(_01556_),
    .B(_01683_),
    .C(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__nand4_2 _07793_ (.A(net5),
    .B(net4),
    .C(net62),
    .D(net61),
    .Y(_01686_));
 sky130_fd_sc_hd__a22o_1 _07794_ (.A1(net4),
    .A2(net62),
    .B1(net61),
    .B2(net5),
    .X(_01687_));
 sky130_fd_sc_hd__nand4_2 _07795_ (.A(_01687_),
    .B(net63),
    .C(net3),
    .D(_01686_),
    .Y(_01688_));
 sky130_fd_sc_hd__nand2_1 _07796_ (.A(_01686_),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _07797_ (.A(_01677_),
    .B(_01678_),
    .Y(_01690_));
 sky130_fd_sc_hd__a22o_1 _07798_ (.A1(net4),
    .A2(net63),
    .B1(_01561_),
    .B2(_01562_),
    .X(_01691_));
 sky130_fd_sc_hd__a21o_1 _07799_ (.A1(_01563_),
    .A2(_01691_),
    .B1(_01690_),
    .X(_01693_));
 sky130_fd_sc_hd__and3_1 _07800_ (.A(_01563_),
    .B(_01690_),
    .C(_01691_),
    .X(_01694_));
 sky130_fd_sc_hd__nand3_1 _07801_ (.A(_01563_),
    .B(_01690_),
    .C(_01691_),
    .Y(_01695_));
 sky130_fd_sc_hd__and3_1 _07802_ (.A(_01689_),
    .B(_01693_),
    .C(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__nand3_1 _07803_ (.A(_01689_),
    .B(_01693_),
    .C(_01695_),
    .Y(_01697_));
 sky130_fd_sc_hd__a21o_1 _07804_ (.A1(_01693_),
    .A2(_01695_),
    .B1(_01689_),
    .X(_01698_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(_01697_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__a21o_1 _07806_ (.A1(_01556_),
    .A2(_01684_),
    .B1(_01683_),
    .X(_01700_));
 sky130_fd_sc_hd__and4_1 _07807_ (.A(_01685_),
    .B(_01697_),
    .C(_01698_),
    .D(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__a31o_1 _07808_ (.A1(_01556_),
    .A2(_01683_),
    .A3(_01684_),
    .B1(_01701_),
    .X(_01702_));
 sky130_fd_sc_hd__a2bb2o_1 _07809_ (.A1_N(_01569_),
    .A2_N(_01570_),
    .B1(_01573_),
    .B2(_01559_),
    .X(_01704_));
 sky130_fd_sc_hd__nand3_1 _07810_ (.A(_01574_),
    .B(_01702_),
    .C(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_1 _07811_ (.A(net34),
    .B(net32),
    .Y(_01706_));
 sky130_fd_sc_hd__nand4_2 _07812_ (.A(net34),
    .B(net2),
    .C(net64),
    .D(net32),
    .Y(_01707_));
 sky130_fd_sc_hd__a22o_1 _07813_ (.A1(net2),
    .A2(net64),
    .B1(net32),
    .B2(net34),
    .X(_01708_));
 sky130_fd_sc_hd__nand4_2 _07814_ (.A(_01708_),
    .B(net31),
    .C(net35),
    .D(_01707_),
    .Y(_01709_));
 sky130_fd_sc_hd__a22oi_1 _07815_ (.A1(net35),
    .A2(net32),
    .B1(_01579_),
    .B2(_01580_),
    .Y(_01710_));
 sky130_fd_sc_hd__a211o_1 _07816_ (.A1(_01707_),
    .A2(_01709_),
    .B1(_01710_),
    .C1(_01581_),
    .X(_01711_));
 sky130_fd_sc_hd__a22o_1 _07817_ (.A1(net38),
    .A2(net29),
    .B1(_01605_),
    .B2(_01606_),
    .X(_01712_));
 sky130_fd_sc_hd__o211ai_1 _07818_ (.A1(_01581_),
    .A2(_01710_),
    .B1(_01709_),
    .C1(_01707_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand4_1 _07819_ (.A(_01607_),
    .B(_01711_),
    .C(_01712_),
    .D(_01713_),
    .Y(_01715_));
 sky130_fd_sc_hd__nand2_1 _07820_ (.A(_01711_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__a22o_1 _07821_ (.A1(_01484_),
    .A2(_01585_),
    .B1(_01586_),
    .B2(_01584_),
    .X(_01717_));
 sky130_fd_sc_hd__a221oi_1 _07822_ (.A1(_01689_),
    .A2(_01693_),
    .B1(_01717_),
    .B2(_01587_),
    .C1(_01694_),
    .Y(_01718_));
 sky130_fd_sc_hd__o211a_1 _07823_ (.A1(_01694_),
    .A2(_01696_),
    .B1(_01717_),
    .C1(_01587_),
    .X(_01719_));
 sky130_fd_sc_hd__nor2_1 _07824_ (.A(_01718_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__xor2_1 _07825_ (.A(_01716_),
    .B(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__a21o_1 _07826_ (.A1(_01574_),
    .A2(_01704_),
    .B1(_01702_),
    .X(_01722_));
 sky130_fd_sc_hd__nand3_1 _07827_ (.A(_01721_),
    .B(_01722_),
    .C(_01705_),
    .Y(_01723_));
 sky130_fd_sc_hd__or2_1 _07828_ (.A(_01595_),
    .B(_01597_),
    .X(_01724_));
 sky130_fd_sc_hd__o41ai_1 _07829_ (.A1(_01577_),
    .A2(_01592_),
    .A3(_01594_),
    .A4(_01596_),
    .B1(_01724_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21o_1 _07830_ (.A1(_01705_),
    .A2(_01723_),
    .B1(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__and4_1 _07831_ (.A(net37),
    .B(net36),
    .C(net30),
    .D(net29),
    .X(_01728_));
 sky130_fd_sc_hd__nand4_1 _07832_ (.A(net37),
    .B(net36),
    .C(net30),
    .D(net29),
    .Y(_01729_));
 sky130_fd_sc_hd__a22o_1 _07833_ (.A1(net36),
    .A2(net30),
    .B1(net29),
    .B2(net37),
    .X(_01730_));
 sky130_fd_sc_hd__and4_1 _07834_ (.A(_01730_),
    .B(net28),
    .C(net38),
    .D(_01729_),
    .X(_01731_));
 sky130_fd_sc_hd__a22o_1 _07835_ (.A1(net41),
    .A2(net26),
    .B1(_01611_),
    .B2(_01612_),
    .X(_01732_));
 sky130_fd_sc_hd__o211ai_2 _07836_ (.A1(_01728_),
    .A2(_01731_),
    .B1(_01732_),
    .C1(_01613_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand4_2 _07837_ (.A(net40),
    .B(net39),
    .C(net27),
    .D(net26),
    .Y(_01734_));
 sky130_fd_sc_hd__a22o_1 _07838_ (.A1(net39),
    .A2(net27),
    .B1(net26),
    .B2(net40),
    .X(_01735_));
 sky130_fd_sc_hd__nand4_2 _07839_ (.A(_01735_),
    .B(net23),
    .C(net41),
    .D(_01734_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_1 _07840_ (.A(_01734_),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__a211o_1 _07841_ (.A1(_01613_),
    .A2(_01732_),
    .B1(_01731_),
    .C1(_01728_),
    .X(_01739_));
 sky130_fd_sc_hd__a21bo_1 _07842_ (.A1(_01738_),
    .A2(_01739_),
    .B1_N(_01733_),
    .X(_01740_));
 sky130_fd_sc_hd__a21o_1 _07843_ (.A1(_01610_),
    .A2(_01616_),
    .B1(_01614_),
    .X(_01741_));
 sky130_fd_sc_hd__nand3_1 _07844_ (.A(_01617_),
    .B(_01740_),
    .C(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand4_1 _07845_ (.A(net43),
    .B(net42),
    .C(net23),
    .D(net12),
    .Y(_01743_));
 sky130_fd_sc_hd__a22o_1 _07846_ (.A1(net42),
    .A2(net23),
    .B1(net12),
    .B2(net43),
    .X(_01744_));
 sky130_fd_sc_hd__and4_1 _07847_ (.A(_01744_),
    .B(net1),
    .C(net45),
    .D(_01743_),
    .X(_01745_));
 sky130_fd_sc_hd__a41o_1 _07848_ (.A1(net43),
    .A2(net42),
    .A3(net23),
    .A4(net12),
    .B1(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__a22o_1 _07849_ (.A1(net45),
    .A2(net12),
    .B1(_01621_),
    .B2(_01622_),
    .X(_01748_));
 sky130_fd_sc_hd__a21oi_1 _07850_ (.A1(_01623_),
    .A2(_01748_),
    .B1(_01746_),
    .Y(_01749_));
 sky130_fd_sc_hd__and3_1 _07851_ (.A(_01623_),
    .B(_01746_),
    .C(_01748_),
    .X(_01750_));
 sky130_fd_sc_hd__nor2_1 _07852_ (.A(_01749_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__o2bb2a_1 _07853_ (.A1_N(net46),
    .A2_N(net1),
    .B1(_01749_),
    .B2(_01750_),
    .X(_01752_));
 sky130_fd_sc_hd__and3_1 _07854_ (.A(net46),
    .B(net1),
    .C(_01751_),
    .X(_01753_));
 sky130_fd_sc_hd__or2_1 _07855_ (.A(_01752_),
    .B(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__a21o_1 _07856_ (.A1(_01617_),
    .A2(_01741_),
    .B1(_01740_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _07857_ (.A(_01742_),
    .B(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__or2_1 _07858_ (.A(_01754_),
    .B(_01756_),
    .X(_01757_));
 sky130_fd_sc_hd__a21oi_1 _07859_ (.A1(_01720_),
    .A2(_01716_),
    .B1(_01719_),
    .Y(_01759_));
 sky130_fd_sc_hd__xnor2_1 _07860_ (.A(_01633_),
    .B(_01635_),
    .Y(_01760_));
 sky130_fd_sc_hd__xnor2_1 _07861_ (.A(_01759_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__a21o_1 _07862_ (.A1(_01742_),
    .A2(_01757_),
    .B1(_01761_),
    .X(_01762_));
 sky130_fd_sc_hd__o211ai_1 _07863_ (.A1(_01754_),
    .A2(_01756_),
    .B1(_01761_),
    .C1(_01742_),
    .Y(_01763_));
 sky130_fd_sc_hd__and2_1 _07864_ (.A(_01762_),
    .B(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__nand3_1 _07865_ (.A(_01705_),
    .B(_01723_),
    .C(_01726_),
    .Y(_01765_));
 sky130_fd_sc_hd__and2_1 _07866_ (.A(_01727_),
    .B(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__nand2_1 _07867_ (.A(_01764_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__or2_1 _07868_ (.A(_01602_),
    .B(_01642_),
    .X(_01768_));
 sky130_fd_sc_hd__nand2_1 _07869_ (.A(_01643_),
    .B(_01768_),
    .Y(_01770_));
 sky130_fd_sc_hd__a21o_1 _07870_ (.A1(_01727_),
    .A2(_01767_),
    .B1(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__nand3_1 _07871_ (.A(_01727_),
    .B(_01767_),
    .C(_01770_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _07872_ (.A(_01771_),
    .B(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__a31o_1 _07873_ (.A1(_01500_),
    .A2(_01624_),
    .A3(_01625_),
    .B1(_01632_),
    .X(_01774_));
 sky130_fd_sc_hd__o21ai_1 _07874_ (.A1(_01759_),
    .A2(_01760_),
    .B1(_01762_),
    .Y(_01775_));
 sky130_fd_sc_hd__o21a_1 _07875_ (.A1(_01628_),
    .A2(_01632_),
    .B1(_01775_),
    .X(_01776_));
 sky130_fd_sc_hd__xor2_1 _07876_ (.A(_01774_),
    .B(_01775_),
    .X(_01777_));
 sky130_fd_sc_hd__xnor2_1 _07877_ (.A(_01629_),
    .B(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__o21ai_2 _07878_ (.A1(_01773_),
    .A2(_01778_),
    .B1(_01771_),
    .Y(_01779_));
 sky130_fd_sc_hd__xnor2_1 _07879_ (.A(_01654_),
    .B(_01656_),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2b_1 _07880_ (.A_N(_01781_),
    .B(_01779_),
    .Y(_01782_));
 sky130_fd_sc_hd__xnor2_1 _07881_ (.A(_01779_),
    .B(_01781_),
    .Y(_01783_));
 sky130_fd_sc_hd__a21oi_1 _07882_ (.A1(_01629_),
    .A2(_01777_),
    .B1(_01776_),
    .Y(_01784_));
 sky130_fd_sc_hd__nand2b_1 _07883_ (.A_N(_01784_),
    .B(_01783_),
    .Y(_01785_));
 sky130_fd_sc_hd__a211o_1 _07884_ (.A1(_01651_),
    .A2(_01646_),
    .B1(_01650_),
    .C1(_01662_),
    .X(_01786_));
 sky130_fd_sc_hd__nand2_1 _07885_ (.A(_01663_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__a21oi_1 _07886_ (.A1(_01782_),
    .A2(_01785_),
    .B1(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__and3_1 _07887_ (.A(_01782_),
    .B(_01785_),
    .C(_01787_),
    .X(_01789_));
 sky130_fd_sc_hd__nand2_1 _07888_ (.A(net8),
    .B(net33),
    .Y(_01790_));
 sky130_fd_sc_hd__nand2_1 _07889_ (.A(net8),
    .B(net44),
    .Y(_01792_));
 sky130_fd_sc_hd__nand4_2 _07890_ (.A(net9),
    .B(net8),
    .C(net44),
    .D(net33),
    .Y(_01793_));
 sky130_fd_sc_hd__a22o_1 _07891_ (.A1(net8),
    .A2(net44),
    .B1(net33),
    .B2(net9),
    .X(_01794_));
 sky130_fd_sc_hd__nand4_2 _07892_ (.A(_01794_),
    .B(net55),
    .C(net7),
    .D(_01793_),
    .Y(_01795_));
 sky130_fd_sc_hd__nand2_1 _07893_ (.A(_01793_),
    .B(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__a22o_1 _07894_ (.A1(net8),
    .A2(net55),
    .B1(_01668_),
    .B2(_01669_),
    .X(_01797_));
 sky130_fd_sc_hd__nand3_2 _07895_ (.A(_01671_),
    .B(_01796_),
    .C(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__a22o_1 _07896_ (.A1(net6),
    .A2(net59),
    .B1(net58),
    .B2(net7),
    .X(_01799_));
 sky130_fd_sc_hd__nand4_2 _07897_ (.A(net7),
    .B(net6),
    .C(net59),
    .D(net58),
    .Y(_01800_));
 sky130_fd_sc_hd__nand4_2 _07898_ (.A(_01799_),
    .B(_01800_),
    .C(net5),
    .D(net60),
    .Y(_01801_));
 sky130_fd_sc_hd__a22o_1 _07899_ (.A1(net5),
    .A2(net60),
    .B1(_01799_),
    .B2(_01800_),
    .X(_01803_));
 sky130_fd_sc_hd__a21o_1 _07900_ (.A1(_01671_),
    .A2(_01797_),
    .B1(_01796_),
    .X(_01804_));
 sky130_fd_sc_hd__nand4_2 _07901_ (.A(_01798_),
    .B(_01801_),
    .C(_01803_),
    .D(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__a21o_1 _07902_ (.A1(_01675_),
    .A2(_01682_),
    .B1(_01680_),
    .X(_01806_));
 sky130_fd_sc_hd__nand3_1 _07903_ (.A(_01675_),
    .B(_01680_),
    .C(_01682_),
    .Y(_01807_));
 sky130_fd_sc_hd__a22o_1 _07904_ (.A1(_01798_),
    .A2(_01805_),
    .B1(_01806_),
    .B2(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__nand4_1 _07905_ (.A(net4),
    .B(net3),
    .C(net62),
    .D(net61),
    .Y(_01809_));
 sky130_fd_sc_hd__a22o_1 _07906_ (.A1(net3),
    .A2(net62),
    .B1(net61),
    .B2(net4),
    .X(_01810_));
 sky130_fd_sc_hd__nand4_1 _07907_ (.A(_01810_),
    .B(net63),
    .C(net2),
    .D(_01809_),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_1 _07908_ (.A(_01809_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _07909_ (.A(_01800_),
    .B(_01801_),
    .Y(_01814_));
 sky130_fd_sc_hd__a22o_1 _07910_ (.A1(net3),
    .A2(net63),
    .B1(_01686_),
    .B2(_01687_),
    .X(_01815_));
 sky130_fd_sc_hd__a21o_1 _07911_ (.A1(_01688_),
    .A2(_01815_),
    .B1(_01814_),
    .X(_01816_));
 sky130_fd_sc_hd__nand3_1 _07912_ (.A(_01688_),
    .B(_01814_),
    .C(_01815_),
    .Y(_01817_));
 sky130_fd_sc_hd__and3_1 _07913_ (.A(_01812_),
    .B(_01816_),
    .C(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__a21oi_1 _07914_ (.A1(_01816_),
    .A2(_01817_),
    .B1(_01812_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand4_1 _07915_ (.A(_01798_),
    .B(_01805_),
    .C(_01806_),
    .D(_01807_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2_1 _07916_ (.A(_01808_),
    .B(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__or3_1 _07917_ (.A(_01818_),
    .B(_01819_),
    .C(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__a21o_1 _07918_ (.A1(_01685_),
    .A2(_01700_),
    .B1(_01699_),
    .X(_01823_));
 sky130_fd_sc_hd__nand3_1 _07919_ (.A(_01685_),
    .B(_01699_),
    .C(_01700_),
    .Y(_01825_));
 sky130_fd_sc_hd__a22o_1 _07920_ (.A1(_01808_),
    .A2(_01822_),
    .B1(_01823_),
    .B2(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _07921_ (.A(net64),
    .B(net31),
    .Y(_01827_));
 sky130_fd_sc_hd__or2_1 _07922_ (.A(_01706_),
    .B(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__a22o_1 _07923_ (.A1(net64),
    .A2(net32),
    .B1(net31),
    .B2(net34),
    .X(_01829_));
 sky130_fd_sc_hd__o2111ai_4 _07924_ (.A1(_01706_),
    .A2(_01827_),
    .B1(net35),
    .C1(net30),
    .D1(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__o21ai_1 _07925_ (.A1(_01706_),
    .A2(_01827_),
    .B1(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__a22o_1 _07926_ (.A1(net35),
    .A2(net31),
    .B1(_01707_),
    .B2(_01708_),
    .X(_01832_));
 sky130_fd_sc_hd__and3_1 _07927_ (.A(_01709_),
    .B(_01831_),
    .C(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__nand3_1 _07928_ (.A(_01709_),
    .B(_01831_),
    .C(_01832_),
    .Y(_01834_));
 sky130_fd_sc_hd__a22oi_1 _07929_ (.A1(net38),
    .A2(net28),
    .B1(_01729_),
    .B2(_01730_),
    .Y(_01836_));
 sky130_fd_sc_hd__a21o_1 _07930_ (.A1(_01709_),
    .A2(_01832_),
    .B1(_01831_),
    .X(_01837_));
 sky130_fd_sc_hd__or4b_2 _07931_ (.A(_01731_),
    .B(_01833_),
    .C(_01836_),
    .D_N(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__nand2_1 _07932_ (.A(_01834_),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__a31o_1 _07933_ (.A1(_01688_),
    .A2(_01814_),
    .A3(_01815_),
    .B1(_01818_),
    .X(_01840_));
 sky130_fd_sc_hd__a22o_1 _07934_ (.A1(_01607_),
    .A2(_01712_),
    .B1(_01713_),
    .B2(_01711_),
    .X(_01841_));
 sky130_fd_sc_hd__a21oi_1 _07935_ (.A1(_01715_),
    .A2(_01841_),
    .B1(_01840_),
    .Y(_01842_));
 sky130_fd_sc_hd__and3_1 _07936_ (.A(_01715_),
    .B(_01840_),
    .C(_01841_),
    .X(_01843_));
 sky130_fd_sc_hd__nor2_1 _07937_ (.A(_01842_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__a211oi_1 _07938_ (.A1(_01834_),
    .A2(_01838_),
    .B1(_01842_),
    .C1(_01843_),
    .Y(_01845_));
 sky130_fd_sc_hd__o211a_1 _07939_ (.A1(_01842_),
    .A2(_01843_),
    .B1(_01834_),
    .C1(_01838_),
    .X(_01847_));
 sky130_fd_sc_hd__nor2_1 _07940_ (.A(_01845_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand4_1 _07941_ (.A(_01808_),
    .B(_01822_),
    .C(_01823_),
    .D(_01825_),
    .Y(_01849_));
 sky130_fd_sc_hd__nand3_1 _07942_ (.A(_01848_),
    .B(_01849_),
    .C(_01826_),
    .Y(_01850_));
 sky130_fd_sc_hd__nand2_1 _07943_ (.A(_01826_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__a21o_1 _07944_ (.A1(_01705_),
    .A2(_01722_),
    .B1(_01721_),
    .X(_01852_));
 sky130_fd_sc_hd__nand3_1 _07945_ (.A(_01723_),
    .B(_01851_),
    .C(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__and4_1 _07946_ (.A(net37),
    .B(net36),
    .C(net29),
    .D(net28),
    .X(_01854_));
 sky130_fd_sc_hd__nand4_1 _07947_ (.A(net37),
    .B(net36),
    .C(net29),
    .D(net28),
    .Y(_01855_));
 sky130_fd_sc_hd__a22o_1 _07948_ (.A1(net36),
    .A2(net29),
    .B1(net28),
    .B2(net37),
    .X(_01856_));
 sky130_fd_sc_hd__and4_1 _07949_ (.A(_01856_),
    .B(net27),
    .C(net38),
    .D(_01855_),
    .X(_01858_));
 sky130_fd_sc_hd__a22o_1 _07950_ (.A1(net41),
    .A2(net23),
    .B1(_01734_),
    .B2(_01735_),
    .X(_01859_));
 sky130_fd_sc_hd__o211ai_2 _07951_ (.A1(_01854_),
    .A2(_01858_),
    .B1(_01859_),
    .C1(_01737_),
    .Y(_01860_));
 sky130_fd_sc_hd__and4_1 _07952_ (.A(net40),
    .B(net39),
    .C(net26),
    .D(net23),
    .X(_01861_));
 sky130_fd_sc_hd__nand4_2 _07953_ (.A(net40),
    .B(net39),
    .C(net26),
    .D(net23),
    .Y(_01862_));
 sky130_fd_sc_hd__a22o_1 _07954_ (.A1(net39),
    .A2(net26),
    .B1(net23),
    .B2(net40),
    .X(_01863_));
 sky130_fd_sc_hd__nand4_2 _07955_ (.A(_01863_),
    .B(net12),
    .C(net41),
    .D(_01862_),
    .Y(_01864_));
 sky130_fd_sc_hd__a31oi_1 _07956_ (.A1(_01863_),
    .A2(net12),
    .A3(net41),
    .B1(_01861_),
    .Y(_01865_));
 sky130_fd_sc_hd__a31o_1 _07957_ (.A1(_01863_),
    .A2(net12),
    .A3(net41),
    .B1(_01861_),
    .X(_01866_));
 sky130_fd_sc_hd__a211o_1 _07958_ (.A1(_01737_),
    .A2(_01859_),
    .B1(_01858_),
    .C1(_01854_),
    .X(_01867_));
 sky130_fd_sc_hd__a21bo_1 _07959_ (.A1(_01866_),
    .A2(_01867_),
    .B1_N(_01860_),
    .X(_01869_));
 sky130_fd_sc_hd__a22o_1 _07960_ (.A1(_01734_),
    .A2(_01737_),
    .B1(_01739_),
    .B2(_01733_),
    .X(_01870_));
 sky130_fd_sc_hd__nand3b_1 _07961_ (.A_N(_01738_),
    .B(_01739_),
    .C(_01733_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21bo_1 _07962_ (.A1(_01870_),
    .A2(_01871_),
    .B1_N(_01869_),
    .X(_01872_));
 sky130_fd_sc_hd__nand2_1 _07963_ (.A(net42),
    .B(net1),
    .Y(_01873_));
 sky130_fd_sc_hd__and4_1 _07964_ (.A(net43),
    .B(net42),
    .C(net12),
    .D(net1),
    .X(_01874_));
 sky130_fd_sc_hd__o2bb2a_1 _07965_ (.A1_N(_01743_),
    .A2_N(_01744_),
    .B1(_01054_),
    .B2(_01263_),
    .X(_01875_));
 sky130_fd_sc_hd__nor2_1 _07966_ (.A(_01745_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__a41o_1 _07967_ (.A1(net43),
    .A2(net42),
    .A3(net12),
    .A4(net1),
    .B1(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__or4b_1 _07968_ (.A(_01065_),
    .B(_01241_),
    .C(_01873_),
    .D_N(_01876_),
    .X(_01878_));
 sky130_fd_sc_hd__and2_1 _07969_ (.A(_01877_),
    .B(_01878_),
    .X(_01880_));
 sky130_fd_sc_hd__nand3b_1 _07970_ (.A_N(_01869_),
    .B(_01870_),
    .C(_01871_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_1 _07971_ (.A(_01872_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__nand3_1 _07972_ (.A(_01872_),
    .B(_01880_),
    .C(_01881_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand2_1 _07973_ (.A(_01754_),
    .B(_01756_),
    .Y(_01884_));
 sky130_fd_sc_hd__a221o_1 _07974_ (.A1(_01844_),
    .A2(_01839_),
    .B1(_01757_),
    .B2(_01884_),
    .C1(_01843_),
    .X(_01885_));
 sky130_fd_sc_hd__o211ai_2 _07975_ (.A1(_01843_),
    .A2(_01845_),
    .B1(_01884_),
    .C1(_01757_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__a21o_1 _07977_ (.A1(_01872_),
    .A2(_01883_),
    .B1(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__nand3_1 _07978_ (.A(_01872_),
    .B(_01883_),
    .C(_01887_),
    .Y(_01889_));
 sky130_fd_sc_hd__and2_1 _07979_ (.A(_01888_),
    .B(_01889_),
    .X(_01891_));
 sky130_fd_sc_hd__a21o_1 _07980_ (.A1(_01723_),
    .A2(_01852_),
    .B1(_01851_),
    .X(_01892_));
 sky130_fd_sc_hd__and2_1 _07981_ (.A(_01853_),
    .B(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__nand2_1 _07982_ (.A(_01891_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__or2_1 _07983_ (.A(_01764_),
    .B(_01766_),
    .X(_01895_));
 sky130_fd_sc_hd__nand2_1 _07984_ (.A(_01767_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__a21o_1 _07985_ (.A1(_01853_),
    .A2(_01894_),
    .B1(_01896_),
    .X(_01897_));
 sky130_fd_sc_hd__a31oi_1 _07986_ (.A1(net46),
    .A2(net1),
    .A3(_01751_),
    .B1(_01750_),
    .Y(_01898_));
 sky130_fd_sc_hd__and3_1 _07987_ (.A(_01886_),
    .B(_01888_),
    .C(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__a21oi_1 _07988_ (.A1(_01886_),
    .A2(_01888_),
    .B1(_01898_),
    .Y(_01900_));
 sky130_fd_sc_hd__or2_1 _07989_ (.A(_01899_),
    .B(_01900_),
    .X(_01902_));
 sky130_fd_sc_hd__nand3_1 _07990_ (.A(_01853_),
    .B(_01894_),
    .C(_01896_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _07991_ (.A(_01897_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__or2_1 _07992_ (.A(_01902_),
    .B(_01904_),
    .X(_01905_));
 sky130_fd_sc_hd__xnor2_1 _07993_ (.A(_01773_),
    .B(_01778_),
    .Y(_01906_));
 sky130_fd_sc_hd__a21o_1 _07994_ (.A1(_01897_),
    .A2(_01905_),
    .B1(_01906_),
    .X(_01907_));
 sky130_fd_sc_hd__o211ai_1 _07995_ (.A1(_01902_),
    .A2(_01904_),
    .B1(_01906_),
    .C1(_01897_),
    .Y(_01908_));
 sky130_fd_sc_hd__and2_1 _07996_ (.A(_01907_),
    .B(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__a21bo_1 _07997_ (.A1(_01900_),
    .A2(_01909_),
    .B1_N(_01907_),
    .X(_01910_));
 sky130_fd_sc_hd__xnor2_1 _07998_ (.A(_01783_),
    .B(_01784_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_1 _07999_ (.A(_01911_),
    .B(_01910_),
    .Y(_01913_));
 sky130_fd_sc_hd__xor2_1 _08000_ (.A(_01910_),
    .B(_01911_),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_1 _08001_ (.A(net7),
    .B(net33),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _08002_ (.A(net7),
    .B(net44),
    .Y(_01916_));
 sky130_fd_sc_hd__and2_1 _08003_ (.A(net6),
    .B(net55),
    .X(_01917_));
 sky130_fd_sc_hd__a22o_1 _08004_ (.A1(net7),
    .A2(net44),
    .B1(net33),
    .B2(net8),
    .X(_01918_));
 sky130_fd_sc_hd__nand3_1 _08005_ (.A(_01916_),
    .B(net33),
    .C(net8),
    .Y(_01919_));
 sky130_fd_sc_hd__nand3_1 _08006_ (.A(_01790_),
    .B(net44),
    .C(net7),
    .Y(_01920_));
 sky130_fd_sc_hd__o2111ai_2 _08007_ (.A1(_01792_),
    .A2(_01915_),
    .B1(net6),
    .C1(net55),
    .D1(_01918_),
    .Y(_01921_));
 sky130_fd_sc_hd__a2bb2o_1 _08008_ (.A1_N(_01792_),
    .A2_N(_01915_),
    .B1(_01917_),
    .B2(_01918_),
    .X(_01922_));
 sky130_fd_sc_hd__a22o_1 _08009_ (.A1(net7),
    .A2(net55),
    .B1(_01793_),
    .B2(_01794_),
    .X(_01924_));
 sky130_fd_sc_hd__nand3_2 _08010_ (.A(_01795_),
    .B(_01922_),
    .C(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand4_2 _08011_ (.A(net6),
    .B(net5),
    .C(net59),
    .D(net58),
    .Y(_01926_));
 sky130_fd_sc_hd__a22o_1 _08012_ (.A1(net5),
    .A2(net59),
    .B1(net58),
    .B2(net6),
    .X(_01927_));
 sky130_fd_sc_hd__nand4_2 _08013_ (.A(_01927_),
    .B(net60),
    .C(net4),
    .D(_01926_),
    .Y(_01928_));
 sky130_fd_sc_hd__a22o_1 _08014_ (.A1(net4),
    .A2(net60),
    .B1(_01926_),
    .B2(_01927_),
    .X(_01929_));
 sky130_fd_sc_hd__nand2_1 _08015_ (.A(_01928_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__a21o_1 _08016_ (.A1(_01795_),
    .A2(_01924_),
    .B1(_01922_),
    .X(_01931_));
 sky130_fd_sc_hd__nand4_1 _08017_ (.A(_01925_),
    .B(_01928_),
    .C(_01929_),
    .D(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_1 _08018_ (.A(_01925_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__a22o_1 _08019_ (.A1(_01801_),
    .A2(_01803_),
    .B1(_01804_),
    .B2(_01798_),
    .X(_01935_));
 sky130_fd_sc_hd__nand3_1 _08020_ (.A(_01805_),
    .B(_01933_),
    .C(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand4_2 _08021_ (.A(net3),
    .B(net2),
    .C(net62),
    .D(net61),
    .Y(_01937_));
 sky130_fd_sc_hd__a22o_1 _08022_ (.A1(net2),
    .A2(net62),
    .B1(net61),
    .B2(net3),
    .X(_01938_));
 sky130_fd_sc_hd__nand4_2 _08023_ (.A(_01938_),
    .B(net63),
    .C(net32),
    .D(_01937_),
    .Y(_01939_));
 sky130_fd_sc_hd__nand2_1 _08024_ (.A(_01937_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__nand2_1 _08025_ (.A(_01926_),
    .B(_01928_),
    .Y(_01941_));
 sky130_fd_sc_hd__a22o_1 _08026_ (.A1(net2),
    .A2(net63),
    .B1(_01809_),
    .B2(_01810_),
    .X(_01942_));
 sky130_fd_sc_hd__nand3_1 _08027_ (.A(_01811_),
    .B(_01941_),
    .C(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21o_1 _08028_ (.A1(_01811_),
    .A2(_01942_),
    .B1(_01941_),
    .X(_01944_));
 sky130_fd_sc_hd__nand3_1 _08029_ (.A(_01940_),
    .B(_01943_),
    .C(_01944_),
    .Y(_01946_));
 sky130_fd_sc_hd__a21o_1 _08030_ (.A1(_01943_),
    .A2(_01944_),
    .B1(_01940_),
    .X(_01947_));
 sky130_fd_sc_hd__and2_1 _08031_ (.A(_01946_),
    .B(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__a21o_1 _08032_ (.A1(_01805_),
    .A2(_01935_),
    .B1(_01933_),
    .X(_01949_));
 sky130_fd_sc_hd__nand2_1 _08033_ (.A(_01936_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__a21bo_1 _08034_ (.A1(_01949_),
    .A2(_01948_),
    .B1_N(_01936_),
    .X(_01951_));
 sky130_fd_sc_hd__a2bb2o_1 _08035_ (.A1_N(_01818_),
    .A2_N(_01819_),
    .B1(_01820_),
    .B2(_01808_),
    .X(_01952_));
 sky130_fd_sc_hd__nand3_1 _08036_ (.A(_01822_),
    .B(_01951_),
    .C(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__nand4_2 _08037_ (.A(net34),
    .B(net64),
    .C(net31),
    .D(net30),
    .Y(_01954_));
 sky130_fd_sc_hd__a22o_1 _08038_ (.A1(net64),
    .A2(net31),
    .B1(net30),
    .B2(net34),
    .X(_01955_));
 sky130_fd_sc_hd__nand4_2 _08039_ (.A(_01955_),
    .B(net29),
    .C(net35),
    .D(_01954_),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _08040_ (.A(_01954_),
    .B(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__a22o_1 _08041_ (.A1(net35),
    .A2(net30),
    .B1(_01828_),
    .B2(_01829_),
    .X(_01959_));
 sky130_fd_sc_hd__and3_1 _08042_ (.A(_01830_),
    .B(_01958_),
    .C(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__nand3_1 _08043_ (.A(_01830_),
    .B(_01958_),
    .C(_01959_),
    .Y(_01961_));
 sky130_fd_sc_hd__o2bb2a_1 _08044_ (.A1_N(_01855_),
    .A2_N(_01856_),
    .B1(_01087_),
    .B2(_01208_),
    .X(_01962_));
 sky130_fd_sc_hd__or2_1 _08045_ (.A(_01858_),
    .B(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__a21o_1 _08046_ (.A1(_01830_),
    .A2(_01959_),
    .B1(_01958_),
    .X(_01964_));
 sky130_fd_sc_hd__and3b_1 _08047_ (.A_N(_01963_),
    .B(_01964_),
    .C(_01961_),
    .X(_01965_));
 sky130_fd_sc_hd__or4b_1 _08048_ (.A(_01858_),
    .B(_01960_),
    .C(_01962_),
    .D_N(_01964_),
    .X(_01966_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(_01943_),
    .B(_01946_),
    .Y(_01968_));
 sky130_fd_sc_hd__a2bb2o_1 _08050_ (.A1_N(_01731_),
    .A2_N(_01836_),
    .B1(_01837_),
    .B2(_01834_),
    .X(_01969_));
 sky130_fd_sc_hd__nand3_1 _08051_ (.A(_01838_),
    .B(_01968_),
    .C(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__a21o_1 _08052_ (.A1(_01838_),
    .A2(_01969_),
    .B1(_01968_),
    .X(_01971_));
 sky130_fd_sc_hd__o211ai_2 _08053_ (.A1(_01960_),
    .A2(_01965_),
    .B1(_01970_),
    .C1(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__a211o_1 _08054_ (.A1(_01970_),
    .A2(_01971_),
    .B1(_01960_),
    .C1(_01965_),
    .X(_01973_));
 sky130_fd_sc_hd__a21o_1 _08055_ (.A1(_01822_),
    .A2(_01952_),
    .B1(_01951_),
    .X(_01974_));
 sky130_fd_sc_hd__nand4_2 _08056_ (.A(_01953_),
    .B(_01972_),
    .C(_01973_),
    .D(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _08057_ (.A(_01953_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__a21o_1 _08058_ (.A1(_01826_),
    .A2(_01849_),
    .B1(_01848_),
    .X(_01977_));
 sky130_fd_sc_hd__nand3_1 _08059_ (.A(_01850_),
    .B(_01976_),
    .C(_01977_),
    .Y(_01979_));
 sky130_fd_sc_hd__and4_1 _08060_ (.A(net37),
    .B(net36),
    .C(net28),
    .D(net27),
    .X(_01980_));
 sky130_fd_sc_hd__nand4_1 _08061_ (.A(net37),
    .B(net36),
    .C(net28),
    .D(net27),
    .Y(_01981_));
 sky130_fd_sc_hd__a22o_1 _08062_ (.A1(net36),
    .A2(net28),
    .B1(net27),
    .B2(net37),
    .X(_01982_));
 sky130_fd_sc_hd__and4_1 _08063_ (.A(_01982_),
    .B(net26),
    .C(net38),
    .D(_01981_),
    .X(_01983_));
 sky130_fd_sc_hd__a22o_1 _08064_ (.A1(net41),
    .A2(net12),
    .B1(_01862_),
    .B2(_01863_),
    .X(_01984_));
 sky130_fd_sc_hd__o211ai_2 _08065_ (.A1(_01980_),
    .A2(_01983_),
    .B1(_01984_),
    .C1(_01864_),
    .Y(_01985_));
 sky130_fd_sc_hd__and4_1 _08066_ (.A(net40),
    .B(net39),
    .C(net23),
    .D(net12),
    .X(_01986_));
 sky130_fd_sc_hd__a22oi_1 _08067_ (.A1(net39),
    .A2(net23),
    .B1(net12),
    .B2(net40),
    .Y(_01987_));
 sky130_fd_sc_hd__a22o_1 _08068_ (.A1(net39),
    .A2(net23),
    .B1(net12),
    .B2(net40),
    .X(_01988_));
 sky130_fd_sc_hd__and4b_1 _08069_ (.A_N(_01986_),
    .B(_01988_),
    .C(net41),
    .D(net1),
    .X(_01990_));
 sky130_fd_sc_hd__a31o_1 _08070_ (.A1(_01988_),
    .A2(net1),
    .A3(net41),
    .B1(_01986_),
    .X(_01991_));
 sky130_fd_sc_hd__a211o_1 _08071_ (.A1(_01864_),
    .A2(_01984_),
    .B1(_01983_),
    .C1(_01980_),
    .X(_01992_));
 sky130_fd_sc_hd__o211ai_2 _08072_ (.A1(_01986_),
    .A2(_01990_),
    .B1(_01992_),
    .C1(_01985_),
    .Y(_01993_));
 sky130_fd_sc_hd__a22o_1 _08073_ (.A1(_01862_),
    .A2(_01864_),
    .B1(_01867_),
    .B2(_01860_),
    .X(_01994_));
 sky130_fd_sc_hd__nand3_1 _08074_ (.A(_01860_),
    .B(_01867_),
    .C(_01865_),
    .Y(_01995_));
 sky130_fd_sc_hd__a22o_1 _08075_ (.A1(_01985_),
    .A2(_01993_),
    .B1(_01994_),
    .B2(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__o2bb2a_1 _08076_ (.A1_N(net42),
    .A2_N(net12),
    .B1(_01263_),
    .B2(_01065_),
    .X(_01997_));
 sky130_fd_sc_hd__nand4_1 _08077_ (.A(_01985_),
    .B(_01993_),
    .C(_01994_),
    .D(_01995_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(_01996_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor3_1 _08079_ (.A(_01874_),
    .B(_01997_),
    .C(_01999_),
    .Y(_02001_));
 sky130_fd_sc_hd__o31a_1 _08080_ (.A1(_01874_),
    .A2(_01997_),
    .A3(_01999_),
    .B1(_01996_),
    .X(_02002_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_01882_),
    .B(_01880_),
    .Y(_02003_));
 sky130_fd_sc_hd__or2_1 _08082_ (.A(_01880_),
    .B(_01882_),
    .X(_02004_));
 sky130_fd_sc_hd__a22oi_1 _08083_ (.A1(_01970_),
    .A2(_01972_),
    .B1(_02003_),
    .B2(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__and4_1 _08084_ (.A(_01970_),
    .B(_01972_),
    .C(_02003_),
    .D(_02004_),
    .X(_02006_));
 sky130_fd_sc_hd__nor2_1 _08085_ (.A(_02005_),
    .B(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__xnor2_1 _08086_ (.A(_02002_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__a21o_1 _08087_ (.A1(_01850_),
    .A2(_01977_),
    .B1(_01976_),
    .X(_02009_));
 sky130_fd_sc_hd__nand3_1 _08088_ (.A(_02008_),
    .B(_02009_),
    .C(_01979_),
    .Y(_02010_));
 sky130_fd_sc_hd__xnor2_1 _08089_ (.A(_01891_),
    .B(_01893_),
    .Y(_02012_));
 sky130_fd_sc_hd__a21o_1 _08090_ (.A1(_01979_),
    .A2(_02010_),
    .B1(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__o21bai_1 _08091_ (.A1(_02002_),
    .A2(_02006_),
    .B1_N(_02005_),
    .Y(_02014_));
 sky130_fd_sc_hd__and3_1 _08092_ (.A(_02014_),
    .B(_01876_),
    .C(_01874_),
    .X(_02015_));
 sky130_fd_sc_hd__xor2_1 _08093_ (.A(_01878_),
    .B(_02014_),
    .X(_02016_));
 sky130_fd_sc_hd__nand3_1 _08094_ (.A(_01979_),
    .B(_02010_),
    .C(_02012_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand2_1 _08095_ (.A(_02013_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__or2_1 _08096_ (.A(_02016_),
    .B(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__nand2_1 _08097_ (.A(_01902_),
    .B(_01904_),
    .Y(_02020_));
 sky130_fd_sc_hd__nand2_1 _08098_ (.A(_01905_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__a21oi_1 _08099_ (.A1(_02013_),
    .A2(_02019_),
    .B1(_02021_),
    .Y(_02023_));
 sky130_fd_sc_hd__and3_1 _08100_ (.A(_02013_),
    .B(_02019_),
    .C(_02021_),
    .X(_02024_));
 sky130_fd_sc_hd__nor2_1 _08101_ (.A(_02023_),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__a21oi_2 _08102_ (.A1(_02015_),
    .A2(_02025_),
    .B1(_02023_),
    .Y(_02026_));
 sky130_fd_sc_hd__xnor2_1 _08103_ (.A(_01900_),
    .B(_01909_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _08104_ (.A(_02026_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__and2_1 _08105_ (.A(_02027_),
    .B(_02026_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _08106_ (.A(net2),
    .B(net44),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _08107_ (.A(net32),
    .B(net33),
    .Y(_02031_));
 sky130_fd_sc_hd__nand2_1 _08108_ (.A(net2),
    .B(net33),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_1 _08109_ (.A(net32),
    .B(net44),
    .Y(_02034_));
 sky130_fd_sc_hd__a22o_1 _08110_ (.A1(net32),
    .A2(net44),
    .B1(net33),
    .B2(net2),
    .X(_02035_));
 sky130_fd_sc_hd__nand3_1 _08111_ (.A(_02034_),
    .B(net33),
    .C(net2),
    .Y(_02036_));
 sky130_fd_sc_hd__nand3_1 _08112_ (.A(_02032_),
    .B(net44),
    .C(net32),
    .Y(_02037_));
 sky130_fd_sc_hd__o2111ai_4 _08113_ (.A1(_02030_),
    .A2(_02031_),
    .B1(net31),
    .C1(net55),
    .D1(_02035_),
    .Y(_02038_));
 sky130_fd_sc_hd__o21ai_1 _08114_ (.A1(_02032_),
    .A2(_02034_),
    .B1(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2_1 _08115_ (.A(net3),
    .B(net44),
    .Y(_02040_));
 sky130_fd_sc_hd__and4_1 _08116_ (.A(net3),
    .B(net2),
    .C(net44),
    .D(net33),
    .X(_02041_));
 sky130_fd_sc_hd__nand4_1 _08117_ (.A(net3),
    .B(net2),
    .C(net44),
    .D(net33),
    .Y(_02042_));
 sky130_fd_sc_hd__a22oi_2 _08118_ (.A1(net2),
    .A2(net44),
    .B1(net33),
    .B2(net3),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _08119_ (.A(net32),
    .B(net55),
    .Y(_02045_));
 sky130_fd_sc_hd__nand4b_1 _08120_ (.A_N(_02043_),
    .B(net55),
    .C(net32),
    .D(_02042_),
    .Y(_02046_));
 sky130_fd_sc_hd__o21ai_1 _08121_ (.A1(_02041_),
    .A2(_02043_),
    .B1(_02045_),
    .Y(_02047_));
 sky130_fd_sc_hd__nand3_1 _08122_ (.A(_02039_),
    .B(_02046_),
    .C(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__a22o_1 _08123_ (.A1(net30),
    .A2(net59),
    .B1(net58),
    .B2(net31),
    .X(_02049_));
 sky130_fd_sc_hd__and4_1 _08124_ (.A(net31),
    .B(net30),
    .C(net59),
    .D(net58),
    .X(_02050_));
 sky130_fd_sc_hd__nand4_1 _08125_ (.A(net31),
    .B(net30),
    .C(net59),
    .D(net58),
    .Y(_02051_));
 sky130_fd_sc_hd__or4b_1 _08126_ (.A(_01186_),
    .B(_02050_),
    .C(_01197_),
    .D_N(_02049_),
    .X(_02052_));
 sky130_fd_sc_hd__a22o_1 _08127_ (.A1(net29),
    .A2(net60),
    .B1(_02049_),
    .B2(_02051_),
    .X(_02053_));
 sky130_fd_sc_hd__a21o_1 _08128_ (.A1(_02046_),
    .A2(_02047_),
    .B1(_02039_),
    .X(_02054_));
 sky130_fd_sc_hd__nand4_2 _08129_ (.A(_02048_),
    .B(_02052_),
    .C(_02053_),
    .D(_02054_),
    .Y(_02056_));
 sky130_fd_sc_hd__nand2_1 _08130_ (.A(_02048_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__a22o_1 _08131_ (.A1(net31),
    .A2(net59),
    .B1(net58),
    .B2(net32),
    .X(_02058_));
 sky130_fd_sc_hd__nand4_1 _08132_ (.A(net32),
    .B(net31),
    .C(net59),
    .D(net58),
    .Y(_02059_));
 sky130_fd_sc_hd__and4_1 _08133_ (.A(_02058_),
    .B(_02059_),
    .C(net30),
    .D(net60),
    .X(_02060_));
 sky130_fd_sc_hd__o2bb2a_1 _08134_ (.A1_N(_02058_),
    .A2_N(_02059_),
    .B1(_01175_),
    .B2(_01197_),
    .X(_02061_));
 sky130_fd_sc_hd__o21ai_1 _08135_ (.A1(_02045_),
    .A2(_02043_),
    .B1(_02042_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _08136_ (.A(net4),
    .B(net33),
    .Y(_02063_));
 sky130_fd_sc_hd__nand4_1 _08137_ (.A(net4),
    .B(net3),
    .C(net44),
    .D(net33),
    .Y(_02064_));
 sky130_fd_sc_hd__a22o_1 _08138_ (.A1(net3),
    .A2(net44),
    .B1(net33),
    .B2(net4),
    .X(_02065_));
 sky130_fd_sc_hd__nand4_2 _08139_ (.A(_02065_),
    .B(net55),
    .C(net2),
    .D(_02064_),
    .Y(_02067_));
 sky130_fd_sc_hd__o2bb2ai_1 _08140_ (.A1_N(_02064_),
    .A2_N(_02065_),
    .B1(_01131_),
    .B2(_01230_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand3_1 _08141_ (.A(_02062_),
    .B(_02067_),
    .C(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21oi_1 _08142_ (.A1(_02067_),
    .A2(_02068_),
    .B1(_02062_),
    .Y(_02070_));
 sky130_fd_sc_hd__a21o_1 _08143_ (.A1(_02067_),
    .A2(_02068_),
    .B1(_02062_),
    .X(_02071_));
 sky130_fd_sc_hd__or4bb_1 _08144_ (.A(_02060_),
    .B(_02061_),
    .C_N(_02069_),
    .D_N(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__a2bb2o_1 _08145_ (.A1_N(_02060_),
    .A2_N(_02061_),
    .B1(_02069_),
    .B2(_02071_),
    .X(_02073_));
 sky130_fd_sc_hd__nand3_1 _08146_ (.A(_02057_),
    .B(_02072_),
    .C(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2_1 _08147_ (.A(net61),
    .B(net28),
    .Y(_02075_));
 sky130_fd_sc_hd__nand4_2 _08148_ (.A(net62),
    .B(net61),
    .C(net28),
    .D(net27),
    .Y(_02076_));
 sky130_fd_sc_hd__a22o_1 _08149_ (.A1(net61),
    .A2(net28),
    .B1(net27),
    .B2(net62),
    .X(_02078_));
 sky130_fd_sc_hd__nand4_2 _08150_ (.A(_02078_),
    .B(net26),
    .C(net63),
    .D(_02076_),
    .Y(_02079_));
 sky130_fd_sc_hd__o31a_1 _08151_ (.A1(_01164_),
    .A2(_01208_),
    .A3(_02075_),
    .B1(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__nand2_1 _08152_ (.A(_02076_),
    .B(_02079_),
    .Y(_02081_));
 sky130_fd_sc_hd__a31o_1 _08153_ (.A1(_02049_),
    .A2(net60),
    .A3(net29),
    .B1(_02050_),
    .X(_02082_));
 sky130_fd_sc_hd__and4_1 _08154_ (.A(net62),
    .B(net61),
    .C(net29),
    .D(net28),
    .X(_02083_));
 sky130_fd_sc_hd__or3_1 _08155_ (.A(_01164_),
    .B(_01186_),
    .C(_02075_),
    .X(_02084_));
 sky130_fd_sc_hd__a22oi_1 _08156_ (.A1(net61),
    .A2(net29),
    .B1(net28),
    .B2(net62),
    .Y(_02085_));
 sky130_fd_sc_hd__or4bb_2 _08157_ (.A(_02083_),
    .B(_02085_),
    .C_N(net63),
    .D_N(net27),
    .X(_02086_));
 sky130_fd_sc_hd__a2bb2o_1 _08158_ (.A1_N(_02083_),
    .A2_N(_02085_),
    .B1(net63),
    .B2(net27),
    .X(_02087_));
 sky130_fd_sc_hd__a21oi_1 _08159_ (.A1(_02086_),
    .A2(_02087_),
    .B1(_02082_),
    .Y(_02089_));
 sky130_fd_sc_hd__a21o_1 _08160_ (.A1(_02086_),
    .A2(_02087_),
    .B1(_02082_),
    .X(_02090_));
 sky130_fd_sc_hd__nand3_1 _08161_ (.A(_02082_),
    .B(_02086_),
    .C(_02087_),
    .Y(_02091_));
 sky130_fd_sc_hd__or3b_1 _08162_ (.A(_02080_),
    .B(_02089_),
    .C_N(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__a21o_1 _08163_ (.A1(_02090_),
    .A2(_02091_),
    .B1(_02081_),
    .X(_02093_));
 sky130_fd_sc_hd__a21o_1 _08164_ (.A1(_02072_),
    .A2(_02073_),
    .B1(_02057_),
    .X(_02094_));
 sky130_fd_sc_hd__nand4_2 _08165_ (.A(_02074_),
    .B(_02092_),
    .C(_02093_),
    .D(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__nand2_1 _08166_ (.A(_02074_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__a41o_1 _08167_ (.A1(net32),
    .A2(net31),
    .A3(net59),
    .A4(net58),
    .B1(_02060_),
    .X(_02097_));
 sky130_fd_sc_hd__and4_1 _08168_ (.A(net62),
    .B(net30),
    .C(net61),
    .D(net29),
    .X(_02098_));
 sky130_fd_sc_hd__nand4_1 _08169_ (.A(net62),
    .B(net30),
    .C(net61),
    .D(net29),
    .Y(_02100_));
 sky130_fd_sc_hd__a22o_1 _08170_ (.A1(net30),
    .A2(net61),
    .B1(net29),
    .B2(net62),
    .X(_02101_));
 sky130_fd_sc_hd__and4_1 _08171_ (.A(_02101_),
    .B(net28),
    .C(net63),
    .D(_02100_),
    .X(_02102_));
 sky130_fd_sc_hd__nand4_1 _08172_ (.A(_02101_),
    .B(net28),
    .C(net63),
    .D(_02100_),
    .Y(_02103_));
 sky130_fd_sc_hd__a22o_1 _08173_ (.A1(net63),
    .A2(net28),
    .B1(_02100_),
    .B2(_02101_),
    .X(_02104_));
 sky130_fd_sc_hd__a21oi_1 _08174_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_02097_),
    .Y(_02105_));
 sky130_fd_sc_hd__and3_1 _08175_ (.A(_02097_),
    .B(_02103_),
    .C(_02104_),
    .X(_02106_));
 sky130_fd_sc_hd__a211oi_2 _08176_ (.A1(_02084_),
    .A2(_02086_),
    .B1(_02105_),
    .C1(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__o211a_1 _08177_ (.A1(_02105_),
    .A2(_02106_),
    .B1(_02084_),
    .C1(_02086_),
    .X(_02108_));
 sky130_fd_sc_hd__o31a_1 _08178_ (.A1(_02060_),
    .A2(_02061_),
    .A3(_02070_),
    .B1(_02069_),
    .X(_02109_));
 sky130_fd_sc_hd__a22o_1 _08179_ (.A1(net32),
    .A2(net59),
    .B1(net58),
    .B2(net2),
    .X(_02111_));
 sky130_fd_sc_hd__nand4_1 _08180_ (.A(net2),
    .B(net32),
    .C(net59),
    .D(net58),
    .Y(_02112_));
 sky130_fd_sc_hd__nand4_1 _08181_ (.A(_02111_),
    .B(_02112_),
    .C(net31),
    .D(net60),
    .Y(_02113_));
 sky130_fd_sc_hd__a22o_1 _08182_ (.A1(net31),
    .A2(net60),
    .B1(_02111_),
    .B2(_02112_),
    .X(_02114_));
 sky130_fd_sc_hd__nand2_1 _08183_ (.A(_02113_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__o21ai_1 _08184_ (.A1(_02040_),
    .A2(_02063_),
    .B1(_02067_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2_1 _08185_ (.A(net5),
    .B(net44),
    .Y(_02117_));
 sky130_fd_sc_hd__and4_1 _08186_ (.A(net5),
    .B(net4),
    .C(net44),
    .D(net33),
    .X(_02118_));
 sky130_fd_sc_hd__nand4_1 _08187_ (.A(net5),
    .B(net4),
    .C(net44),
    .D(net33),
    .Y(_02119_));
 sky130_fd_sc_hd__a22o_1 _08188_ (.A1(net4),
    .A2(net44),
    .B1(net33),
    .B2(net5),
    .X(_02120_));
 sky130_fd_sc_hd__o2111ai_2 _08189_ (.A1(_02063_),
    .A2(_02117_),
    .B1(net3),
    .C1(net55),
    .D1(_02120_),
    .Y(_02122_));
 sky130_fd_sc_hd__a22o_1 _08190_ (.A1(net3),
    .A2(net55),
    .B1(_02119_),
    .B2(_02120_),
    .X(_02123_));
 sky130_fd_sc_hd__nand3_1 _08191_ (.A(_02116_),
    .B(_02122_),
    .C(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__a21oi_1 _08192_ (.A1(_02122_),
    .A2(_02123_),
    .B1(_02116_),
    .Y(_02125_));
 sky130_fd_sc_hd__a21o_1 _08193_ (.A1(_02122_),
    .A2(_02123_),
    .B1(_02116_),
    .X(_02126_));
 sky130_fd_sc_hd__a21oi_1 _08194_ (.A1(_02124_),
    .A2(_02126_),
    .B1(_02115_),
    .Y(_02127_));
 sky130_fd_sc_hd__and3_1 _08195_ (.A(_02115_),
    .B(_02124_),
    .C(_02126_),
    .X(_02128_));
 sky130_fd_sc_hd__o21bai_1 _08196_ (.A1(_02127_),
    .A2(_02128_),
    .B1_N(_02109_),
    .Y(_02129_));
 sky130_fd_sc_hd__or3b_1 _08197_ (.A(_02127_),
    .B(_02128_),
    .C_N(_02109_),
    .X(_02130_));
 sky130_fd_sc_hd__or4bb_1 _08198_ (.A(_02107_),
    .B(_02108_),
    .C_N(_02129_),
    .D_N(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__a2bb2o_1 _08199_ (.A1_N(_02107_),
    .A2_N(_02108_),
    .B1(_02129_),
    .B2(_02130_),
    .X(_02133_));
 sky130_fd_sc_hd__nand3_2 _08200_ (.A(_02096_),
    .B(_02131_),
    .C(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__and4_1 _08201_ (.A(net34),
    .B(net64),
    .C(net23),
    .D(net12),
    .X(_02135_));
 sky130_fd_sc_hd__a22oi_2 _08202_ (.A1(net64),
    .A2(net23),
    .B1(net12),
    .B2(net34),
    .Y(_02136_));
 sky130_fd_sc_hd__nor4_2 _08203_ (.A(_01109_),
    .B(_02136_),
    .C(_01263_),
    .D(_02135_),
    .Y(_02137_));
 sky130_fd_sc_hd__a41o_1 _08204_ (.A1(net34),
    .A2(net64),
    .A3(net23),
    .A4(net12),
    .B1(_02137_),
    .X(_02138_));
 sky130_fd_sc_hd__nand4_2 _08205_ (.A(net34),
    .B(net64),
    .C(net26),
    .D(net23),
    .Y(_02139_));
 sky130_fd_sc_hd__a22o_1 _08206_ (.A1(net64),
    .A2(net26),
    .B1(net23),
    .B2(net34),
    .X(_02140_));
 sky130_fd_sc_hd__nand4_2 _08207_ (.A(_02140_),
    .B(net12),
    .C(net35),
    .D(_02139_),
    .Y(_02141_));
 sky130_fd_sc_hd__a22o_1 _08208_ (.A1(net35),
    .A2(net12),
    .B1(_02139_),
    .B2(_02140_),
    .X(_02142_));
 sky130_fd_sc_hd__o211ai_2 _08209_ (.A1(_02135_),
    .A2(_02137_),
    .B1(_02141_),
    .C1(_02142_),
    .Y(_02144_));
 sky130_fd_sc_hd__nand2_1 _08210_ (.A(net36),
    .B(net1),
    .Y(_02145_));
 sky130_fd_sc_hd__a21oi_1 _08211_ (.A1(_02141_),
    .A2(_02142_),
    .B1(_02138_),
    .Y(_02146_));
 sky130_fd_sc_hd__a211o_1 _08212_ (.A1(_02141_),
    .A2(_02142_),
    .B1(_02135_),
    .C1(_02137_),
    .X(_02147_));
 sky130_fd_sc_hd__o21a_1 _08213_ (.A1(_02145_),
    .A2(_02146_),
    .B1(_02144_),
    .X(_02148_));
 sky130_fd_sc_hd__o21ai_1 _08214_ (.A1(_02080_),
    .A2(_02089_),
    .B1(_02091_),
    .Y(_02149_));
 sky130_fd_sc_hd__and4_1 _08215_ (.A(net37),
    .B(net36),
    .C(net12),
    .D(net1),
    .X(_02150_));
 sky130_fd_sc_hd__a22oi_1 _08216_ (.A1(net36),
    .A2(net12),
    .B1(net1),
    .B2(net37),
    .Y(_02151_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_02139_),
    .B(_02141_),
    .Y(_02152_));
 sky130_fd_sc_hd__nand4_1 _08218_ (.A(net34),
    .B(net64),
    .C(net27),
    .D(net26),
    .Y(_02153_));
 sky130_fd_sc_hd__a22o_1 _08219_ (.A1(net64),
    .A2(net27),
    .B1(net26),
    .B2(net34),
    .X(_02155_));
 sky130_fd_sc_hd__nand4_1 _08220_ (.A(_02155_),
    .B(net23),
    .C(net35),
    .D(_02153_),
    .Y(_02156_));
 sky130_fd_sc_hd__a22o_1 _08221_ (.A1(net35),
    .A2(net23),
    .B1(_02153_),
    .B2(_02155_),
    .X(_02157_));
 sky130_fd_sc_hd__nand3_1 _08222_ (.A(_02152_),
    .B(_02156_),
    .C(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21o_1 _08223_ (.A1(_02156_),
    .A2(_02157_),
    .B1(_02152_),
    .X(_02159_));
 sky130_fd_sc_hd__or4bb_1 _08224_ (.A(_02150_),
    .B(_02151_),
    .C_N(_02158_),
    .D_N(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__a2bb2o_1 _08225_ (.A1_N(_02150_),
    .A2_N(_02151_),
    .B1(_02158_),
    .B2(_02159_),
    .X(_02161_));
 sky130_fd_sc_hd__a21oi_1 _08226_ (.A1(_02160_),
    .A2(_02161_),
    .B1(_02149_),
    .Y(_02162_));
 sky130_fd_sc_hd__nand3_1 _08227_ (.A(_02149_),
    .B(_02160_),
    .C(_02161_),
    .Y(_02163_));
 sky130_fd_sc_hd__nand2b_1 _08228_ (.A_N(_02162_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__xor2_1 _08229_ (.A(_02148_),
    .B(_02164_),
    .X(_02166_));
 sky130_fd_sc_hd__a21o_1 _08230_ (.A1(_02131_),
    .A2(_02133_),
    .B1(_02096_),
    .X(_02167_));
 sky130_fd_sc_hd__nand3_2 _08231_ (.A(_02166_),
    .B(_02167_),
    .C(_02134_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _08232_ (.A(_02158_),
    .B(_02160_),
    .Y(_02169_));
 sky130_fd_sc_hd__nand4_2 _08233_ (.A(net37),
    .B(net36),
    .C(net23),
    .D(net12),
    .Y(_02170_));
 sky130_fd_sc_hd__a22o_1 _08234_ (.A1(net36),
    .A2(net23),
    .B1(net12),
    .B2(net37),
    .X(_02171_));
 sky130_fd_sc_hd__nand4_2 _08235_ (.A(_02171_),
    .B(net1),
    .C(net38),
    .D(_02170_),
    .Y(_02172_));
 sky130_fd_sc_hd__a22o_1 _08236_ (.A1(net38),
    .A2(net1),
    .B1(_02170_),
    .B2(_02171_),
    .X(_02173_));
 sky130_fd_sc_hd__nand2_1 _08237_ (.A(_02153_),
    .B(_02156_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand4_2 _08238_ (.A(net34),
    .B(net64),
    .C(net28),
    .D(net27),
    .Y(_02175_));
 sky130_fd_sc_hd__a22o_1 _08239_ (.A1(net64),
    .A2(net28),
    .B1(net27),
    .B2(net34),
    .X(_02177_));
 sky130_fd_sc_hd__nand4_2 _08240_ (.A(_02177_),
    .B(net26),
    .C(net35),
    .D(_02175_),
    .Y(_02178_));
 sky130_fd_sc_hd__a22o_1 _08241_ (.A1(net35),
    .A2(net26),
    .B1(_02175_),
    .B2(_02177_),
    .X(_02179_));
 sky130_fd_sc_hd__and3_1 _08242_ (.A(_02174_),
    .B(_02178_),
    .C(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__nand3_1 _08243_ (.A(_02174_),
    .B(_02178_),
    .C(_02179_),
    .Y(_02181_));
 sky130_fd_sc_hd__a21o_1 _08244_ (.A1(_02178_),
    .A2(_02179_),
    .B1(_02174_),
    .X(_02182_));
 sky130_fd_sc_hd__nand4_1 _08245_ (.A(_02172_),
    .B(_02173_),
    .C(_02181_),
    .D(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__a22o_1 _08246_ (.A1(_02172_),
    .A2(_02173_),
    .B1(_02181_),
    .B2(_02182_),
    .X(_02184_));
 sky130_fd_sc_hd__a211o_1 _08247_ (.A1(_02183_),
    .A2(_02184_),
    .B1(_02106_),
    .C1(_02107_),
    .X(_02185_));
 sky130_fd_sc_hd__o211ai_1 _08248_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_02183_),
    .C1(_02184_),
    .Y(_02186_));
 sky130_fd_sc_hd__and3_1 _08249_ (.A(_02169_),
    .B(_02185_),
    .C(_02186_),
    .X(_02188_));
 sky130_fd_sc_hd__a21oi_1 _08250_ (.A1(_02185_),
    .A2(_02186_),
    .B1(_02169_),
    .Y(_02189_));
 sky130_fd_sc_hd__nand2_1 _08251_ (.A(_02129_),
    .B(_02131_),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _08252_ (.A(_02112_),
    .B(_02113_),
    .Y(_02191_));
 sky130_fd_sc_hd__or4b_4 _08253_ (.A(_01153_),
    .B(_01164_),
    .C(_01175_),
    .D_N(net61),
    .X(_02192_));
 sky130_fd_sc_hd__a22o_1 _08254_ (.A1(net62),
    .A2(net30),
    .B1(net61),
    .B2(net31),
    .X(_02193_));
 sky130_fd_sc_hd__nand4_4 _08255_ (.A(_02193_),
    .B(net29),
    .C(net63),
    .D(_02192_),
    .Y(_02194_));
 sky130_fd_sc_hd__a22o_1 _08256_ (.A1(net63),
    .A2(net29),
    .B1(_02192_),
    .B2(_02193_),
    .X(_02195_));
 sky130_fd_sc_hd__a21o_1 _08257_ (.A1(_02194_),
    .A2(_02195_),
    .B1(_02191_),
    .X(_02196_));
 sky130_fd_sc_hd__nand3_1 _08258_ (.A(_02191_),
    .B(_02194_),
    .C(_02195_),
    .Y(_02197_));
 sky130_fd_sc_hd__o211a_1 _08259_ (.A1(_02098_),
    .A2(_02102_),
    .B1(_02196_),
    .C1(_02197_),
    .X(_02199_));
 sky130_fd_sc_hd__a211oi_1 _08260_ (.A1(_02196_),
    .A2(_02197_),
    .B1(_02098_),
    .C1(_02102_),
    .Y(_02200_));
 sky130_fd_sc_hd__o21ai_1 _08261_ (.A1(_02115_),
    .A2(_02125_),
    .B1(_02124_),
    .Y(_02201_));
 sky130_fd_sc_hd__a22o_1 _08262_ (.A1(net2),
    .A2(net59),
    .B1(net58),
    .B2(net3),
    .X(_02202_));
 sky130_fd_sc_hd__nand4_2 _08263_ (.A(net3),
    .B(net2),
    .C(net59),
    .D(net58),
    .Y(_02203_));
 sky130_fd_sc_hd__nand4_2 _08264_ (.A(_02202_),
    .B(_02203_),
    .C(net32),
    .D(net60),
    .Y(_02204_));
 sky130_fd_sc_hd__a22o_1 _08265_ (.A1(net32),
    .A2(net60),
    .B1(_02202_),
    .B2(_02203_),
    .X(_02205_));
 sky130_fd_sc_hd__a31o_1 _08266_ (.A1(_02120_),
    .A2(net55),
    .A3(net3),
    .B1(_02118_),
    .X(_02206_));
 sky130_fd_sc_hd__nand2_1 _08267_ (.A(net6),
    .B(net33),
    .Y(_02207_));
 sky130_fd_sc_hd__nand4_1 _08268_ (.A(net6),
    .B(net5),
    .C(net44),
    .D(net33),
    .Y(_02208_));
 sky130_fd_sc_hd__a22o_1 _08269_ (.A1(net5),
    .A2(net44),
    .B1(net33),
    .B2(net6),
    .X(_02210_));
 sky130_fd_sc_hd__nand4_2 _08270_ (.A(_02210_),
    .B(net55),
    .C(net4),
    .D(_02208_),
    .Y(_02211_));
 sky130_fd_sc_hd__a22o_1 _08271_ (.A1(net4),
    .A2(net55),
    .B1(_02208_),
    .B2(_02210_),
    .X(_02212_));
 sky130_fd_sc_hd__nand3_2 _08272_ (.A(_02206_),
    .B(_02211_),
    .C(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__a21o_1 _08273_ (.A1(_02211_),
    .A2(_02212_),
    .B1(_02206_),
    .X(_02214_));
 sky130_fd_sc_hd__nand4_2 _08274_ (.A(_02204_),
    .B(_02205_),
    .C(_02213_),
    .D(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__a22o_1 _08275_ (.A1(_02204_),
    .A2(_02205_),
    .B1(_02213_),
    .B2(_02214_),
    .X(_02216_));
 sky130_fd_sc_hd__nand3_1 _08276_ (.A(_02201_),
    .B(_02215_),
    .C(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__a21o_1 _08277_ (.A1(_02215_),
    .A2(_02216_),
    .B1(_02201_),
    .X(_02218_));
 sky130_fd_sc_hd__or4bb_2 _08278_ (.A(_02199_),
    .B(_02200_),
    .C_N(_02217_),
    .D_N(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__a2bb2o_1 _08279_ (.A1_N(_02199_),
    .A2_N(_02200_),
    .B1(_02217_),
    .B2(_02218_),
    .X(_02221_));
 sky130_fd_sc_hd__nand3_2 _08280_ (.A(_02190_),
    .B(_02219_),
    .C(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__a21o_1 _08281_ (.A1(_02219_),
    .A2(_02221_),
    .B1(_02190_),
    .X(_02223_));
 sky130_fd_sc_hd__or4bb_1 _08282_ (.A(_02188_),
    .B(_02189_),
    .C_N(_02222_),
    .D_N(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__a211o_1 _08283_ (.A1(_02222_),
    .A2(_02223_),
    .B1(_02188_),
    .C1(_02189_),
    .X(_02225_));
 sky130_fd_sc_hd__o211ai_2 _08284_ (.A1(_02188_),
    .A2(_02189_),
    .B1(_02222_),
    .C1(_02223_),
    .Y(_02226_));
 sky130_fd_sc_hd__a22oi_2 _08285_ (.A1(_02134_),
    .A2(_02168_),
    .B1(_02225_),
    .B2(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__o21ai_1 _08286_ (.A1(_02148_),
    .A2(_02162_),
    .B1(_02163_),
    .Y(_02228_));
 sky130_fd_sc_hd__and2_1 _08287_ (.A(_02228_),
    .B(_02150_),
    .X(_02229_));
 sky130_fd_sc_hd__xor2_1 _08288_ (.A(_02150_),
    .B(_02228_),
    .X(_02230_));
 sky130_fd_sc_hd__nand4_1 _08289_ (.A(_02134_),
    .B(_02168_),
    .C(_02225_),
    .D(_02226_),
    .Y(_02232_));
 sky130_fd_sc_hd__and2b_1 _08290_ (.A_N(_02227_),
    .B(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__a21o_1 _08291_ (.A1(_02232_),
    .A2(_02230_),
    .B1(_02227_),
    .X(_02234_));
 sky130_fd_sc_hd__a21bo_1 _08292_ (.A1(_02169_),
    .A2(_02185_),
    .B1_N(_02186_),
    .X(_02235_));
 sky130_fd_sc_hd__nand2_1 _08293_ (.A(_02170_),
    .B(_02172_),
    .Y(_02236_));
 sky130_fd_sc_hd__and3_1 _08294_ (.A(_02236_),
    .B(net1),
    .C(net39),
    .X(_02237_));
 sky130_fd_sc_hd__a21oi_1 _08295_ (.A1(net39),
    .A2(net1),
    .B1(_02236_),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_1 _08296_ (.A(_02237_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _08297_ (.A(_02239_),
    .B(_02235_),
    .Y(_02240_));
 sky130_fd_sc_hd__and2_1 _08298_ (.A(_02235_),
    .B(_02239_),
    .X(_02241_));
 sky130_fd_sc_hd__nor2_1 _08299_ (.A(_02240_),
    .B(_02241_),
    .Y(_02243_));
 sky130_fd_sc_hd__a31o_1 _08300_ (.A1(_02172_),
    .A2(_02173_),
    .A3(_02182_),
    .B1(_02180_),
    .X(_02244_));
 sky130_fd_sc_hd__a31oi_1 _08301_ (.A1(_02191_),
    .A2(_02194_),
    .A3(_02195_),
    .B1(_02199_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand4_2 _08302_ (.A(net37),
    .B(net36),
    .C(net26),
    .D(net23),
    .Y(_02246_));
 sky130_fd_sc_hd__a22o_1 _08303_ (.A1(net36),
    .A2(net26),
    .B1(net23),
    .B2(net37),
    .X(_02247_));
 sky130_fd_sc_hd__nand4_2 _08304_ (.A(_02247_),
    .B(net12),
    .C(net38),
    .D(_02246_),
    .Y(_02248_));
 sky130_fd_sc_hd__a22o_1 _08305_ (.A1(net38),
    .A2(net12),
    .B1(_02246_),
    .B2(_02247_),
    .X(_02249_));
 sky130_fd_sc_hd__nand2_1 _08306_ (.A(_02175_),
    .B(_02178_),
    .Y(_02250_));
 sky130_fd_sc_hd__nand4_1 _08307_ (.A(net34),
    .B(net64),
    .C(net29),
    .D(net28),
    .Y(_02251_));
 sky130_fd_sc_hd__a22o_1 _08308_ (.A1(net64),
    .A2(net29),
    .B1(net28),
    .B2(net34),
    .X(_02252_));
 sky130_fd_sc_hd__nand4_1 _08309_ (.A(_02252_),
    .B(net27),
    .C(net35),
    .D(_02251_),
    .Y(_02254_));
 sky130_fd_sc_hd__a22o_1 _08310_ (.A1(net35),
    .A2(net27),
    .B1(_02251_),
    .B2(_02252_),
    .X(_02255_));
 sky130_fd_sc_hd__and3_1 _08311_ (.A(_02250_),
    .B(_02254_),
    .C(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__a21oi_1 _08312_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02250_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _08313_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__and3_1 _08314_ (.A(_02258_),
    .B(_02249_),
    .C(_02248_),
    .X(_02259_));
 sky130_fd_sc_hd__o211ai_1 _08315_ (.A1(_02256_),
    .A2(_02257_),
    .B1(_02248_),
    .C1(_02249_),
    .Y(_02260_));
 sky130_fd_sc_hd__a211o_1 _08316_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02256_),
    .C1(_02257_),
    .X(_02261_));
 sky130_fd_sc_hd__nand3_1 _08317_ (.A(_02245_),
    .B(_02260_),
    .C(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__a21o_1 _08318_ (.A1(_02260_),
    .A2(_02261_),
    .B1(_02245_),
    .X(_02263_));
 sky130_fd_sc_hd__nand3_2 _08319_ (.A(_02244_),
    .B(_02262_),
    .C(_02263_),
    .Y(_02265_));
 sky130_fd_sc_hd__a21o_1 _08320_ (.A1(_02262_),
    .A2(_02263_),
    .B1(_02244_),
    .X(_02266_));
 sky130_fd_sc_hd__nand2_1 _08321_ (.A(_02265_),
    .B(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__nand2_1 _08322_ (.A(_02203_),
    .B(_02204_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand4_2 _08323_ (.A(net32),
    .B(net31),
    .C(net62),
    .D(net61),
    .Y(_02269_));
 sky130_fd_sc_hd__a22o_1 _08324_ (.A1(net31),
    .A2(net62),
    .B1(net61),
    .B2(net32),
    .X(_02270_));
 sky130_fd_sc_hd__nand4_2 _08325_ (.A(_02270_),
    .B(net30),
    .C(net63),
    .D(_02269_),
    .Y(_02271_));
 sky130_fd_sc_hd__a22o_1 _08326_ (.A1(net63),
    .A2(net30),
    .B1(_02269_),
    .B2(_02270_),
    .X(_02272_));
 sky130_fd_sc_hd__a21oi_2 _08327_ (.A1(_02271_),
    .A2(_02272_),
    .B1(_02268_),
    .Y(_02273_));
 sky130_fd_sc_hd__and3_2 _08328_ (.A(_02268_),
    .B(_02271_),
    .C(_02272_),
    .X(_02274_));
 sky130_fd_sc_hd__a211oi_4 _08329_ (.A1(_02192_),
    .A2(_02194_),
    .B1(_02273_),
    .C1(_02274_),
    .Y(_02276_));
 sky130_fd_sc_hd__o211a_1 _08330_ (.A1(_02273_),
    .A2(_02274_),
    .B1(_02192_),
    .C1(_02194_),
    .X(_02277_));
 sky130_fd_sc_hd__nand2_1 _08331_ (.A(_02213_),
    .B(_02215_),
    .Y(_02278_));
 sky130_fd_sc_hd__a22o_1 _08332_ (.A1(net3),
    .A2(net59),
    .B1(net58),
    .B2(net4),
    .X(_02279_));
 sky130_fd_sc_hd__nand4_1 _08333_ (.A(net4),
    .B(net3),
    .C(net59),
    .D(net58),
    .Y(_02280_));
 sky130_fd_sc_hd__o2bb2a_1 _08334_ (.A1_N(_02279_),
    .A2_N(_02280_),
    .B1(_01131_),
    .B2(_01197_),
    .X(_02281_));
 sky130_fd_sc_hd__and4_1 _08335_ (.A(_02279_),
    .B(_02280_),
    .C(net2),
    .D(net60),
    .X(_02282_));
 sky130_fd_sc_hd__nor2_1 _08336_ (.A(_02281_),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__o21ai_1 _08337_ (.A1(_02117_),
    .A2(_02207_),
    .B1(_02211_),
    .Y(_02284_));
 sky130_fd_sc_hd__and4_1 _08338_ (.A(net7),
    .B(net6),
    .C(net44),
    .D(net33),
    .X(_02285_));
 sky130_fd_sc_hd__or2_1 _08339_ (.A(_01916_),
    .B(_02207_),
    .X(_02287_));
 sky130_fd_sc_hd__a22o_1 _08340_ (.A1(net6),
    .A2(net44),
    .B1(net33),
    .B2(net7),
    .X(_02288_));
 sky130_fd_sc_hd__and2_1 _08341_ (.A(net5),
    .B(net55),
    .X(_02289_));
 sky130_fd_sc_hd__o2111ai_4 _08342_ (.A1(_01916_),
    .A2(_02207_),
    .B1(net5),
    .C1(net55),
    .D1(_02288_),
    .Y(_02290_));
 sky130_fd_sc_hd__a22o_1 _08343_ (.A1(net5),
    .A2(net55),
    .B1(_02287_),
    .B2(_02288_),
    .X(_02291_));
 sky130_fd_sc_hd__and3_1 _08344_ (.A(_02284_),
    .B(_02290_),
    .C(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__nand3_1 _08345_ (.A(_02284_),
    .B(_02290_),
    .C(_02291_),
    .Y(_02293_));
 sky130_fd_sc_hd__a21oi_1 _08346_ (.A1(_02290_),
    .A2(_02291_),
    .B1(_02284_),
    .Y(_02294_));
 sky130_fd_sc_hd__a21o_1 _08347_ (.A1(_02290_),
    .A2(_02291_),
    .B1(_02284_),
    .X(_02295_));
 sky130_fd_sc_hd__nand3_1 _08348_ (.A(_02295_),
    .B(_02283_),
    .C(_02293_),
    .Y(_02296_));
 sky130_fd_sc_hd__a2bb2o_1 _08349_ (.A1_N(_02281_),
    .A2_N(_02282_),
    .B1(_02293_),
    .B2(_02295_),
    .X(_02298_));
 sky130_fd_sc_hd__a211o_1 _08350_ (.A1(_02293_),
    .A2(_02295_),
    .B1(_02281_),
    .C1(_02282_),
    .X(_02299_));
 sky130_fd_sc_hd__or3_1 _08351_ (.A(_02283_),
    .B(_02292_),
    .C(_02294_),
    .X(_02300_));
 sky130_fd_sc_hd__a22o_1 _08352_ (.A1(_02213_),
    .A2(_02215_),
    .B1(_02299_),
    .B2(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__and4_1 _08353_ (.A(_02213_),
    .B(_02215_),
    .C(_02299_),
    .D(_02300_),
    .X(_02302_));
 sky130_fd_sc_hd__a21o_1 _08354_ (.A1(_02296_),
    .A2(_02298_),
    .B1(_02278_),
    .X(_02303_));
 sky130_fd_sc_hd__a211o_1 _08355_ (.A1(_02301_),
    .A2(_02303_),
    .B1(_02276_),
    .C1(_02277_),
    .X(_02304_));
 sky130_fd_sc_hd__o211ai_2 _08356_ (.A1(_02276_),
    .A2(_02277_),
    .B1(_02301_),
    .C1(_02303_),
    .Y(_02305_));
 sky130_fd_sc_hd__a22oi_1 _08357_ (.A1(_02217_),
    .A2(_02219_),
    .B1(_02304_),
    .B2(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__a22o_1 _08358_ (.A1(_02217_),
    .A2(_02219_),
    .B1(_02304_),
    .B2(_02305_),
    .X(_02307_));
 sky130_fd_sc_hd__nand4_1 _08359_ (.A(_02217_),
    .B(_02219_),
    .C(_02304_),
    .D(_02305_),
    .Y(_02309_));
 sky130_fd_sc_hd__a21o_1 _08360_ (.A1(_02307_),
    .A2(_02309_),
    .B1(_02267_),
    .X(_02310_));
 sky130_fd_sc_hd__nand3_1 _08361_ (.A(_02267_),
    .B(_02307_),
    .C(_02309_),
    .Y(_02311_));
 sky130_fd_sc_hd__a22o_1 _08362_ (.A1(_02222_),
    .A2(_02224_),
    .B1(_02310_),
    .B2(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__nand4_1 _08363_ (.A(_02222_),
    .B(_02224_),
    .C(_02310_),
    .D(_02311_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand3_1 _08364_ (.A(_02312_),
    .B(_02313_),
    .C(_02243_),
    .Y(_02314_));
 sky130_fd_sc_hd__a21o_1 _08365_ (.A1(_02312_),
    .A2(_02313_),
    .B1(_02243_),
    .X(_02315_));
 sky130_fd_sc_hd__nand3_1 _08366_ (.A(_02234_),
    .B(_02314_),
    .C(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__a221o_1 _08367_ (.A1(_02232_),
    .A2(_02230_),
    .B1(_02315_),
    .B2(_02314_),
    .C1(_02227_),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_1 _08368_ (.A(_02316_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__a21boi_1 _08369_ (.A1(_02317_),
    .A2(_02229_),
    .B1_N(_02316_),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_2 _08370_ (.A(_02312_),
    .B(_02314_),
    .Y(_02321_));
 sky130_fd_sc_hd__and4_1 _08371_ (.A(net40),
    .B(net39),
    .C(net12),
    .D(net1),
    .X(_02322_));
 sky130_fd_sc_hd__nand4_1 _08372_ (.A(net40),
    .B(net39),
    .C(net12),
    .D(net1),
    .Y(_02323_));
 sky130_fd_sc_hd__a22oi_1 _08373_ (.A1(net39),
    .A2(net12),
    .B1(net1),
    .B2(net40),
    .Y(_02324_));
 sky130_fd_sc_hd__a211o_1 _08374_ (.A1(_02246_),
    .A2(_02248_),
    .B1(_02322_),
    .C1(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__o211ai_1 _08375_ (.A1(_02322_),
    .A2(_02324_),
    .B1(_02246_),
    .C1(_02248_),
    .Y(_02326_));
 sky130_fd_sc_hd__and3_1 _08376_ (.A(_02237_),
    .B(_02325_),
    .C(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__a21oi_1 _08377_ (.A1(_02325_),
    .A2(_02326_),
    .B1(_02237_),
    .Y(_02328_));
 sky130_fd_sc_hd__o211a_1 _08378_ (.A1(_02327_),
    .A2(_02328_),
    .B1(_02263_),
    .C1(_02265_),
    .X(_02329_));
 sky130_fd_sc_hd__a211oi_2 _08379_ (.A1(_02263_),
    .A2(_02265_),
    .B1(_02327_),
    .C1(_02328_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_1 _08380_ (.A(_02329_),
    .B(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__a31o_1 _08381_ (.A1(_02265_),
    .A2(_02266_),
    .A3(_02309_),
    .B1(_02306_),
    .X(_02333_));
 sky130_fd_sc_hd__a31o_1 _08382_ (.A1(_02268_),
    .A2(_02271_),
    .A3(_02272_),
    .B1(_02276_),
    .X(_02334_));
 sky130_fd_sc_hd__nand4_2 _08383_ (.A(net37),
    .B(net36),
    .C(net27),
    .D(net26),
    .Y(_02335_));
 sky130_fd_sc_hd__a22o_1 _08384_ (.A1(net36),
    .A2(net27),
    .B1(net26),
    .B2(net37),
    .X(_02336_));
 sky130_fd_sc_hd__nand4_2 _08385_ (.A(_02336_),
    .B(net23),
    .C(net38),
    .D(_02335_),
    .Y(_02337_));
 sky130_fd_sc_hd__a22o_1 _08386_ (.A1(net38),
    .A2(net23),
    .B1(_02335_),
    .B2(_02336_),
    .X(_02338_));
 sky130_fd_sc_hd__nand2_1 _08387_ (.A(_02251_),
    .B(_02254_),
    .Y(_02339_));
 sky130_fd_sc_hd__nand4_1 _08388_ (.A(net34),
    .B(net64),
    .C(net30),
    .D(net29),
    .Y(_02340_));
 sky130_fd_sc_hd__a22o_1 _08389_ (.A1(net64),
    .A2(net30),
    .B1(net29),
    .B2(net34),
    .X(_02342_));
 sky130_fd_sc_hd__nand4_1 _08390_ (.A(_02342_),
    .B(net28),
    .C(net35),
    .D(_02340_),
    .Y(_02343_));
 sky130_fd_sc_hd__a22o_1 _08391_ (.A1(net35),
    .A2(net28),
    .B1(_02340_),
    .B2(_02342_),
    .X(_02344_));
 sky130_fd_sc_hd__nand3_1 _08392_ (.A(_02339_),
    .B(_02343_),
    .C(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__a21o_1 _08393_ (.A1(_02343_),
    .A2(_02344_),
    .B1(_02339_),
    .X(_02346_));
 sky130_fd_sc_hd__nand4_2 _08394_ (.A(_02337_),
    .B(_02338_),
    .C(_02345_),
    .D(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__a22o_1 _08395_ (.A1(_02337_),
    .A2(_02338_),
    .B1(_02345_),
    .B2(_02346_),
    .X(_02348_));
 sky130_fd_sc_hd__a211o_1 _08396_ (.A1(_02347_),
    .A2(_02348_),
    .B1(_02274_),
    .C1(_02276_),
    .X(_02349_));
 sky130_fd_sc_hd__o211ai_1 _08397_ (.A1(_02274_),
    .A2(_02276_),
    .B1(_02347_),
    .C1(_02348_),
    .Y(_02350_));
 sky130_fd_sc_hd__o211a_1 _08398_ (.A1(_02256_),
    .A2(_02259_),
    .B1(_02349_),
    .C1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__a211oi_1 _08399_ (.A1(_02349_),
    .A2(_02350_),
    .B1(_02256_),
    .C1(_02259_),
    .Y(_02353_));
 sky130_fd_sc_hd__o31ai_1 _08400_ (.A1(_02276_),
    .A2(_02277_),
    .A3(_02302_),
    .B1(_02301_),
    .Y(_02354_));
 sky130_fd_sc_hd__a41o_1 _08401_ (.A1(net4),
    .A2(net3),
    .A3(net59),
    .A4(net58),
    .B1(_02282_),
    .X(_02355_));
 sky130_fd_sc_hd__nand4_1 _08402_ (.A(net2),
    .B(net32),
    .C(net62),
    .D(net61),
    .Y(_02356_));
 sky130_fd_sc_hd__a22o_1 _08403_ (.A1(net32),
    .A2(net62),
    .B1(net61),
    .B2(net2),
    .X(_02357_));
 sky130_fd_sc_hd__nand4_1 _08404_ (.A(_02357_),
    .B(net31),
    .C(net63),
    .D(_02356_),
    .Y(_02358_));
 sky130_fd_sc_hd__a22o_1 _08405_ (.A1(net63),
    .A2(net31),
    .B1(_02356_),
    .B2(_02357_),
    .X(_02359_));
 sky130_fd_sc_hd__a21oi_1 _08406_ (.A1(_02358_),
    .A2(_02359_),
    .B1(_02355_),
    .Y(_02360_));
 sky130_fd_sc_hd__and3_1 _08407_ (.A(_02355_),
    .B(_02358_),
    .C(_02359_),
    .X(_02361_));
 sky130_fd_sc_hd__a211oi_1 _08408_ (.A1(_02269_),
    .A2(_02271_),
    .B1(_02360_),
    .C1(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__o211a_1 _08409_ (.A1(_02360_),
    .A2(_02361_),
    .B1(_02269_),
    .C1(_02271_),
    .X(_02364_));
 sky130_fd_sc_hd__a22o_1 _08410_ (.A1(net4),
    .A2(net59),
    .B1(net58),
    .B2(net5),
    .X(_02365_));
 sky130_fd_sc_hd__nand4_2 _08411_ (.A(net5),
    .B(net4),
    .C(net59),
    .D(net58),
    .Y(_02366_));
 sky130_fd_sc_hd__a22o_1 _08412_ (.A1(net3),
    .A2(net60),
    .B1(_02365_),
    .B2(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__nand4_2 _08413_ (.A(_02365_),
    .B(_02366_),
    .C(net3),
    .D(net60),
    .Y(_02368_));
 sky130_fd_sc_hd__a21o_1 _08414_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_02285_),
    .X(_02369_));
 sky130_fd_sc_hd__nand3b_1 _08415_ (.A_N(_01917_),
    .B(_01919_),
    .C(_01920_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand3_2 _08416_ (.A(_01921_),
    .B(_02369_),
    .C(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__a21o_1 _08417_ (.A1(_01921_),
    .A2(_02370_),
    .B1(_02369_),
    .X(_02372_));
 sky130_fd_sc_hd__nand4_2 _08418_ (.A(_02367_),
    .B(_02368_),
    .C(_02371_),
    .D(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__a22o_1 _08419_ (.A1(_02367_),
    .A2(_02368_),
    .B1(_02371_),
    .B2(_02372_),
    .X(_02375_));
 sky130_fd_sc_hd__nand2_1 _08420_ (.A(_02373_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _08421_ (.A1(_02293_),
    .A2(_02296_),
    .B1(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__a221o_1 _08422_ (.A1(_02295_),
    .A2(_02283_),
    .B1(_02375_),
    .B2(_02373_),
    .C1(_02292_),
    .X(_02378_));
 sky130_fd_sc_hd__or4bb_2 _08423_ (.A(_02362_),
    .B(_02364_),
    .C_N(_02377_),
    .D_N(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__a2bb2o_1 _08424_ (.A1_N(_02362_),
    .A2_N(_02364_),
    .B1(_02377_),
    .B2(_02378_),
    .X(_02380_));
 sky130_fd_sc_hd__nand3_1 _08425_ (.A(_02354_),
    .B(_02379_),
    .C(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__a21o_1 _08426_ (.A1(_02379_),
    .A2(_02380_),
    .B1(_02354_),
    .X(_02382_));
 sky130_fd_sc_hd__or4bb_2 _08427_ (.A(_02351_),
    .B(_02353_),
    .C_N(_02381_),
    .D_N(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__a2bb2o_1 _08428_ (.A1_N(_02351_),
    .A2_N(_02353_),
    .B1(_02381_),
    .B2(_02382_),
    .X(_02384_));
 sky130_fd_sc_hd__nand3_1 _08429_ (.A(_02333_),
    .B(_02383_),
    .C(_02384_),
    .Y(_02386_));
 sky130_fd_sc_hd__a21o_1 _08430_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_02333_),
    .X(_02387_));
 sky130_fd_sc_hd__nand3_1 _08431_ (.A(_02387_),
    .B(_02332_),
    .C(_02386_),
    .Y(_02388_));
 sky130_fd_sc_hd__a21o_1 _08432_ (.A1(_02386_),
    .A2(_02387_),
    .B1(_02332_),
    .X(_02389_));
 sky130_fd_sc_hd__and2_2 _08433_ (.A(_02388_),
    .B(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__xor2_2 _08434_ (.A(_02321_),
    .B(_02390_),
    .X(_02391_));
 sky130_fd_sc_hd__xnor2_1 _08435_ (.A(_02241_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__nand2_1 _08436_ (.A(net31),
    .B(net44),
    .Y(_02393_));
 sky130_fd_sc_hd__nand4_1 _08437_ (.A(net32),
    .B(net31),
    .C(net44),
    .D(net33),
    .Y(_02394_));
 sky130_fd_sc_hd__nand2_1 _08438_ (.A(net30),
    .B(net55),
    .Y(_02395_));
 sky130_fd_sc_hd__a22oi_1 _08439_ (.A1(net31),
    .A2(net44),
    .B1(net33),
    .B2(net32),
    .Y(_02397_));
 sky130_fd_sc_hd__nand3_1 _08440_ (.A(_02393_),
    .B(net33),
    .C(net32),
    .Y(_02398_));
 sky130_fd_sc_hd__nand3_1 _08441_ (.A(_02031_),
    .B(net44),
    .C(net31),
    .Y(_02399_));
 sky130_fd_sc_hd__nand4b_1 _08442_ (.A_N(_02397_),
    .B(net55),
    .C(net30),
    .D(_02394_),
    .Y(_02400_));
 sky130_fd_sc_hd__o21ai_1 _08443_ (.A1(_02395_),
    .A2(_02397_),
    .B1(_02394_),
    .Y(_02401_));
 sky130_fd_sc_hd__o211ai_2 _08444_ (.A1(_01153_),
    .A2(_01230_),
    .B1(_02036_),
    .C1(_02037_),
    .Y(_02402_));
 sky130_fd_sc_hd__and3_1 _08445_ (.A(_02038_),
    .B(_02401_),
    .C(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__a22o_1 _08446_ (.A1(net29),
    .A2(net59),
    .B1(net58),
    .B2(net30),
    .X(_02404_));
 sky130_fd_sc_hd__nand4_2 _08447_ (.A(net30),
    .B(net29),
    .C(net59),
    .D(net58),
    .Y(_02405_));
 sky130_fd_sc_hd__nand4_2 _08448_ (.A(_02404_),
    .B(_02405_),
    .C(net60),
    .D(net28),
    .Y(_02406_));
 sky130_fd_sc_hd__a22o_1 _08449_ (.A1(net60),
    .A2(net28),
    .B1(_02404_),
    .B2(_02405_),
    .X(_02408_));
 sky130_fd_sc_hd__a21oi_1 _08450_ (.A1(_02038_),
    .A2(_02402_),
    .B1(_02401_),
    .Y(_02409_));
 sky130_fd_sc_hd__a21o_1 _08451_ (.A1(_02038_),
    .A2(_02402_),
    .B1(_02401_),
    .X(_02410_));
 sky130_fd_sc_hd__a31o_1 _08452_ (.A1(_02406_),
    .A2(_02408_),
    .A3(_02410_),
    .B1(_02403_),
    .X(_02411_));
 sky130_fd_sc_hd__a22o_1 _08453_ (.A1(_02052_),
    .A2(_02053_),
    .B1(_02054_),
    .B2(_02048_),
    .X(_02412_));
 sky130_fd_sc_hd__and3_1 _08454_ (.A(_02056_),
    .B(_02411_),
    .C(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__nand3_1 _08455_ (.A(_02056_),
    .B(_02411_),
    .C(_02412_),
    .Y(_02414_));
 sky130_fd_sc_hd__nand4_4 _08456_ (.A(net62),
    .B(net61),
    .C(net27),
    .D(net26),
    .Y(_02415_));
 sky130_fd_sc_hd__a22o_1 _08457_ (.A1(net61),
    .A2(net27),
    .B1(net26),
    .B2(net62),
    .X(_02416_));
 sky130_fd_sc_hd__nand4_4 _08458_ (.A(_02416_),
    .B(net23),
    .C(net63),
    .D(_02415_),
    .Y(_02417_));
 sky130_fd_sc_hd__nand2_1 _08459_ (.A(_02405_),
    .B(_02406_),
    .Y(_02419_));
 sky130_fd_sc_hd__a22o_1 _08460_ (.A1(net63),
    .A2(net26),
    .B1(_02076_),
    .B2(_02078_),
    .X(_02420_));
 sky130_fd_sc_hd__a21oi_1 _08461_ (.A1(_02079_),
    .A2(_02420_),
    .B1(_02419_),
    .Y(_02421_));
 sky130_fd_sc_hd__and3_1 _08462_ (.A(_02079_),
    .B(_02419_),
    .C(_02420_),
    .X(_02422_));
 sky130_fd_sc_hd__nand3_1 _08463_ (.A(_02079_),
    .B(_02419_),
    .C(_02420_),
    .Y(_02423_));
 sky130_fd_sc_hd__a211o_1 _08464_ (.A1(_02415_),
    .A2(_02417_),
    .B1(_02421_),
    .C1(_02422_),
    .X(_02424_));
 sky130_fd_sc_hd__o211ai_1 _08465_ (.A1(_02421_),
    .A2(_02422_),
    .B1(_02415_),
    .C1(_02417_),
    .Y(_02425_));
 sky130_fd_sc_hd__nand2_1 _08466_ (.A(_02424_),
    .B(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__a21o_1 _08467_ (.A1(_02056_),
    .A2(_02412_),
    .B1(_02411_),
    .X(_02427_));
 sky130_fd_sc_hd__a31o_1 _08468_ (.A1(_02424_),
    .A2(_02425_),
    .A3(_02427_),
    .B1(_02413_),
    .X(_02428_));
 sky130_fd_sc_hd__a22o_1 _08469_ (.A1(_02092_),
    .A2(_02093_),
    .B1(_02094_),
    .B2(_02074_),
    .X(_02430_));
 sky130_fd_sc_hd__nand3_1 _08470_ (.A(_02095_),
    .B(_02428_),
    .C(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__nand2_1 _08471_ (.A(net64),
    .B(net1),
    .Y(_02432_));
 sky130_fd_sc_hd__and4_1 _08472_ (.A(net34),
    .B(net64),
    .C(net12),
    .D(net1),
    .X(_02433_));
 sky130_fd_sc_hd__o22a_1 _08473_ (.A1(_01109_),
    .A2(_01263_),
    .B1(_02135_),
    .B2(_02136_),
    .X(_02434_));
 sky130_fd_sc_hd__nor3b_2 _08474_ (.A(_02137_),
    .B(_02434_),
    .C_N(_02433_),
    .Y(_02435_));
 sky130_fd_sc_hd__a21o_1 _08475_ (.A1(_02144_),
    .A2(_02147_),
    .B1(_02145_),
    .X(_02436_));
 sky130_fd_sc_hd__nand3_1 _08476_ (.A(_02144_),
    .B(_02145_),
    .C(_02147_),
    .Y(_02437_));
 sky130_fd_sc_hd__nand4_1 _08477_ (.A(_02423_),
    .B(_02424_),
    .C(_02436_),
    .D(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__a22o_1 _08478_ (.A1(_02423_),
    .A2(_02424_),
    .B1(_02436_),
    .B2(_02437_),
    .X(_02439_));
 sky130_fd_sc_hd__a21o_1 _08479_ (.A1(_02438_),
    .A2(_02439_),
    .B1(_02435_),
    .X(_02441_));
 sky130_fd_sc_hd__nand3_1 _08480_ (.A(_02438_),
    .B(_02439_),
    .C(_02435_),
    .Y(_02442_));
 sky130_fd_sc_hd__a21o_1 _08481_ (.A1(_02095_),
    .A2(_02430_),
    .B1(_02428_),
    .X(_02443_));
 sky130_fd_sc_hd__and4_1 _08482_ (.A(_02431_),
    .B(_02441_),
    .C(_02442_),
    .D(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__a31o_1 _08483_ (.A1(_02095_),
    .A2(_02428_),
    .A3(_02430_),
    .B1(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__a21o_1 _08484_ (.A1(_02134_),
    .A2(_02167_),
    .B1(_02166_),
    .X(_02446_));
 sky130_fd_sc_hd__nand3_1 _08485_ (.A(_02168_),
    .B(_02445_),
    .C(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__a21o_1 _08486_ (.A1(_02168_),
    .A2(_02446_),
    .B1(_02445_),
    .X(_02448_));
 sky130_fd_sc_hd__nand2_1 _08487_ (.A(_02447_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__and2_1 _08488_ (.A(_02439_),
    .B(_02442_),
    .X(_02450_));
 sky130_fd_sc_hd__a21o_1 _08489_ (.A1(_02439_),
    .A2(_02442_),
    .B1(_02449_),
    .X(_02452_));
 sky130_fd_sc_hd__xnor2_1 _08490_ (.A(_02230_),
    .B(_02233_),
    .Y(_02453_));
 sky130_fd_sc_hd__a21o_1 _08491_ (.A1(_02447_),
    .A2(_02452_),
    .B1(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__xor2_1 _08492_ (.A(_02229_),
    .B(_02318_),
    .X(_02455_));
 sky130_fd_sc_hd__o22a_1 _08493_ (.A1(_02454_),
    .A2(_02455_),
    .B1(_02320_),
    .B2(_02392_),
    .X(_02456_));
 sky130_fd_sc_hd__nand4_2 _08494_ (.A(net59),
    .B(net27),
    .C(net58),
    .D(net26),
    .Y(_02457_));
 sky130_fd_sc_hd__a22o_1 _08495_ (.A1(net27),
    .A2(net58),
    .B1(net26),
    .B2(net59),
    .X(_02458_));
 sky130_fd_sc_hd__nand4_2 _08496_ (.A(_02458_),
    .B(net23),
    .C(net60),
    .D(_02457_),
    .Y(_02459_));
 sky130_fd_sc_hd__nand2_1 _08497_ (.A(_02457_),
    .B(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__nand4_2 _08498_ (.A(net62),
    .B(net61),
    .C(net23),
    .D(net12),
    .Y(_02461_));
 sky130_fd_sc_hd__a22o_1 _08499_ (.A1(net61),
    .A2(net23),
    .B1(net12),
    .B2(net62),
    .X(_02463_));
 sky130_fd_sc_hd__nand4_2 _08500_ (.A(_02463_),
    .B(net1),
    .C(net63),
    .D(_02461_),
    .Y(_02464_));
 sky130_fd_sc_hd__a22o_1 _08501_ (.A1(net63),
    .A2(net1),
    .B1(_02461_),
    .B2(_02463_),
    .X(_02465_));
 sky130_fd_sc_hd__nand3_1 _08502_ (.A(_02460_),
    .B(_02464_),
    .C(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__and4_2 _08503_ (.A(net62),
    .B(net61),
    .C(net12),
    .D(net1),
    .X(_02467_));
 sky130_fd_sc_hd__a21o_1 _08504_ (.A1(_02464_),
    .A2(_02465_),
    .B1(_02460_),
    .X(_02468_));
 sky130_fd_sc_hd__and3_1 _08505_ (.A(_02466_),
    .B(_02468_),
    .C(_02467_),
    .X(_02469_));
 sky130_fd_sc_hd__a31oi_2 _08506_ (.A1(_02460_),
    .A2(_02464_),
    .A3(_02465_),
    .B1(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_2 _08507_ (.A(net28),
    .B(net44),
    .Y(_02471_));
 sky130_fd_sc_hd__and4_1 _08508_ (.A(net29),
    .B(net28),
    .C(net44),
    .D(net33),
    .X(_02472_));
 sky130_fd_sc_hd__nand4_2 _08509_ (.A(net29),
    .B(net28),
    .C(net44),
    .D(net33),
    .Y(_02474_));
 sky130_fd_sc_hd__a22o_1 _08510_ (.A1(net28),
    .A2(net44),
    .B1(net33),
    .B2(net29),
    .X(_02475_));
 sky130_fd_sc_hd__and4_2 _08511_ (.A(_02475_),
    .B(net55),
    .C(net27),
    .D(_02474_),
    .X(_02476_));
 sky130_fd_sc_hd__a31o_1 _08512_ (.A1(_02475_),
    .A2(net55),
    .A3(net27),
    .B1(_02472_),
    .X(_02477_));
 sky130_fd_sc_hd__and4_1 _08513_ (.A(net30),
    .B(net29),
    .C(net44),
    .D(net33),
    .X(_02478_));
 sky130_fd_sc_hd__nand4_1 _08514_ (.A(net30),
    .B(net29),
    .C(net44),
    .D(net33),
    .Y(_02479_));
 sky130_fd_sc_hd__a22o_1 _08515_ (.A1(net29),
    .A2(net44),
    .B1(net33),
    .B2(net30),
    .X(_02480_));
 sky130_fd_sc_hd__nand4_2 _08516_ (.A(_02480_),
    .B(net55),
    .C(net28),
    .D(_02479_),
    .Y(_02481_));
 sky130_fd_sc_hd__a22o_1 _08517_ (.A1(net28),
    .A2(net55),
    .B1(_02479_),
    .B2(_02480_),
    .X(_02482_));
 sky130_fd_sc_hd__o211ai_4 _08518_ (.A1(_02472_),
    .A2(_02476_),
    .B1(_02481_),
    .C1(_02482_),
    .Y(_02483_));
 sky130_fd_sc_hd__a22o_1 _08519_ (.A1(net60),
    .A2(net23),
    .B1(_02457_),
    .B2(_02458_),
    .X(_02485_));
 sky130_fd_sc_hd__nand2_1 _08520_ (.A(_02459_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__a21oi_1 _08521_ (.A1(_02481_),
    .A2(_02482_),
    .B1(_02477_),
    .Y(_02487_));
 sky130_fd_sc_hd__a21o_1 _08522_ (.A1(_02481_),
    .A2(_02482_),
    .B1(_02477_),
    .X(_02488_));
 sky130_fd_sc_hd__nor3b_1 _08523_ (.A(_02486_),
    .B(_02487_),
    .C_N(_02483_),
    .Y(_02489_));
 sky130_fd_sc_hd__o21ai_2 _08524_ (.A1(_02486_),
    .A2(_02487_),
    .B1(_02483_),
    .Y(_02490_));
 sky130_fd_sc_hd__a22o_1 _08525_ (.A1(net59),
    .A2(net27),
    .B1(net58),
    .B2(net28),
    .X(_02491_));
 sky130_fd_sc_hd__nand4_2 _08526_ (.A(net28),
    .B(net59),
    .C(net27),
    .D(net58),
    .Y(_02492_));
 sky130_fd_sc_hd__nand4_2 _08527_ (.A(_02491_),
    .B(_02492_),
    .C(net60),
    .D(net26),
    .Y(_02493_));
 sky130_fd_sc_hd__a22o_1 _08528_ (.A1(net60),
    .A2(net26),
    .B1(_02491_),
    .B2(_02492_),
    .X(_02494_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(_02493_),
    .B(_02494_),
    .Y(_02496_));
 sky130_fd_sc_hd__a31o_1 _08530_ (.A1(_02480_),
    .A2(net55),
    .A3(net28),
    .B1(_02478_),
    .X(_02497_));
 sky130_fd_sc_hd__nand4_2 _08531_ (.A(net31),
    .B(net30),
    .C(net44),
    .D(net33),
    .Y(_02498_));
 sky130_fd_sc_hd__a22oi_1 _08532_ (.A1(net30),
    .A2(net44),
    .B1(net33),
    .B2(net31),
    .Y(_02499_));
 sky130_fd_sc_hd__a22o_1 _08533_ (.A1(net30),
    .A2(net44),
    .B1(net33),
    .B2(net31),
    .X(_02500_));
 sky130_fd_sc_hd__nand4_1 _08534_ (.A(_02500_),
    .B(net55),
    .C(net29),
    .D(_02498_),
    .Y(_02501_));
 sky130_fd_sc_hd__o2bb2ai_1 _08535_ (.A1_N(_02498_),
    .A2_N(_02500_),
    .B1(_01186_),
    .B2(_01230_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand3_1 _08536_ (.A(_02497_),
    .B(_02501_),
    .C(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__a21oi_1 _08537_ (.A1(_02501_),
    .A2(_02502_),
    .B1(_02497_),
    .Y(_02504_));
 sky130_fd_sc_hd__a21o_1 _08538_ (.A1(_02501_),
    .A2(_02502_),
    .B1(_02497_),
    .X(_02505_));
 sky130_fd_sc_hd__nand4_1 _08539_ (.A(_02493_),
    .B(_02494_),
    .C(_02503_),
    .D(_02505_),
    .Y(_02507_));
 sky130_fd_sc_hd__a22o_1 _08540_ (.A1(_02493_),
    .A2(_02494_),
    .B1(_02503_),
    .B2(_02505_),
    .X(_02508_));
 sky130_fd_sc_hd__nand3_2 _08541_ (.A(_02490_),
    .B(_02507_),
    .C(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__a21oi_1 _08542_ (.A1(_02466_),
    .A2(_02468_),
    .B1(_02467_),
    .Y(_02510_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_02469_),
    .B(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__a21o_1 _08544_ (.A1(_02507_),
    .A2(_02508_),
    .B1(_02490_),
    .X(_02512_));
 sky130_fd_sc_hd__nand3_1 _08545_ (.A(_02511_),
    .B(_02512_),
    .C(_02509_),
    .Y(_02513_));
 sky130_fd_sc_hd__nand2_1 _08546_ (.A(_02461_),
    .B(_02464_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand2_1 _08547_ (.A(_02492_),
    .B(_02493_),
    .Y(_02515_));
 sky130_fd_sc_hd__and4_1 _08548_ (.A(net62),
    .B(net61),
    .C(net26),
    .D(net23),
    .X(_02516_));
 sky130_fd_sc_hd__nand4_1 _08549_ (.A(net62),
    .B(net61),
    .C(net26),
    .D(net23),
    .Y(_02518_));
 sky130_fd_sc_hd__a22o_1 _08550_ (.A1(net61),
    .A2(net26),
    .B1(net23),
    .B2(net62),
    .X(_02519_));
 sky130_fd_sc_hd__and4_1 _08551_ (.A(_02519_),
    .B(net12),
    .C(net63),
    .D(_02518_),
    .X(_02520_));
 sky130_fd_sc_hd__nand4_1 _08552_ (.A(_02519_),
    .B(net12),
    .C(net63),
    .D(_02518_),
    .Y(_02521_));
 sky130_fd_sc_hd__a22o_1 _08553_ (.A1(net63),
    .A2(net12),
    .B1(_02518_),
    .B2(_02519_),
    .X(_02522_));
 sky130_fd_sc_hd__a21o_1 _08554_ (.A1(_02521_),
    .A2(_02522_),
    .B1(_02515_),
    .X(_02523_));
 sky130_fd_sc_hd__nand3_2 _08555_ (.A(_02515_),
    .B(_02521_),
    .C(_02522_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand3_2 _08556_ (.A(_02514_),
    .B(_02523_),
    .C(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__a21o_1 _08557_ (.A1(_02523_),
    .A2(_02524_),
    .B1(_02514_),
    .X(_02526_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(_02525_),
    .B(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__o21ai_1 _08559_ (.A1(_02496_),
    .A2(_02504_),
    .B1(_02503_),
    .Y(_02529_));
 sky130_fd_sc_hd__a22o_1 _08560_ (.A1(net28),
    .A2(net59),
    .B1(net58),
    .B2(net29),
    .X(_02530_));
 sky130_fd_sc_hd__and4_1 _08561_ (.A(net29),
    .B(net28),
    .C(net59),
    .D(net58),
    .X(_02531_));
 sky130_fd_sc_hd__nand4_1 _08562_ (.A(net29),
    .B(net28),
    .C(net59),
    .D(net58),
    .Y(_02532_));
 sky130_fd_sc_hd__o2bb2a_1 _08563_ (.A1_N(_02530_),
    .A2_N(_02532_),
    .B1(_01197_),
    .B2(_01208_),
    .X(_02533_));
 sky130_fd_sc_hd__and4_2 _08564_ (.A(_02530_),
    .B(_02532_),
    .C(net60),
    .D(net27),
    .X(_02534_));
 sky130_fd_sc_hd__nor2_1 _08565_ (.A(_02533_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__o31ai_2 _08566_ (.A1(_01186_),
    .A2(_01230_),
    .A3(_02499_),
    .B1(_02498_),
    .Y(_02536_));
 sky130_fd_sc_hd__o211ai_2 _08567_ (.A1(_01175_),
    .A2(_01230_),
    .B1(_02398_),
    .C1(_02399_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand3_2 _08568_ (.A(_02400_),
    .B(_02536_),
    .C(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__a21o_1 _08569_ (.A1(_02400_),
    .A2(_02537_),
    .B1(_02536_),
    .X(_02540_));
 sky130_fd_sc_hd__nand3_2 _08570_ (.A(_02540_),
    .B(_02535_),
    .C(_02538_),
    .Y(_02541_));
 sky130_fd_sc_hd__a2bb2o_1 _08571_ (.A1_N(_02533_),
    .A2_N(_02534_),
    .B1(_02538_),
    .B2(_02540_),
    .X(_02542_));
 sky130_fd_sc_hd__and3_1 _08572_ (.A(_02529_),
    .B(_02541_),
    .C(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__nand3_1 _08573_ (.A(_02529_),
    .B(_02541_),
    .C(_02542_),
    .Y(_02544_));
 sky130_fd_sc_hd__a21o_1 _08574_ (.A1(_02541_),
    .A2(_02542_),
    .B1(_02529_),
    .X(_02545_));
 sky130_fd_sc_hd__a21o_1 _08575_ (.A1(_02544_),
    .A2(_02545_),
    .B1(_02527_),
    .X(_02546_));
 sky130_fd_sc_hd__nand3_1 _08576_ (.A(_02527_),
    .B(_02544_),
    .C(_02545_),
    .Y(_02547_));
 sky130_fd_sc_hd__a22o_1 _08577_ (.A1(_02509_),
    .A2(_02513_),
    .B1(_02546_),
    .B2(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__xor2_2 _08578_ (.A(_02432_),
    .B(_02470_),
    .X(_02549_));
 sky130_fd_sc_hd__nand4_1 _08579_ (.A(_02509_),
    .B(_02513_),
    .C(_02546_),
    .D(_02547_),
    .Y(_02551_));
 sky130_fd_sc_hd__nand2_1 _08580_ (.A(_02548_),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__a21bo_1 _08581_ (.A1(_02549_),
    .A2(_02551_),
    .B1_N(_02548_),
    .X(_02553_));
 sky130_fd_sc_hd__a22oi_2 _08582_ (.A1(net64),
    .A2(net12),
    .B1(net1),
    .B2(net34),
    .Y(_02554_));
 sky130_fd_sc_hd__a211oi_2 _08583_ (.A1(_02524_),
    .A2(_02525_),
    .B1(_02554_),
    .C1(_02433_),
    .Y(_02555_));
 sky130_fd_sc_hd__o211a_1 _08584_ (.A1(_02433_),
    .A2(_02554_),
    .B1(_02525_),
    .C1(_02524_),
    .X(_02556_));
 sky130_fd_sc_hd__nor2_1 _08585_ (.A(_02555_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__a31o_1 _08586_ (.A1(_02525_),
    .A2(_02526_),
    .A3(_02545_),
    .B1(_02543_),
    .X(_02558_));
 sky130_fd_sc_hd__a31o_1 _08587_ (.A1(_02519_),
    .A2(net12),
    .A3(net63),
    .B1(_02516_),
    .X(_02559_));
 sky130_fd_sc_hd__a22o_1 _08588_ (.A1(net63),
    .A2(net23),
    .B1(_02415_),
    .B2(_02416_),
    .X(_02560_));
 sky130_fd_sc_hd__a211o_1 _08589_ (.A1(_02417_),
    .A2(_02560_),
    .B1(_02534_),
    .C1(_02531_),
    .X(_02562_));
 sky130_fd_sc_hd__o211ai_4 _08590_ (.A1(_02531_),
    .A2(_02534_),
    .B1(_02560_),
    .C1(_02417_),
    .Y(_02563_));
 sky130_fd_sc_hd__and3_1 _08591_ (.A(_02559_),
    .B(_02562_),
    .C(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__o211ai_2 _08592_ (.A1(_02516_),
    .A2(_02520_),
    .B1(_02562_),
    .C1(_02563_),
    .Y(_02565_));
 sky130_fd_sc_hd__a21oi_1 _08593_ (.A1(_02562_),
    .A2(_02563_),
    .B1(_02559_),
    .Y(_02566_));
 sky130_fd_sc_hd__a211o_1 _08594_ (.A1(_02562_),
    .A2(_02563_),
    .B1(_02516_),
    .C1(_02520_),
    .X(_02567_));
 sky130_fd_sc_hd__o211ai_1 _08595_ (.A1(_02403_),
    .A2(_02409_),
    .B1(_02408_),
    .C1(_02406_),
    .Y(_02568_));
 sky130_fd_sc_hd__a211o_1 _08596_ (.A1(_02406_),
    .A2(_02408_),
    .B1(_02409_),
    .C1(_02403_),
    .X(_02569_));
 sky130_fd_sc_hd__a22o_1 _08597_ (.A1(_02538_),
    .A2(_02541_),
    .B1(_02568_),
    .B2(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__nand4_1 _08598_ (.A(_02538_),
    .B(_02541_),
    .C(_02568_),
    .D(_02569_),
    .Y(_02571_));
 sky130_fd_sc_hd__nand4_1 _08599_ (.A(_02565_),
    .B(_02567_),
    .C(_02570_),
    .D(_02571_),
    .Y(_02573_));
 sky130_fd_sc_hd__a2bb2o_1 _08600_ (.A1_N(_02564_),
    .A2_N(_02566_),
    .B1(_02570_),
    .B2(_02571_),
    .X(_02574_));
 sky130_fd_sc_hd__nand3_1 _08601_ (.A(_02558_),
    .B(_02573_),
    .C(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__a21o_1 _08602_ (.A1(_02573_),
    .A2(_02574_),
    .B1(_02558_),
    .X(_02576_));
 sky130_fd_sc_hd__a211o_1 _08603_ (.A1(_02575_),
    .A2(_02576_),
    .B1(_02555_),
    .C1(_02556_),
    .X(_02577_));
 sky130_fd_sc_hd__o211ai_1 _08604_ (.A1(_02555_),
    .A2(_02556_),
    .B1(_02575_),
    .C1(_02576_),
    .Y(_02578_));
 sky130_fd_sc_hd__a21bo_1 _08605_ (.A1(_02577_),
    .A2(_02578_),
    .B1_N(_02553_),
    .X(_02579_));
 sky130_fd_sc_hd__nand3b_1 _08606_ (.A_N(_02553_),
    .B(_02577_),
    .C(_02578_),
    .Y(_02580_));
 sky130_fd_sc_hd__or4bb_2 _08607_ (.A(_02432_),
    .B(_02470_),
    .C_N(_02579_),
    .D_N(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__a2bb2o_1 _08608_ (.A1_N(_02470_),
    .A2_N(_02432_),
    .B1(_02580_),
    .B2(_02579_),
    .X(_02582_));
 sky130_fd_sc_hd__nand2_2 _08609_ (.A(net27),
    .B(net33),
    .Y(_02584_));
 sky130_fd_sc_hd__or2_1 _08610_ (.A(_02471_),
    .B(_02584_),
    .X(_02585_));
 sky130_fd_sc_hd__a22o_1 _08611_ (.A1(net27),
    .A2(net44),
    .B1(net33),
    .B2(net28),
    .X(_02586_));
 sky130_fd_sc_hd__o2111ai_4 _08612_ (.A1(_02471_),
    .A2(_02584_),
    .B1(net26),
    .C1(net55),
    .D1(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__a22oi_4 _08613_ (.A1(net27),
    .A2(net55),
    .B1(_02474_),
    .B2(_02475_),
    .Y(_02588_));
 sky130_fd_sc_hd__a21o_1 _08614_ (.A1(_02585_),
    .A2(_02587_),
    .B1(_02476_),
    .X(_02589_));
 sky130_fd_sc_hd__a211oi_1 _08615_ (.A1(_02585_),
    .A2(_02587_),
    .B1(_02588_),
    .C1(_02476_),
    .Y(_02590_));
 sky130_fd_sc_hd__a211o_1 _08616_ (.A1(_02585_),
    .A2(_02587_),
    .B1(_02588_),
    .C1(_02476_),
    .X(_02591_));
 sky130_fd_sc_hd__a22o_1 _08617_ (.A1(net58),
    .A2(net26),
    .B1(net23),
    .B2(net59),
    .X(_02592_));
 sky130_fd_sc_hd__nand4_4 _08618_ (.A(net59),
    .B(net58),
    .C(net26),
    .D(net23),
    .Y(_02593_));
 sky130_fd_sc_hd__nand4_4 _08619_ (.A(_02592_),
    .B(_02593_),
    .C(net60),
    .D(net12),
    .Y(_02595_));
 sky130_fd_sc_hd__a22o_1 _08620_ (.A1(net60),
    .A2(net12),
    .B1(_02592_),
    .B2(_02593_),
    .X(_02596_));
 sky130_fd_sc_hd__o221ai_4 _08621_ (.A1(_02471_),
    .A2(_02584_),
    .B1(_02588_),
    .B2(_02476_),
    .C1(_02587_),
    .Y(_02597_));
 sky130_fd_sc_hd__o2111ai_4 _08622_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02595_),
    .C1(_02596_),
    .D1(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__a31o_1 _08623_ (.A1(_02595_),
    .A2(_02596_),
    .A3(_02597_),
    .B1(_02590_),
    .X(_02599_));
 sky130_fd_sc_hd__a22oi_2 _08624_ (.A1(_02459_),
    .A2(_02485_),
    .B1(_02488_),
    .B2(_02483_),
    .Y(_02600_));
 sky130_fd_sc_hd__a22o_1 _08625_ (.A1(_02459_),
    .A2(_02485_),
    .B1(_02488_),
    .B2(_02483_),
    .X(_02601_));
 sky130_fd_sc_hd__nand3b_2 _08626_ (.A_N(_02489_),
    .B(_02599_),
    .C(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__o2bb2a_1 _08627_ (.A1_N(net61),
    .A2_N(net12),
    .B1(_01263_),
    .B2(_01164_),
    .X(_02603_));
 sky130_fd_sc_hd__a211oi_4 _08628_ (.A1(_02593_),
    .A2(_02595_),
    .B1(_02603_),
    .C1(_02467_),
    .Y(_02604_));
 sky130_fd_sc_hd__inv_2 _08629_ (.A(_02604_),
    .Y(_02606_));
 sky130_fd_sc_hd__o211a_1 _08630_ (.A1(_02467_),
    .A2(_02603_),
    .B1(_02595_),
    .C1(_02593_),
    .X(_02607_));
 sky130_fd_sc_hd__o221ai_4 _08631_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02600_),
    .B2(_02489_),
    .C1(_02598_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(_02602_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__or3_1 _08633_ (.A(_02604_),
    .B(_02607_),
    .C(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__a211o_1 _08634_ (.A1(_02509_),
    .A2(_02512_),
    .B1(_02510_),
    .C1(_02469_),
    .X(_02611_));
 sky130_fd_sc_hd__o211ai_2 _08635_ (.A1(_02469_),
    .A2(_02510_),
    .B1(_02512_),
    .C1(_02509_),
    .Y(_02612_));
 sky130_fd_sc_hd__a22o_1 _08636_ (.A1(_02602_),
    .A2(_02610_),
    .B1(_02611_),
    .B2(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__nand4_2 _08637_ (.A(_02602_),
    .B(_02610_),
    .C(_02611_),
    .D(_02612_),
    .Y(_02614_));
 sky130_fd_sc_hd__nand3_1 _08638_ (.A(_02613_),
    .B(_02614_),
    .C(_02604_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _08639_ (.A(_02613_),
    .B(_02615_),
    .Y(_02617_));
 sky130_fd_sc_hd__xnor2_2 _08640_ (.A(_02549_),
    .B(_02552_),
    .Y(_02618_));
 sky130_fd_sc_hd__nand4_1 _08641_ (.A(_02582_),
    .B(_02618_),
    .C(_02617_),
    .D(_02581_),
    .Y(_02619_));
 sky130_fd_sc_hd__a22o_1 _08642_ (.A1(_02618_),
    .A2(_02617_),
    .B1(_02582_),
    .B2(_02581_),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_1 _08643_ (.A(_02619_),
    .B(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__nand4_1 _08644_ (.A(net27),
    .B(net26),
    .C(net44),
    .D(net33),
    .Y(_02622_));
 sky130_fd_sc_hd__a22o_1 _08645_ (.A1(net26),
    .A2(net44),
    .B1(net33),
    .B2(net27),
    .X(_02623_));
 sky130_fd_sc_hd__and4_1 _08646_ (.A(_02623_),
    .B(net55),
    .C(net23),
    .D(_02622_),
    .X(_02624_));
 sky130_fd_sc_hd__a41o_1 _08647_ (.A1(net27),
    .A2(net26),
    .A3(net44),
    .A4(net33),
    .B1(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__a22o_1 _08648_ (.A1(net26),
    .A2(net55),
    .B1(_02585_),
    .B2(_02586_),
    .X(_02626_));
 sky130_fd_sc_hd__and3_1 _08649_ (.A(_02587_),
    .B(_02625_),
    .C(_02626_),
    .X(_02628_));
 sky130_fd_sc_hd__a22o_1 _08650_ (.A1(net58),
    .A2(net23),
    .B1(net12),
    .B2(net59),
    .X(_02629_));
 sky130_fd_sc_hd__and4_1 _08651_ (.A(net59),
    .B(net58),
    .C(net23),
    .D(net12),
    .X(_02630_));
 sky130_fd_sc_hd__nand4_1 _08652_ (.A(net59),
    .B(net58),
    .C(net23),
    .D(net12),
    .Y(_02631_));
 sky130_fd_sc_hd__and4_1 _08653_ (.A(_02629_),
    .B(_02631_),
    .C(net60),
    .D(net1),
    .X(_02632_));
 sky130_fd_sc_hd__o2bb2a_1 _08654_ (.A1_N(_02629_),
    .A2_N(_02631_),
    .B1(_01197_),
    .B2(_01263_),
    .X(_02633_));
 sky130_fd_sc_hd__or2_1 _08655_ (.A(_02632_),
    .B(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__a21oi_1 _08656_ (.A1(_02587_),
    .A2(_02626_),
    .B1(_02625_),
    .Y(_02635_));
 sky130_fd_sc_hd__o21bai_1 _08657_ (.A1(_02634_),
    .A2(_02635_),
    .B1_N(_02628_),
    .Y(_02636_));
 sky130_fd_sc_hd__a22o_1 _08658_ (.A1(_02595_),
    .A2(_02596_),
    .B1(_02597_),
    .B2(_02591_),
    .X(_02637_));
 sky130_fd_sc_hd__nand3_1 _08659_ (.A(_02598_),
    .B(_02636_),
    .C(_02637_),
    .Y(_02639_));
 sky130_fd_sc_hd__a211oi_1 _08660_ (.A1(net61),
    .A2(net1),
    .B1(_02630_),
    .C1(_02632_),
    .Y(_02640_));
 sky130_fd_sc_hd__o211a_1 _08661_ (.A1(_02630_),
    .A2(_02632_),
    .B1(net61),
    .C1(net1),
    .X(_02641_));
 sky130_fd_sc_hd__nor2_1 _08662_ (.A(_02640_),
    .B(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__a21o_1 _08663_ (.A1(_02598_),
    .A2(_02637_),
    .B1(_02636_),
    .X(_02643_));
 sky130_fd_sc_hd__and3_1 _08664_ (.A(_02639_),
    .B(_02643_),
    .C(_02642_),
    .X(_02644_));
 sky130_fd_sc_hd__a21boi_1 _08665_ (.A1(_02643_),
    .A2(_02642_),
    .B1_N(_02639_),
    .Y(_02645_));
 sky130_fd_sc_hd__a211o_1 _08666_ (.A1(_02602_),
    .A2(_02608_),
    .B1(_02607_),
    .C1(_02604_),
    .X(_02646_));
 sky130_fd_sc_hd__o211ai_1 _08667_ (.A1(_02604_),
    .A2(_02607_),
    .B1(_02608_),
    .C1(_02602_),
    .Y(_02647_));
 sky130_fd_sc_hd__a21o_1 _08668_ (.A1(_02646_),
    .A2(_02647_),
    .B1(_02645_),
    .X(_02648_));
 sky130_fd_sc_hd__nand3_1 _08669_ (.A(_02646_),
    .B(_02647_),
    .C(_02645_),
    .Y(_02650_));
 sky130_fd_sc_hd__and3_1 _08670_ (.A(_02648_),
    .B(_02650_),
    .C(_02641_),
    .X(_02651_));
 sky130_fd_sc_hd__a21bo_1 _08671_ (.A1(_02641_),
    .A2(_02650_),
    .B1_N(_02648_),
    .X(_02652_));
 sky130_fd_sc_hd__a21o_1 _08672_ (.A1(_02613_),
    .A2(_02614_),
    .B1(_02604_),
    .X(_02653_));
 sky130_fd_sc_hd__a21oi_1 _08673_ (.A1(_02613_),
    .A2(_02614_),
    .B1(_02606_),
    .Y(_02654_));
 sky130_fd_sc_hd__and3_1 _08674_ (.A(_02606_),
    .B(_02613_),
    .C(_02614_),
    .X(_02655_));
 sky130_fd_sc_hd__o21ai_1 _08675_ (.A1(_02654_),
    .A2(_02655_),
    .B1(_02652_),
    .Y(_02656_));
 sky130_fd_sc_hd__xnor2_2 _08676_ (.A(_02617_),
    .B(_02618_),
    .Y(_02657_));
 sky130_fd_sc_hd__a21oi_1 _08677_ (.A1(_02648_),
    .A2(_02650_),
    .B1(_02641_),
    .Y(_02658_));
 sky130_fd_sc_hd__a311oi_1 _08678_ (.A1(_02615_),
    .A2(_02652_),
    .A3(_02653_),
    .B1(_02658_),
    .C1(_02651_),
    .Y(_02659_));
 sky130_fd_sc_hd__o31ai_1 _08679_ (.A1(_02652_),
    .A2(_02654_),
    .A3(_02655_),
    .B1(_02659_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand4_2 _08680_ (.A(net26),
    .B(net23),
    .C(net44),
    .D(net33),
    .Y(_02662_));
 sky130_fd_sc_hd__a22o_1 _08681_ (.A1(net23),
    .A2(net44),
    .B1(net33),
    .B2(net26),
    .X(_02663_));
 sky130_fd_sc_hd__and4_1 _08682_ (.A(_02663_),
    .B(net12),
    .C(net55),
    .D(_02662_),
    .X(_02664_));
 sky130_fd_sc_hd__nand4_1 _08683_ (.A(_02663_),
    .B(net12),
    .C(net55),
    .D(_02662_),
    .Y(_02665_));
 sky130_fd_sc_hd__a22oi_1 _08684_ (.A1(net23),
    .A2(net55),
    .B1(_02622_),
    .B2(_02623_),
    .Y(_02666_));
 sky130_fd_sc_hd__a211o_1 _08685_ (.A1(_02662_),
    .A2(_02665_),
    .B1(_02666_),
    .C1(_02624_),
    .X(_02667_));
 sky130_fd_sc_hd__a22oi_1 _08686_ (.A1(net58),
    .A2(net12),
    .B1(net1),
    .B2(net59),
    .Y(_02668_));
 sky130_fd_sc_hd__and4_1 _08687_ (.A(net59),
    .B(net58),
    .C(net12),
    .D(net1),
    .X(_02669_));
 sky130_fd_sc_hd__nor2_1 _08688_ (.A(_02668_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__o211ai_1 _08689_ (.A1(_02624_),
    .A2(_02666_),
    .B1(_02665_),
    .C1(_02662_),
    .Y(_02672_));
 sky130_fd_sc_hd__and2_1 _08690_ (.A(_02667_),
    .B(_02672_),
    .X(_02673_));
 sky130_fd_sc_hd__a21bo_1 _08691_ (.A1(_02670_),
    .A2(_02672_),
    .B1_N(_02667_),
    .X(_02674_));
 sky130_fd_sc_hd__o21ai_1 _08692_ (.A1(_02628_),
    .A2(_02635_),
    .B1(_02634_),
    .Y(_02675_));
 sky130_fd_sc_hd__o41a_1 _08693_ (.A1(_02628_),
    .A2(_02632_),
    .A3(_02633_),
    .A4(_02635_),
    .B1(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_1 _08694_ (.A(_02676_),
    .B(_02674_),
    .Y(_02677_));
 sky130_fd_sc_hd__xor2_1 _08695_ (.A(_02674_),
    .B(_02676_),
    .X(_02678_));
 sky130_fd_sc_hd__nand2_1 _08696_ (.A(_02669_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__a21oi_1 _08697_ (.A1(_02639_),
    .A2(_02643_),
    .B1(_02642_),
    .Y(_02680_));
 sky130_fd_sc_hd__or2_1 _08698_ (.A(_02644_),
    .B(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__a21o_1 _08699_ (.A1(_02677_),
    .A2(_02679_),
    .B1(_02681_),
    .X(_02683_));
 sky130_fd_sc_hd__o22a_1 _08700_ (.A1(_02656_),
    .A2(_02657_),
    .B1(_02661_),
    .B2(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__o2bb2a_1 _08701_ (.A1_N(_02662_),
    .A2_N(_02663_),
    .B1(_01230_),
    .B2(_01241_),
    .X(_02685_));
 sky130_fd_sc_hd__and4_1 _08702_ (.A(net23),
    .B(net12),
    .C(net44),
    .D(net33),
    .X(_02686_));
 sky130_fd_sc_hd__a22o_1 _08703_ (.A1(net12),
    .A2(net44),
    .B1(net33),
    .B2(net23),
    .X(_02687_));
 sky130_fd_sc_hd__and2b_1 _08704_ (.A_N(_02686_),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__a31o_1 _08705_ (.A1(_02687_),
    .A2(net1),
    .A3(net55),
    .B1(_02686_),
    .X(_02689_));
 sky130_fd_sc_hd__or3b_1 _08706_ (.A(_02664_),
    .B(_02685_),
    .C_N(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__o21bai_1 _08707_ (.A1(_02664_),
    .A2(_02685_),
    .B1_N(_02689_),
    .Y(_02691_));
 sky130_fd_sc_hd__and2_1 _08708_ (.A(_02690_),
    .B(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__nand4_1 _08709_ (.A(_02690_),
    .B(_02691_),
    .C(net58),
    .D(net1),
    .Y(_02694_));
 sky130_fd_sc_hd__and2_1 _08710_ (.A(_02690_),
    .B(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__xnor2_1 _08711_ (.A(_02670_),
    .B(_02673_),
    .Y(_02696_));
 sky130_fd_sc_hd__o2111a_1 _08712_ (.A1(net23),
    .A2(_01230_),
    .B1(net12),
    .C1(net44),
    .D1(net33),
    .X(_02697_));
 sky130_fd_sc_hd__o2111a_1 _08713_ (.A1(net55),
    .A2(_02688_),
    .B1(_02697_),
    .C1(net1),
    .D1(_02694_),
    .X(_02698_));
 sky130_fd_sc_hd__o21ai_1 _08714_ (.A1(net58),
    .A2(_02692_),
    .B1(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__a21o_1 _08715_ (.A1(_02695_),
    .A2(_02696_),
    .B1(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__o22a_1 _08716_ (.A1(_02695_),
    .A2(_02696_),
    .B1(_02700_),
    .B2(_02657_),
    .X(_02701_));
 sky130_fd_sc_hd__nand3_1 _08717_ (.A(_02677_),
    .B(_02679_),
    .C(_02681_),
    .Y(_02702_));
 sky130_fd_sc_hd__o2bb2a_1 _08718_ (.A1_N(_02669_),
    .A2_N(_02678_),
    .B1(_02681_),
    .B2(_02677_),
    .X(_02703_));
 sky130_fd_sc_hd__a21boi_1 _08719_ (.A1(_02576_),
    .A2(_02557_),
    .B1_N(_02575_),
    .Y(_02705_));
 sky130_fd_sc_hd__o21ba_1 _08720_ (.A1(_02137_),
    .A2(_02434_),
    .B1_N(_02433_),
    .X(_02706_));
 sky130_fd_sc_hd__a211oi_2 _08721_ (.A1(_02563_),
    .A2(_02565_),
    .B1(_02706_),
    .C1(_02435_),
    .Y(_02707_));
 sky130_fd_sc_hd__o211a_1 _08722_ (.A1(_02435_),
    .A2(_02706_),
    .B1(_02565_),
    .C1(_02563_),
    .X(_02708_));
 sky130_fd_sc_hd__nor2_1 _08723_ (.A(_02707_),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__nand2_1 _08724_ (.A(_02570_),
    .B(_02573_),
    .Y(_02710_));
 sky130_fd_sc_hd__a21oi_1 _08725_ (.A1(_02414_),
    .A2(_02427_),
    .B1(_02426_),
    .Y(_02711_));
 sky130_fd_sc_hd__and3_1 _08726_ (.A(_02414_),
    .B(_02426_),
    .C(_02427_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_1 _08727_ (.A1(_02711_),
    .A2(_02712_),
    .B1(_02710_),
    .Y(_02713_));
 sky130_fd_sc_hd__or3_1 _08728_ (.A(_02711_),
    .B(_02712_),
    .C(_02710_),
    .X(_02714_));
 sky130_fd_sc_hd__a211o_1 _08729_ (.A1(_02713_),
    .A2(_02714_),
    .B1(_02707_),
    .C1(_02708_),
    .X(_02716_));
 sky130_fd_sc_hd__o211ai_1 _08730_ (.A1(_02707_),
    .A2(_02708_),
    .B1(_02713_),
    .C1(_02714_),
    .Y(_02717_));
 sky130_fd_sc_hd__a21o_1 _08731_ (.A1(_02716_),
    .A2(_02717_),
    .B1(_02705_),
    .X(_02718_));
 sky130_fd_sc_hd__nand3_1 _08732_ (.A(_02705_),
    .B(_02716_),
    .C(_02717_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand3_1 _08733_ (.A(_02718_),
    .B(_02719_),
    .C(_02555_),
    .Y(_02720_));
 sky130_fd_sc_hd__a21o_1 _08734_ (.A1(_02718_),
    .A2(_02719_),
    .B1(_02555_),
    .X(_02721_));
 sky130_fd_sc_hd__nand2_1 _08735_ (.A(_02720_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__and2_1 _08736_ (.A(_02579_),
    .B(_02581_),
    .X(_02723_));
 sky130_fd_sc_hd__nand2_1 _08737_ (.A(_02579_),
    .B(_02581_),
    .Y(_02724_));
 sky130_fd_sc_hd__a21o_1 _08738_ (.A1(_02579_),
    .A2(_02581_),
    .B1(_02722_),
    .X(_02725_));
 sky130_fd_sc_hd__a21o_1 _08739_ (.A1(_02720_),
    .A2(_02721_),
    .B1(_02724_),
    .X(_02727_));
 sky130_fd_sc_hd__nand2_1 _08740_ (.A(_02725_),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__o21ba_1 _08741_ (.A1(_02695_),
    .A2(_02696_),
    .B1_N(_02700_),
    .X(_02729_));
 sky130_fd_sc_hd__nor3_1 _08742_ (.A(_02656_),
    .B(_02729_),
    .C(_02657_),
    .Y(_02730_));
 sky130_fd_sc_hd__o21ai_1 _08743_ (.A1(_02684_),
    .A2(_02730_),
    .B1(_02621_),
    .Y(_02731_));
 sky130_fd_sc_hd__a22o_1 _08744_ (.A1(_02656_),
    .A2(_02657_),
    .B1(_02728_),
    .B2(_02619_),
    .X(_02732_));
 sky130_fd_sc_hd__o2111ai_1 _08745_ (.A1(_02669_),
    .A2(_02678_),
    .B1(_02702_),
    .C1(_02703_),
    .D1(_02731_),
    .Y(_02733_));
 sky130_fd_sc_hd__o32a_1 _08746_ (.A1(_02661_),
    .A2(_02701_),
    .A3(_02733_),
    .B1(_02684_),
    .B2(_02621_),
    .X(_02734_));
 sky130_fd_sc_hd__a21bo_1 _08747_ (.A1(_02709_),
    .A2(_02714_),
    .B1_N(_02713_),
    .X(_02735_));
 sky130_fd_sc_hd__a22oi_1 _08748_ (.A1(_02441_),
    .A2(_02442_),
    .B1(_02443_),
    .B2(_02431_),
    .Y(_02736_));
 sky130_fd_sc_hd__nor2_1 _08749_ (.A(_02444_),
    .B(_02736_),
    .Y(_02738_));
 sky130_fd_sc_hd__nand2_1 _08750_ (.A(_02738_),
    .B(_02735_),
    .Y(_02739_));
 sky130_fd_sc_hd__xor2_1 _08751_ (.A(_02735_),
    .B(_02738_),
    .X(_02740_));
 sky130_fd_sc_hd__nand2_1 _08752_ (.A(_02707_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__xnor2_1 _08753_ (.A(_02707_),
    .B(_02740_),
    .Y(_02742_));
 sky130_fd_sc_hd__a21o_1 _08754_ (.A1(_02718_),
    .A2(_02720_),
    .B1(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__nand3_1 _08755_ (.A(_02718_),
    .B(_02720_),
    .C(_02742_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand2_1 _08756_ (.A(_02743_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__o32a_1 _08757_ (.A1(_02722_),
    .A2(_02723_),
    .A3(_02745_),
    .B1(_02728_),
    .B2(_02619_),
    .X(_02746_));
 sky130_fd_sc_hd__o21a_1 _08758_ (.A1(_02732_),
    .A2(_02734_),
    .B1(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__xnor2_1 _08759_ (.A(_02449_),
    .B(_02450_),
    .Y(_02749_));
 sky130_fd_sc_hd__a21o_1 _08760_ (.A1(_02739_),
    .A2(_02741_),
    .B1(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__nand3_1 _08761_ (.A(_02739_),
    .B(_02741_),
    .C(_02749_),
    .Y(_02751_));
 sky130_fd_sc_hd__nand2_1 _08762_ (.A(_02750_),
    .B(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__a22o_1 _08763_ (.A1(_02725_),
    .A2(_02745_),
    .B1(_02752_),
    .B2(_02743_),
    .X(_02753_));
 sky130_fd_sc_hd__o211ai_1 _08764_ (.A1(_02450_),
    .A2(_02449_),
    .B1(_02447_),
    .C1(_02453_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _08765_ (.A(_02454_),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__a211o_1 _08766_ (.A1(_02739_),
    .A2(_02741_),
    .B1(_02749_),
    .C1(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__o221a_1 _08767_ (.A1(_02743_),
    .A2(_02752_),
    .B1(_02753_),
    .B2(_02747_),
    .C1(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__a22o_1 _08768_ (.A1(_02454_),
    .A2(_02455_),
    .B1(_02750_),
    .B2(_02755_),
    .X(_02758_));
 sky130_fd_sc_hd__o21ai_1 _08769_ (.A1(_02758_),
    .A2(_02757_),
    .B1(_02456_),
    .Y(_02760_));
 sky130_fd_sc_hd__nand2_1 _08770_ (.A(_02392_),
    .B(_02320_),
    .Y(_02761_));
 sky130_fd_sc_hd__a32oi_4 _08771_ (.A1(_02391_),
    .A2(_02235_),
    .A3(_02239_),
    .B1(_02390_),
    .B2(_02321_),
    .Y(_02762_));
 sky130_fd_sc_hd__a31o_1 _08772_ (.A1(_02334_),
    .A2(_02347_),
    .A3(_02348_),
    .B1(_02351_),
    .X(_02763_));
 sky130_fd_sc_hd__o2bb2a_1 _08773_ (.A1_N(net41),
    .A2_N(net1),
    .B1(_01986_),
    .B2(_01987_),
    .X(_02764_));
 sky130_fd_sc_hd__a211oi_2 _08774_ (.A1(_02335_),
    .A2(_02337_),
    .B1(_02764_),
    .C1(_01990_),
    .Y(_02765_));
 sky130_fd_sc_hd__o211a_1 _08775_ (.A1(_01990_),
    .A2(_02764_),
    .B1(_02337_),
    .C1(_02335_),
    .X(_02766_));
 sky130_fd_sc_hd__o211ai_1 _08776_ (.A1(_02765_),
    .A2(_02766_),
    .B1(_02323_),
    .C1(_02325_),
    .Y(_02767_));
 sky130_fd_sc_hd__a211o_1 _08777_ (.A1(_02323_),
    .A2(_02325_),
    .B1(_02765_),
    .C1(_02766_),
    .X(_02768_));
 sky130_fd_sc_hd__and2_1 _08778_ (.A(_02767_),
    .B(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__a311o_1 _08779_ (.A1(_02334_),
    .A2(_02347_),
    .A3(_02348_),
    .B1(_02351_),
    .C1(_02769_),
    .X(_02771_));
 sky130_fd_sc_hd__nand2_1 _08780_ (.A(_02763_),
    .B(_02769_),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2_1 _08781_ (.A(_02771_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__xnor2_1 _08782_ (.A(_02327_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _08783_ (.A(_02345_),
    .B(_02347_),
    .Y(_02775_));
 sky130_fd_sc_hd__o2bb2a_1 _08784_ (.A1_N(_01981_),
    .A2_N(_01982_),
    .B1(_01087_),
    .B2(_01219_),
    .X(_02776_));
 sky130_fd_sc_hd__nor2_1 _08785_ (.A(_01983_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _08786_ (.A(_02340_),
    .B(_02343_),
    .Y(_02778_));
 sky130_fd_sc_hd__a22o_1 _08787_ (.A1(net35),
    .A2(net29),
    .B1(_01954_),
    .B2(_01955_),
    .X(_02779_));
 sky130_fd_sc_hd__and3_1 _08788_ (.A(_01957_),
    .B(_02778_),
    .C(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__nand3_1 _08789_ (.A(_01957_),
    .B(_02778_),
    .C(_02779_),
    .Y(_02782_));
 sky130_fd_sc_hd__a21oi_1 _08790_ (.A1(_01957_),
    .A2(_02779_),
    .B1(_02778_),
    .Y(_02783_));
 sky130_fd_sc_hd__a21o_1 _08791_ (.A1(_01957_),
    .A2(_02779_),
    .B1(_02778_),
    .X(_02784_));
 sky130_fd_sc_hd__and3_1 _08792_ (.A(_02784_),
    .B(_02777_),
    .C(_02782_),
    .X(_02785_));
 sky130_fd_sc_hd__a211o_1 _08793_ (.A1(_02782_),
    .A2(_02784_),
    .B1(_01983_),
    .C1(_02776_),
    .X(_02786_));
 sky130_fd_sc_hd__or3_1 _08794_ (.A(_02777_),
    .B(_02780_),
    .C(_02783_),
    .X(_02787_));
 sky130_fd_sc_hd__or4bb_1 _08795_ (.A(_02361_),
    .B(_02362_),
    .C_N(_02786_),
    .D_N(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__a2bb2o_1 _08796_ (.A1_N(_02361_),
    .A2_N(_02362_),
    .B1(_02786_),
    .B2(_02787_),
    .X(_02789_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_02788_),
    .B(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__xnor2_1 _08798_ (.A(_02775_),
    .B(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__inv_2 _08799_ (.A(_02791_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand2_1 _08800_ (.A(_02356_),
    .B(_02358_),
    .Y(_02794_));
 sky130_fd_sc_hd__nand2_1 _08801_ (.A(_02366_),
    .B(_02368_),
    .Y(_02795_));
 sky130_fd_sc_hd__a22o_1 _08802_ (.A1(net32),
    .A2(net63),
    .B1(_01937_),
    .B2(_01938_),
    .X(_02796_));
 sky130_fd_sc_hd__a21o_1 _08803_ (.A1(_01939_),
    .A2(_02796_),
    .B1(_02795_),
    .X(_02797_));
 sky130_fd_sc_hd__nand3_1 _08804_ (.A(_01939_),
    .B(_02795_),
    .C(_02796_),
    .Y(_02798_));
 sky130_fd_sc_hd__and3_1 _08805_ (.A(_02794_),
    .B(_02797_),
    .C(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__a21oi_1 _08806_ (.A1(_02797_),
    .A2(_02798_),
    .B1(_02794_),
    .Y(_02800_));
 sky130_fd_sc_hd__nor2_1 _08807_ (.A(_02799_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__nand2_1 _08808_ (.A(_02371_),
    .B(_02373_),
    .Y(_02802_));
 sky130_fd_sc_hd__a22o_1 _08809_ (.A1(_01928_),
    .A2(_01929_),
    .B1(_01931_),
    .B2(_01925_),
    .X(_02804_));
 sky130_fd_sc_hd__a21o_1 _08810_ (.A1(_01925_),
    .A2(_01931_),
    .B1(_01930_),
    .X(_02805_));
 sky130_fd_sc_hd__nand3_1 _08811_ (.A(_01925_),
    .B(_01930_),
    .C(_01931_),
    .Y(_02806_));
 sky130_fd_sc_hd__nand3_2 _08812_ (.A(_01932_),
    .B(_02802_),
    .C(_02804_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand4_1 _08813_ (.A(_02371_),
    .B(_02373_),
    .C(_02805_),
    .D(_02806_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _08814_ (.A(_02807_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__or3_1 _08815_ (.A(_02799_),
    .B(_02800_),
    .C(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__a211o_1 _08816_ (.A1(_02807_),
    .A2(_02808_),
    .B1(_02799_),
    .C1(_02800_),
    .X(_02811_));
 sky130_fd_sc_hd__or2_1 _08817_ (.A(_02801_),
    .B(_02809_),
    .X(_02812_));
 sky130_fd_sc_hd__a22oi_1 _08818_ (.A1(_02377_),
    .A2(_02379_),
    .B1(_02811_),
    .B2(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__a22o_1 _08819_ (.A1(_02377_),
    .A2(_02379_),
    .B1(_02811_),
    .B2(_02812_),
    .X(_02815_));
 sky130_fd_sc_hd__and4_1 _08820_ (.A(_02377_),
    .B(_02379_),
    .C(_02811_),
    .D(_02812_),
    .X(_02816_));
 sky130_fd_sc_hd__nor2_1 _08821_ (.A(_02813_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__or3_1 _08822_ (.A(_02813_),
    .B(_02816_),
    .C(_02793_),
    .X(_02818_));
 sky130_fd_sc_hd__xnor2_1 _08823_ (.A(_02791_),
    .B(_02817_),
    .Y(_02819_));
 sky130_fd_sc_hd__a21o_1 _08824_ (.A1(_02381_),
    .A2(_02383_),
    .B1(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__nand3_1 _08825_ (.A(_02381_),
    .B(_02383_),
    .C(_02819_),
    .Y(_02821_));
 sky130_fd_sc_hd__and2_1 _08826_ (.A(_02820_),
    .B(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__nand2_1 _08827_ (.A(_02774_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__or2_1 _08828_ (.A(_02774_),
    .B(_02822_),
    .X(_02824_));
 sky130_fd_sc_hd__nand2_1 _08829_ (.A(_02823_),
    .B(_02824_),
    .Y(_02826_));
 sky130_fd_sc_hd__a21oi_1 _08830_ (.A1(_02386_),
    .A2(_02388_),
    .B1(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__and3_1 _08831_ (.A(_02386_),
    .B(_02388_),
    .C(_02826_),
    .X(_02828_));
 sky130_fd_sc_hd__nor2_1 _08832_ (.A(_02827_),
    .B(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__xnor2_1 _08833_ (.A(_02331_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand2_1 _08834_ (.A(_02830_),
    .B(_02762_),
    .Y(_02831_));
 sky130_fd_sc_hd__and3_1 _08835_ (.A(_02760_),
    .B(_02761_),
    .C(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__a21oi_1 _08836_ (.A1(_02331_),
    .A2(_02829_),
    .B1(_02827_),
    .Y(_02833_));
 sky130_fd_sc_hd__a21boi_1 _08837_ (.A1(_02771_),
    .A2(_02327_),
    .B1_N(_02772_),
    .Y(_02834_));
 sky130_fd_sc_hd__or3_1 _08838_ (.A(_02325_),
    .B(_02765_),
    .C(_02766_),
    .X(_02835_));
 sky130_fd_sc_hd__a21bo_1 _08839_ (.A1(_02775_),
    .A2(_02788_),
    .B1_N(_02789_),
    .X(_02837_));
 sky130_fd_sc_hd__a21o_1 _08840_ (.A1(_01985_),
    .A2(_01992_),
    .B1(_01991_),
    .X(_02838_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(_01993_),
    .B(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__o21bai_1 _08842_ (.A1(_02323_),
    .A2(_02766_),
    .B1_N(_02765_),
    .Y(_02840_));
 sky130_fd_sc_hd__nand3_1 _08843_ (.A(_02840_),
    .B(_02838_),
    .C(_01993_),
    .Y(_02841_));
 sky130_fd_sc_hd__xor2_1 _08844_ (.A(_02839_),
    .B(_02840_),
    .X(_02842_));
 sky130_fd_sc_hd__xor2_1 _08845_ (.A(_01873_),
    .B(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__nor2_1 _08846_ (.A(_02837_),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__nand2_1 _08847_ (.A(_02843_),
    .B(_02837_),
    .Y(_02845_));
 sky130_fd_sc_hd__and2b_1 _08848_ (.A_N(_02844_),
    .B(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__xnor2_1 _08849_ (.A(_02835_),
    .B(_02846_),
    .Y(_02848_));
 sky130_fd_sc_hd__a31o_1 _08850_ (.A1(_01939_),
    .A2(_02795_),
    .A3(_02796_),
    .B1(_02799_),
    .X(_02849_));
 sky130_fd_sc_hd__a2bb2o_1 _08851_ (.A1_N(_01858_),
    .A2_N(_01962_),
    .B1(_01964_),
    .B2(_01961_),
    .X(_02850_));
 sky130_fd_sc_hd__a21o_1 _08852_ (.A1(_01966_),
    .A2(_02850_),
    .B1(_02849_),
    .X(_02851_));
 sky130_fd_sc_hd__nand3_2 _08853_ (.A(_01966_),
    .B(_02849_),
    .C(_02850_),
    .Y(_02852_));
 sky130_fd_sc_hd__o211ai_2 _08854_ (.A1(_02780_),
    .A2(_02785_),
    .B1(_02851_),
    .C1(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__a221o_1 _08855_ (.A1(_02777_),
    .A2(_02784_),
    .B1(_02851_),
    .B2(_02852_),
    .C1(_02780_),
    .X(_02854_));
 sky130_fd_sc_hd__and2_1 _08856_ (.A(_02853_),
    .B(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__nand2_1 _08857_ (.A(_01950_),
    .B(_01948_),
    .Y(_02856_));
 sky130_fd_sc_hd__a21o_1 _08858_ (.A1(_01946_),
    .A2(_01947_),
    .B1(_01950_),
    .X(_02857_));
 sky130_fd_sc_hd__a22oi_2 _08859_ (.A1(_02807_),
    .A2(_02810_),
    .B1(_02856_),
    .B2(_02857_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand4_1 _08860_ (.A(_02807_),
    .B(_02810_),
    .C(_02856_),
    .D(_02857_),
    .Y(_02860_));
 sky130_fd_sc_hd__and2b_1 _08861_ (.A_N(_02859_),
    .B(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__xnor2_1 _08862_ (.A(_02855_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__a21o_1 _08863_ (.A1(_02815_),
    .A2(_02818_),
    .B1(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__o211ai_1 _08864_ (.A1(_02816_),
    .A2(_02793_),
    .B1(_02815_),
    .C1(_02862_),
    .Y(_02864_));
 sky130_fd_sc_hd__and2_1 _08865_ (.A(_02863_),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_02848_),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__or2_1 _08867_ (.A(_02848_),
    .B(_02865_),
    .X(_02867_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(_02866_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__a21o_1 _08869_ (.A1(_02820_),
    .A2(_02823_),
    .B1(_02868_),
    .X(_02870_));
 sky130_fd_sc_hd__nand3_1 _08870_ (.A(_02820_),
    .B(_02823_),
    .C(_02868_),
    .Y(_02871_));
 sky130_fd_sc_hd__and2_1 _08871_ (.A(_02870_),
    .B(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__nand2b_1 _08872_ (.A_N(_02834_),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__nand2b_1 _08873_ (.A_N(_02872_),
    .B(_02834_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(_02873_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__o22ai_1 _08875_ (.A1(_02762_),
    .A2(_02830_),
    .B1(_02833_),
    .B2(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__o21ai_1 _08876_ (.A1(_01873_),
    .A2(_02842_),
    .B1(_02841_),
    .Y(_02877_));
 sky130_fd_sc_hd__o21a_1 _08877_ (.A1(_01874_),
    .A2(_01997_),
    .B1(_01999_),
    .X(_02878_));
 sky130_fd_sc_hd__o211a_1 _08878_ (.A1(_02001_),
    .A2(_02878_),
    .B1(_02853_),
    .C1(_02852_),
    .X(_02879_));
 sky130_fd_sc_hd__a211oi_2 _08879_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_02878_),
    .C1(_02001_),
    .Y(_02881_));
 sky130_fd_sc_hd__nor2_1 _08880_ (.A(_02879_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__xor2_1 _08881_ (.A(_02877_),
    .B(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__a31o_1 _08882_ (.A1(_02853_),
    .A2(_02854_),
    .A3(_02860_),
    .B1(_02859_),
    .X(_02884_));
 sky130_fd_sc_hd__a22o_1 _08883_ (.A1(_01972_),
    .A2(_01973_),
    .B1(_01974_),
    .B2(_01953_),
    .X(_02885_));
 sky130_fd_sc_hd__nand3_1 _08884_ (.A(_01975_),
    .B(_02884_),
    .C(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__a221o_1 _08885_ (.A1(_02855_),
    .A2(_02860_),
    .B1(_02885_),
    .B2(_01975_),
    .C1(_02859_),
    .X(_02887_));
 sky130_fd_sc_hd__and2_1 _08886_ (.A(_02886_),
    .B(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__nand2_1 _08887_ (.A(_02883_),
    .B(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__or2_1 _08888_ (.A(_02883_),
    .B(_02888_),
    .X(_02890_));
 sky130_fd_sc_hd__nand2_1 _08889_ (.A(_02889_),
    .B(_02890_),
    .Y(_02892_));
 sky130_fd_sc_hd__a21oi_1 _08890_ (.A1(_02863_),
    .A2(_02866_),
    .B1(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__o21ai_1 _08891_ (.A1(_02835_),
    .A2(_02844_),
    .B1(_02845_),
    .Y(_02894_));
 sky130_fd_sc_hd__and3_1 _08892_ (.A(_02863_),
    .B(_02866_),
    .C(_02892_),
    .X(_02895_));
 sky130_fd_sc_hd__nor2_1 _08893_ (.A(_02893_),
    .B(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__a21o_1 _08894_ (.A1(_02896_),
    .A2(_02894_),
    .B1(_02893_),
    .X(_02897_));
 sky130_fd_sc_hd__a21oi_1 _08895_ (.A1(_02882_),
    .A2(_02877_),
    .B1(_02881_),
    .Y(_02898_));
 sky130_fd_sc_hd__a21o_1 _08896_ (.A1(_01979_),
    .A2(_02009_),
    .B1(_02008_),
    .X(_02899_));
 sky130_fd_sc_hd__nand2_1 _08897_ (.A(_02010_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__a21oi_1 _08898_ (.A1(_02886_),
    .A2(_02889_),
    .B1(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__and3_1 _08899_ (.A(_02886_),
    .B(_02889_),
    .C(_02900_),
    .X(_02903_));
 sky130_fd_sc_hd__nor2_1 _08900_ (.A(_02901_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__and2b_1 _08901_ (.A_N(_02898_),
    .B(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__a211oi_1 _08902_ (.A1(_02882_),
    .A2(_02877_),
    .B1(_02881_),
    .C1(_02904_),
    .Y(_02906_));
 sky130_fd_sc_hd__or2_1 _08903_ (.A(_02905_),
    .B(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__nand2b_1 _08904_ (.A_N(_02907_),
    .B(_02897_),
    .Y(_02908_));
 sky130_fd_sc_hd__xnor2_1 _08905_ (.A(_02897_),
    .B(_02907_),
    .Y(_02909_));
 sky130_fd_sc_hd__xnor2_1 _08906_ (.A(_02894_),
    .B(_02896_),
    .Y(_02910_));
 sky130_fd_sc_hd__a21oi_1 _08907_ (.A1(_02870_),
    .A2(_02873_),
    .B1(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__and3_1 _08908_ (.A(_02870_),
    .B(_02873_),
    .C(_02910_),
    .X(_02912_));
 sky130_fd_sc_hd__nor2_1 _08909_ (.A(_02911_),
    .B(_02912_),
    .Y(_02914_));
 sky130_fd_sc_hd__nand2_1 _08910_ (.A(_02875_),
    .B(_02833_),
    .Y(_02915_));
 sky130_fd_sc_hd__o2111ai_2 _08911_ (.A1(_02832_),
    .A2(_02876_),
    .B1(_02909_),
    .C1(_02915_),
    .D1(_02914_),
    .Y(_02916_));
 sky130_fd_sc_hd__nand2_1 _08912_ (.A(_02016_),
    .B(_02018_),
    .Y(_02917_));
 sky130_fd_sc_hd__nand2_1 _08913_ (.A(_02019_),
    .B(_02917_),
    .Y(_02918_));
 sky130_fd_sc_hd__o21bai_2 _08914_ (.A1(_02901_),
    .A2(_02905_),
    .B1_N(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__or3b_1 _08915_ (.A(_02901_),
    .B(_02905_),
    .C_N(_02918_),
    .X(_02920_));
 sky130_fd_sc_hd__nand2_1 _08916_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__nand2_1 _08917_ (.A(_02909_),
    .B(_02911_),
    .Y(_02922_));
 sky130_fd_sc_hd__o211a_1 _08918_ (.A1(_02908_),
    .A2(_02921_),
    .B1(_02922_),
    .C1(_02916_),
    .X(_02923_));
 sky130_fd_sc_hd__xnor2_2 _08919_ (.A(_02015_),
    .B(_02025_),
    .Y(_02925_));
 sky130_fd_sc_hd__a22o_1 _08920_ (.A1(_02908_),
    .A2(_02921_),
    .B1(_02925_),
    .B2(_02919_),
    .X(_02926_));
 sky130_fd_sc_hd__o22ai_4 _08921_ (.A1(_02919_),
    .A2(_02925_),
    .B1(_02926_),
    .B2(_02923_),
    .Y(_02927_));
 sky130_fd_sc_hd__o21ba_1 _08922_ (.A1(_02028_),
    .A2(_02927_),
    .B1_N(_02029_),
    .X(_02928_));
 sky130_fd_sc_hd__nand2_1 _08923_ (.A(_02928_),
    .B(_01914_),
    .Y(_02929_));
 sky130_fd_sc_hd__a211oi_1 _08924_ (.A1(_01913_),
    .A2(_02929_),
    .B1(_01788_),
    .C1(_01789_),
    .Y(_02930_));
 sky130_fd_sc_hd__o21ai_1 _08925_ (.A1(_01788_),
    .A2(_02930_),
    .B1(_01667_),
    .Y(_02931_));
 sky130_fd_sc_hd__and2b_1 _08926_ (.A_N(_01540_),
    .B(_01541_),
    .X(_02932_));
 sky130_fd_sc_hd__or2_1 _08927_ (.A(_01542_),
    .B(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__a21oi_1 _08928_ (.A1(_01665_),
    .A2(_02931_),
    .B1(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__nor2_1 _08929_ (.A(_01542_),
    .B(_02934_),
    .Y(_02936_));
 sky130_fd_sc_hd__nor2_1 _08930_ (.A(_01419_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__o21a_1 _08931_ (.A1(_01418_),
    .A2(_02937_),
    .B1(_01293_),
    .X(_02938_));
 sky130_fd_sc_hd__o21a_1 _08932_ (.A1(_01291_),
    .A2(_02938_),
    .B1(_01156_),
    .X(_02939_));
 sky130_fd_sc_hd__o21a_1 _08933_ (.A1(_01154_),
    .A2(_02939_),
    .B1(_01023_),
    .X(_02940_));
 sky130_fd_sc_hd__o21a_1 _08934_ (.A1(_01022_),
    .A2(_02940_),
    .B1(_00903_),
    .X(_02941_));
 sky130_fd_sc_hd__xor2_1 _08935_ (.A(_00792_),
    .B(_00794_),
    .X(_02942_));
 sky130_fd_sc_hd__o21a_1 _08936_ (.A1(_00901_),
    .A2(_02941_),
    .B1(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__a21oi_1 _08937_ (.A1(_00792_),
    .A2(_00794_),
    .B1(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__o21ai_1 _08938_ (.A1(_00692_),
    .A2(_02944_),
    .B1(_00690_),
    .Y(_02945_));
 sky130_fd_sc_hd__nand2_1 _08939_ (.A(_02945_),
    .B(_00601_),
    .Y(_02947_));
 sky130_fd_sc_hd__a21oi_1 _08940_ (.A1(_00599_),
    .A2(_02947_),
    .B1(_00509_),
    .Y(_02948_));
 sky130_fd_sc_hd__a21oi_1 _08941_ (.A1(_00506_),
    .A2(_00508_),
    .B1(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__nor2_1 _08942_ (.A(_00424_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__a21oi_1 _08943_ (.A1(_00422_),
    .A2(_00423_),
    .B1(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__a211oi_1 _08944_ (.A1(_00337_),
    .A2(_00335_),
    .B1(_00334_),
    .C1(_00340_),
    .Y(_02952_));
 sky130_fd_sc_hd__or2_1 _08945_ (.A(_00341_),
    .B(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__o21bai_1 _08946_ (.A1(_02953_),
    .A2(_02951_),
    .B1_N(_00341_),
    .Y(_02954_));
 sky130_fd_sc_hd__nand2b_1 _08947_ (.A_N(_00263_),
    .B(_00264_),
    .Y(_02955_));
 sky130_fd_sc_hd__a21oi_1 _08948_ (.A1(_00264_),
    .A2(_02954_),
    .B1(_00263_),
    .Y(_02956_));
 sky130_fd_sc_hd__or2_1 _08949_ (.A(_00197_),
    .B(_02956_),
    .X(_02958_));
 sky130_fd_sc_hd__a21oi_1 _08950_ (.A1(_00195_),
    .A2(_02958_),
    .B1(_00136_),
    .Y(_02959_));
 sky130_fd_sc_hd__o21a_1 _08951_ (.A1(_00134_),
    .A2(_02959_),
    .B1(_00083_),
    .X(_02960_));
 sky130_fd_sc_hd__o21ai_1 _08952_ (.A1(_00081_),
    .A2(_02960_),
    .B1(_05392_),
    .Y(_02961_));
 sky130_fd_sc_hd__inv_2 _08953_ (.A(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__a31o_1 _08954_ (.A1(_05344_),
    .A2(_05388_),
    .A3(_05390_),
    .B1(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__a21o_2 _08955_ (.A1(_02963_),
    .A2(_05349_),
    .B1(_05346_),
    .X(_02964_));
 sky130_fd_sc_hd__nor2_1 _08956_ (.A(_05304_),
    .B(_05298_),
    .Y(_02965_));
 sky130_fd_sc_hd__or2_1 _08957_ (.A(_05305_),
    .B(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__inv_2 _08958_ (.A(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__nand2_1 _08959_ (.A(_02964_),
    .B(_02967_),
    .Y(_02969_));
 sky130_fd_sc_hd__a21oi_4 _08960_ (.A1(_02964_),
    .A2(_02967_),
    .B1(_05305_),
    .Y(_02970_));
 sky130_fd_sc_hd__a21o_4 _08961_ (.A1(_02964_),
    .A2(_02967_),
    .B1(_05305_),
    .X(_02971_));
 sky130_fd_sc_hd__a31o_4 _08962_ (.A1(net46),
    .A2(net14),
    .A3(_05227_),
    .B1(_05226_),
    .X(_02972_));
 sky130_fd_sc_hd__a21boi_4 _08963_ (.A1(_05284_),
    .A2(_05291_),
    .B1_N(_05300_),
    .Y(_02973_));
 sky130_fd_sc_hd__nor2_2 _08964_ (.A(_02972_),
    .B(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__a2bb2o_1 _08965_ (.A1_N(_02972_),
    .A2_N(_02973_),
    .B1(_02967_),
    .B2(_02964_),
    .X(_02975_));
 sky130_fd_sc_hd__and3b_4 _08966_ (.A_N(_05305_),
    .B(_02969_),
    .C(_02974_),
    .X(_02976_));
 sky130_fd_sc_hd__or3_4 _08967_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .X(_02977_));
 sky130_fd_sc_hd__nor3_1 _08968_ (.A(_02028_),
    .B(_02029_),
    .C(_02927_),
    .Y(_02978_));
 sky130_fd_sc_hd__o21ai_1 _08969_ (.A1(_02028_),
    .A2(_02029_),
    .B1(_02927_),
    .Y(_02980_));
 sky130_fd_sc_hd__or3b_1 _08970_ (.A(_02977_),
    .B(_02978_),
    .C_N(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__xor2_1 _08971_ (.A(_01914_),
    .B(_02928_),
    .X(_02982_));
 sky130_fd_sc_hd__a21o_1 _08972_ (.A1(_02970_),
    .A2(_02974_),
    .B1(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__nor4_1 _08973_ (.A(net19),
    .B(net18),
    .C(net17),
    .D(net16),
    .Y(_02984_));
 sky130_fd_sc_hd__nor3_1 _08974_ (.A(net24),
    .B(net22),
    .C(net21),
    .Y(_02985_));
 sky130_fd_sc_hd__or4_1 _08975_ (.A(net51),
    .B(net50),
    .C(net49),
    .D(net48),
    .X(_02986_));
 sky130_fd_sc_hd__or4_1 _08976_ (.A(net56),
    .B(net54),
    .C(net53),
    .D(net52),
    .X(_02987_));
 sky130_fd_sc_hd__nor2_1 _08977_ (.A(_02986_),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__a311o_4 _08978_ (.A1(_00977_),
    .A2(_02984_),
    .A3(_02985_),
    .B1(_02988_),
    .C1(net65),
    .X(_02989_));
 sky130_fd_sc_hd__and4_1 _08979_ (.A(net51),
    .B(net50),
    .C(net49),
    .D(net48),
    .X(_02991_));
 sky130_fd_sc_hd__and3_1 _08980_ (.A(net56),
    .B(net54),
    .C(net53),
    .X(_02992_));
 sky130_fd_sc_hd__and3_1 _08981_ (.A(net52),
    .B(_02991_),
    .C(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__and4_1 _08982_ (.A(net19),
    .B(net18),
    .C(net17),
    .D(net16),
    .X(_02994_));
 sky130_fd_sc_hd__and3_1 _08983_ (.A(net24),
    .B(net22),
    .C(net21),
    .X(_02995_));
 sky130_fd_sc_hd__a31o_4 _08984_ (.A1(net20),
    .A2(_02994_),
    .A3(_02995_),
    .B1(_02993_),
    .X(_02996_));
 sky130_fd_sc_hd__nor2_8 _08985_ (.A(_02989_),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__nand3_1 _08986_ (.A(_05004_),
    .B(_05005_),
    .C(\adder_inst.fraction1_32neg[0] ),
    .Y(_02998_));
 sky130_fd_sc_hd__xor2_1 _08987_ (.A(\adder_inst.fraction1_32neg[0] ),
    .B(\adder_inst.fraction2[0] ),
    .X(_02999_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(\adder_inst.fraction1[0] ),
    .B(\adder_inst.fraction2[0] ),
    .Y(_03000_));
 sky130_fd_sc_hd__a21o_1 _08989_ (.A1(_05004_),
    .A2(_05005_),
    .B1(\adder_inst.fraction1[0] ),
    .X(_03002_));
 sky130_fd_sc_hd__and2_1 _08990_ (.A(_03000_),
    .B(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__a221o_1 _08991_ (.A1(_01263_),
    .A2(_02088_),
    .B1(_05002_),
    .B2(_03847_),
    .C1(_01274_),
    .X(_03004_));
 sky130_fd_sc_hd__nand2_1 _08992_ (.A(_01274_),
    .B(_05003_),
    .Y(_03005_));
 sky130_fd_sc_hd__a211o_1 _08993_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_05230_),
    .C1(_05232_),
    .X(_03006_));
 sky130_fd_sc_hd__o221a_2 _08994_ (.A1(_00000_),
    .A2(_02999_),
    .B1(_03003_),
    .B2(_05233_),
    .C1(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__nand2_1 _08995_ (.A(_04623_),
    .B(_04634_),
    .Y(_03008_));
 sky130_fd_sc_hd__o21ai_1 _08996_ (.A1(_05008_),
    .A2(_05029_),
    .B1(_05034_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand2_1 _08997_ (.A(_04975_),
    .B(\adder_inst.fraction2[0] ),
    .Y(_03010_));
 sky130_fd_sc_hd__and3_1 _08998_ (.A(_04975_),
    .B(\adder_inst.fraction1[0] ),
    .C(\adder_inst.fraction2[0] ),
    .X(_03011_));
 sky130_fd_sc_hd__a21oi_1 _08999_ (.A1(\adder_inst.fraction1[0] ),
    .A2(\adder_inst.fraction2[0] ),
    .B1(_04975_),
    .Y(_03013_));
 sky130_fd_sc_hd__xnor2_1 _09000_ (.A(_04979_),
    .B(\adder_inst.fraction1[0] ),
    .Y(_00034_));
 sky130_fd_sc_hd__a211oi_1 _09001_ (.A1(_04936_),
    .A2(_04943_),
    .B1(_03011_),
    .C1(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__o22ai_2 _09002_ (.A1(_05003_),
    .A2(_03010_),
    .B1(_04956_),
    .B2(_03013_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand2_1 _09003_ (.A(_05031_),
    .B(_05033_),
    .Y(_03016_));
 sky130_fd_sc_hd__a21boi_2 _09004_ (.A1(_03015_),
    .A2(_03016_),
    .B1_N(_03009_),
    .Y(_03017_));
 sky130_fd_sc_hd__nand2_1 _09005_ (.A(_04612_),
    .B(_04645_),
    .Y(_03018_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(_03009_),
    .B(_03016_),
    .Y(_03019_));
 sky130_fd_sc_hd__xor2_1 _09007_ (.A(_04949_),
    .B(_04979_),
    .X(_03020_));
 sky130_fd_sc_hd__nand4_1 _09008_ (.A(_03000_),
    .B(_03002_),
    .C(_03009_),
    .D(_03016_),
    .Y(_03021_));
 sky130_fd_sc_hd__o21ai_1 _09009_ (.A1(_03021_),
    .A2(_03020_),
    .B1(_03018_),
    .Y(_03023_));
 sky130_fd_sc_hd__and2_1 _09010_ (.A(_03008_),
    .B(_03018_),
    .X(_03024_));
 sky130_fd_sc_hd__a2bb2o_1 _09011_ (.A1_N(_03017_),
    .A2_N(_03023_),
    .B1(_04623_),
    .B2(_04634_),
    .X(_03025_));
 sky130_fd_sc_hd__a221o_1 _09012_ (.A1(net27),
    .A2(_02088_),
    .B1(_03902_),
    .B2(_04295_),
    .C1(_04339_),
    .X(_03026_));
 sky130_fd_sc_hd__nand2_1 _09013_ (.A(_04317_),
    .B(_04339_),
    .Y(_03027_));
 sky130_fd_sc_hd__nand2_1 _09014_ (.A(_03026_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_05049_),
    .B(_05051_),
    .Y(_03029_));
 sky130_fd_sc_hd__o211ai_2 _09016_ (.A1(_03017_),
    .A2(_03023_),
    .B1(_03027_),
    .C1(_03008_),
    .Y(_03030_));
 sky130_fd_sc_hd__o211ai_2 _09017_ (.A1(_04317_),
    .A2(_04339_),
    .B1(_03880_),
    .C1(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__a2bb2oi_1 _09018_ (.A1_N(_03836_),
    .A2_N(_03869_),
    .B1(_03026_),
    .B2(_03030_),
    .Y(_03032_));
 sky130_fd_sc_hd__a2bb2o_1 _09019_ (.A1_N(_03836_),
    .A2_N(_03869_),
    .B1(_03026_),
    .B2(_03030_),
    .X(_03034_));
 sky130_fd_sc_hd__nand2_1 _09020_ (.A(_03031_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__o21ai_2 _09021_ (.A1(_03825_),
    .A2(_03032_),
    .B1(_03031_),
    .Y(_03036_));
 sky130_fd_sc_hd__o21ai_2 _09022_ (.A1(_05049_),
    .A2(_05051_),
    .B1(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__a2bb2oi_2 _09023_ (.A1_N(_05064_),
    .A2_N(_05065_),
    .B1(_03029_),
    .B2(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__nand3_1 _09024_ (.A(_03037_),
    .B(_05068_),
    .C(_03029_),
    .Y(_03039_));
 sky130_fd_sc_hd__a31oi_2 _09025_ (.A1(_03037_),
    .A2(_05068_),
    .A3(_03029_),
    .B1(_05063_),
    .Y(_03040_));
 sky130_fd_sc_hd__and4_1 _09026_ (.A(_05083_),
    .B(_05094_),
    .C(_05103_),
    .D(_05113_),
    .X(_03041_));
 sky130_fd_sc_hd__o21ai_1 _09027_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__o22ai_2 _09028_ (.A1(_05097_),
    .A2(_05099_),
    .B1(_03038_),
    .B2(_03040_),
    .Y(_03043_));
 sky130_fd_sc_hd__a22oi_2 _09029_ (.A1(_05106_),
    .A2(_05107_),
    .B1(_03043_),
    .B2(_05101_),
    .Y(_03045_));
 sky130_fd_sc_hd__o211ai_2 _09030_ (.A1(_05098_),
    .A2(_05100_),
    .B1(_05110_),
    .C1(_03043_),
    .Y(_03046_));
 sky130_fd_sc_hd__and2b_1 _09031_ (.A_N(_03045_),
    .B(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__a21oi_2 _09032_ (.A1(_05111_),
    .A2(_03046_),
    .B1(_03045_),
    .Y(_03048_));
 sky130_fd_sc_hd__o21a_1 _09033_ (.A1(_05081_),
    .A2(_03048_),
    .B1(_05082_),
    .X(_03049_));
 sky130_fd_sc_hd__o211ai_1 _09034_ (.A1(_05081_),
    .A2(_03048_),
    .B1(_05093_),
    .C1(_05082_),
    .Y(_03050_));
 sky130_fd_sc_hd__a21oi_1 _09035_ (.A1(_05088_),
    .A2(_05092_),
    .B1(_03041_),
    .Y(_03051_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(_03050_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__a21boi_1 _09037_ (.A1(_03050_),
    .A2(_03051_),
    .B1_N(_03042_),
    .Y(_03053_));
 sky130_fd_sc_hd__o2bb2ai_1 _09038_ (.A1_N(_03042_),
    .A2_N(_03052_),
    .B1(_05124_),
    .B2(_05125_),
    .Y(_03054_));
 sky130_fd_sc_hd__a22oi_1 _09039_ (.A1(_05150_),
    .A2(_05151_),
    .B1(_03054_),
    .B2(_05128_),
    .Y(_03056_));
 sky130_fd_sc_hd__a221o_1 _09040_ (.A1(_01098_),
    .A2(_02088_),
    .B1(_05128_),
    .B2(_03054_),
    .C1(_05152_),
    .X(_03057_));
 sky130_fd_sc_hd__o211ai_2 _09041_ (.A1(_05127_),
    .A2(_03053_),
    .B1(_05154_),
    .C1(_05128_),
    .Y(_03058_));
 sky130_fd_sc_hd__and3_1 _09042_ (.A(_03057_),
    .B(_03058_),
    .C(_05148_),
    .X(_03059_));
 sky130_fd_sc_hd__a21oi_1 _09043_ (.A1(_05148_),
    .A2(_03058_),
    .B1(_03056_),
    .Y(_03060_));
 sky130_fd_sc_hd__o21bai_1 _09044_ (.A1(_05136_),
    .A2(_03060_),
    .B1_N(_05137_),
    .Y(_03061_));
 sky130_fd_sc_hd__or4bb_1 _09045_ (.A(_05136_),
    .B(_05137_),
    .C_N(_05156_),
    .D_N(_05129_),
    .X(_03062_));
 sky130_fd_sc_hd__o21a_1 _09046_ (.A1(_05140_),
    .A2(_05143_),
    .B1(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__nand2_1 _09047_ (.A(_03061_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__a2bb2o_1 _09048_ (.A1_N(_03062_),
    .A2_N(_03053_),
    .B1(_05143_),
    .B2(_05140_),
    .X(_03065_));
 sky130_fd_sc_hd__o21ai_1 _09049_ (.A1(_05140_),
    .A2(_05143_),
    .B1(_03065_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _09050_ (.A(_03064_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__inv_2 _09051_ (.A(_03068_),
    .Y(_03069_));
 sky130_fd_sc_hd__or4b_2 _09052_ (.A(_05169_),
    .B(_05175_),
    .C(_05190_),
    .D_N(_05183_),
    .X(_03070_));
 sky130_fd_sc_hd__nand3_1 _09053_ (.A(_05188_),
    .B(_03064_),
    .C(_03067_),
    .Y(_03071_));
 sky130_fd_sc_hd__o21ai_1 _09054_ (.A1(_05185_),
    .A2(_05187_),
    .B1(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__o211ai_1 _09055_ (.A1(_05185_),
    .A2(_05187_),
    .B1(_03071_),
    .C1(_05179_),
    .Y(_03073_));
 sky130_fd_sc_hd__a21oi_1 _09056_ (.A1(_05189_),
    .A2(_03071_),
    .B1(_05179_),
    .Y(_03074_));
 sky130_fd_sc_hd__xor2_1 _09057_ (.A(_05178_),
    .B(_03072_),
    .X(_03075_));
 sky130_fd_sc_hd__o21ai_2 _09058_ (.A1(_05181_),
    .A2(_03074_),
    .B1(_03073_),
    .Y(_03076_));
 sky130_fd_sc_hd__a21o_1 _09059_ (.A1(_05166_),
    .A2(_03076_),
    .B1(_05168_),
    .X(_03078_));
 sky130_fd_sc_hd__a221oi_2 _09060_ (.A1(_05171_),
    .A2(_05174_),
    .B1(_03076_),
    .B2(_05166_),
    .C1(_05168_),
    .Y(_03079_));
 sky130_fd_sc_hd__o21ai_1 _09061_ (.A1(_05171_),
    .A2(_05174_),
    .B1(_03070_),
    .Y(_03080_));
 sky130_fd_sc_hd__o22ai_4 _09062_ (.A1(_03069_),
    .A2(_03070_),
    .B1(_03080_),
    .B2(_03079_),
    .Y(_03081_));
 sky130_fd_sc_hd__o21bai_4 _09063_ (.A1(_05221_),
    .A2(_03081_),
    .B1_N(_05220_),
    .Y(_03082_));
 sky130_fd_sc_hd__nor2_2 _09064_ (.A(_05206_),
    .B(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__nand2_1 _09065_ (.A(_03082_),
    .B(_05206_),
    .Y(_03084_));
 sky130_fd_sc_hd__a21o_1 _09066_ (.A1(_03082_),
    .A2(_05206_),
    .B1(net114),
    .X(_03085_));
 sky130_fd_sc_hd__nand2b_4 _09067_ (.A_N(_03083_),
    .B(_03084_),
    .Y(_03086_));
 sky130_fd_sc_hd__a211o_4 _09068_ (.A1(_05206_),
    .A2(_03082_),
    .B1(net114),
    .C1(_03083_),
    .X(_03087_));
 sky130_fd_sc_hd__and2_1 _09069_ (.A(_05163_),
    .B(\adder_inst.fraction1_32neg[18] ),
    .X(_03089_));
 sky130_fd_sc_hd__nand2_1 _09070_ (.A(_05163_),
    .B(\adder_inst.fraction1_32neg[18] ),
    .Y(_03090_));
 sky130_fd_sc_hd__nor2_2 _09071_ (.A(\adder_inst.fraction1_32neg[18] ),
    .B(_05163_),
    .Y(_03091_));
 sky130_fd_sc_hd__nor2_1 _09072_ (.A(\adder_inst.fraction1_32neg[16] ),
    .B(_05187_),
    .Y(_03092_));
 sky130_fd_sc_hd__or2_1 _09073_ (.A(\adder_inst.fraction1_32neg[16] ),
    .B(_05187_),
    .X(_03093_));
 sky130_fd_sc_hd__nand2_1 _09074_ (.A(_01296_),
    .B(_04612_),
    .Y(_03094_));
 sky130_fd_sc_hd__and2_1 _09075_ (.A(_05034_),
    .B(\adder_inst.fraction1_32neg[2] ),
    .X(_03095_));
 sky130_fd_sc_hd__nand2_1 _09076_ (.A(_05034_),
    .B(\adder_inst.fraction1_32neg[2] ),
    .Y(_03096_));
 sky130_fd_sc_hd__and4_1 _09077_ (.A(_05004_),
    .B(_05005_),
    .C(\adder_inst.fraction1_32neg[0] ),
    .D(\adder_inst.fraction1_32neg[1] ),
    .X(_03097_));
 sky130_fd_sc_hd__a21oi_1 _09078_ (.A1(\adder_inst.fraction1_32neg[0] ),
    .A2(\adder_inst.fraction2[0] ),
    .B1(\adder_inst.fraction1_32neg[1] ),
    .Y(_03098_));
 sky130_fd_sc_hd__nor2_1 _09079_ (.A(_03097_),
    .B(_03098_),
    .Y(_03100_));
 sky130_fd_sc_hd__a22oi_2 _09080_ (.A1(_04936_),
    .A2(_04943_),
    .B1(_02998_),
    .B2(_01285_),
    .Y(_03101_));
 sky130_fd_sc_hd__a221o_1 _09081_ (.A1(net55),
    .A2(_02077_),
    .B1(_05028_),
    .B2(_04328_),
    .C1(\adder_inst.fraction1_32neg[2] ),
    .X(_03102_));
 sky130_fd_sc_hd__o22ai_1 _09082_ (.A1(\adder_inst.fraction1_32neg[2] ),
    .A2(_05034_),
    .B1(_03097_),
    .B2(_03101_),
    .Y(_03103_));
 sky130_fd_sc_hd__nand2_1 _09083_ (.A(_03096_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__or2_1 _09084_ (.A(_01296_),
    .B(_04612_),
    .X(_03105_));
 sky130_fd_sc_hd__o211ai_1 _09085_ (.A1(_01296_),
    .A2(_04612_),
    .B1(_03096_),
    .C1(_03103_),
    .Y(_03106_));
 sky130_fd_sc_hd__o21ai_1 _09086_ (.A1(\adder_inst.fraction1_32neg[3] ),
    .A2(_04623_),
    .B1(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__and2_1 _09087_ (.A(_05051_),
    .B(\adder_inst.fraction1_32neg[6] ),
    .X(_03108_));
 sky130_fd_sc_hd__nand2_1 _09088_ (.A(_05051_),
    .B(\adder_inst.fraction1_32neg[6] ),
    .Y(_03109_));
 sky130_fd_sc_hd__nor2_1 _09089_ (.A(\adder_inst.fraction1_32neg[6] ),
    .B(_05051_),
    .Y(_03111_));
 sky130_fd_sc_hd__nor2_1 _09090_ (.A(\adder_inst.fraction1_32neg[4] ),
    .B(_04339_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(_04339_),
    .B(\adder_inst.fraction1_32neg[4] ),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2b_1 _09092_ (.A_N(_03112_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__a22oi_1 _09093_ (.A1(_04339_),
    .A2(\adder_inst.fraction1_32neg[4] ),
    .B1(_03106_),
    .B2(_03094_),
    .Y(_03115_));
 sky130_fd_sc_hd__a211oi_2 _09094_ (.A1(_03107_),
    .A2(_03113_),
    .B1(_03112_),
    .C1(_01307_),
    .Y(_03116_));
 sky130_fd_sc_hd__o21bai_1 _09095_ (.A1(_03112_),
    .A2(_03115_),
    .B1_N(\adder_inst.fraction1_32neg[5] ),
    .Y(_03117_));
 sky130_fd_sc_hd__and2b_1 _09096_ (.A_N(_03116_),
    .B(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__and3b_1 _09097_ (.A_N(_03116_),
    .B(_03117_),
    .C(_03814_),
    .X(_03119_));
 sky130_fd_sc_hd__a21oi_1 _09098_ (.A1(_03117_),
    .A2(_03814_),
    .B1(_03116_),
    .Y(_03120_));
 sky130_fd_sc_hd__o21ai_1 _09099_ (.A1(_03111_),
    .A2(_03120_),
    .B1(_03109_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_2 _09100_ (.A(_03122_),
    .B(\adder_inst.fraction1_32neg[7] ),
    .Y(_03123_));
 sky130_fd_sc_hd__o211ai_2 _09101_ (.A1(_03111_),
    .A2(_03120_),
    .B1(_01318_),
    .C1(_03109_),
    .Y(_03124_));
 sky130_fd_sc_hd__o21ai_2 _09102_ (.A1(_05060_),
    .A2(_05061_),
    .B1(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__or2_1 _09103_ (.A(\adder_inst.fraction1_32neg[10] ),
    .B(_05079_),
    .X(_03126_));
 sky130_fd_sc_hd__nor2_2 _09104_ (.A(_01340_),
    .B(_05080_),
    .Y(_03127_));
 sky130_fd_sc_hd__nand2_1 _09105_ (.A(_05079_),
    .B(\adder_inst.fraction1_32neg[10] ),
    .Y(_03128_));
 sky130_fd_sc_hd__nand2_1 _09106_ (.A(_03126_),
    .B(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__nor2_1 _09107_ (.A(\adder_inst.fraction1_32neg[8] ),
    .B(_05099_),
    .Y(_03130_));
 sky130_fd_sc_hd__or2_1 _09108_ (.A(\adder_inst.fraction1_32neg[8] ),
    .B(_05099_),
    .X(_03131_));
 sky130_fd_sc_hd__nand2_1 _09109_ (.A(_05099_),
    .B(\adder_inst.fraction1_32neg[8] ),
    .Y(_03133_));
 sky130_fd_sc_hd__nand2_1 _09110_ (.A(_03131_),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__o211ai_2 _09111_ (.A1(_01329_),
    .A2(_05100_),
    .B1(_03123_),
    .C1(_03125_),
    .Y(_03135_));
 sky130_fd_sc_hd__a31oi_2 _09112_ (.A1(_03123_),
    .A2(_03125_),
    .A3(_03133_),
    .B1(_03130_),
    .Y(_03136_));
 sky130_fd_sc_hd__nand2_2 _09113_ (.A(\adder_inst.fraction1_32neg[9] ),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__a21oi_1 _09114_ (.A1(_03131_),
    .A2(_03135_),
    .B1(\adder_inst.fraction1_32neg[9] ),
    .Y(_03138_));
 sky130_fd_sc_hd__a21o_1 _09115_ (.A1(_03131_),
    .A2(_03135_),
    .B1(\adder_inst.fraction1_32neg[9] ),
    .X(_03139_));
 sky130_fd_sc_hd__a31oi_1 _09116_ (.A1(_03135_),
    .A2(\adder_inst.fraction1_32neg[9] ),
    .A3(_03131_),
    .B1(_05112_),
    .Y(_03140_));
 sky130_fd_sc_hd__o21ai_2 _09117_ (.A1(\adder_inst.fraction1_32neg[9] ),
    .A2(_03136_),
    .B1(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__o21ai_2 _09118_ (.A1(_05112_),
    .A2(_03138_),
    .B1(_03137_),
    .Y(_03142_));
 sky130_fd_sc_hd__a22oi_4 _09119_ (.A1(_05080_),
    .A2(_01340_),
    .B1(_03141_),
    .B2(_03137_),
    .Y(_03144_));
 sky130_fd_sc_hd__o21ai_1 _09120_ (.A1(\adder_inst.fraction1_32neg[10] ),
    .A2(_05079_),
    .B1(_03142_),
    .Y(_03145_));
 sky130_fd_sc_hd__a21oi_1 _09121_ (.A1(_03126_),
    .A2(_03142_),
    .B1(_03127_),
    .Y(_03146_));
 sky130_fd_sc_hd__a21oi_2 _09122_ (.A1(_03128_),
    .A2(_03145_),
    .B1(_01351_),
    .Y(_03147_));
 sky130_fd_sc_hd__o21ai_1 _09123_ (.A1(_03127_),
    .A2(_03144_),
    .B1(\adder_inst.fraction1_32neg[11] ),
    .Y(_03148_));
 sky130_fd_sc_hd__o211ai_1 _09124_ (.A1(_05080_),
    .A2(_01340_),
    .B1(_01351_),
    .C1(_03145_),
    .Y(_03149_));
 sky130_fd_sc_hd__o31a_1 _09125_ (.A1(\adder_inst.fraction1_32neg[11] ),
    .A2(_03127_),
    .A3(_03144_),
    .B1(_05091_),
    .X(_03150_));
 sky130_fd_sc_hd__o31ai_4 _09126_ (.A1(\adder_inst.fraction1_32neg[11] ),
    .A2(_03127_),
    .A3(_03144_),
    .B1(_05091_),
    .Y(_03151_));
 sky130_fd_sc_hd__nor2_1 _09127_ (.A(\adder_inst.fraction1_32neg[12] ),
    .B(_05125_),
    .Y(_03152_));
 sky130_fd_sc_hd__or2_2 _09128_ (.A(\adder_inst.fraction1_32neg[12] ),
    .B(_05125_),
    .X(_03153_));
 sky130_fd_sc_hd__nand2_2 _09129_ (.A(_05125_),
    .B(\adder_inst.fraction1_32neg[12] ),
    .Y(_03155_));
 sky130_fd_sc_hd__and2_1 _09130_ (.A(_03153_),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__nor2_1 _09131_ (.A(_01362_),
    .B(_05134_),
    .Y(_03157_));
 sky130_fd_sc_hd__nand2_1 _09132_ (.A(_05133_),
    .B(\adder_inst.fraction1_32neg[14] ),
    .Y(_03158_));
 sky130_fd_sc_hd__nor2_1 _09133_ (.A(\adder_inst.fraction1_32neg[14] ),
    .B(_05133_),
    .Y(_03159_));
 sky130_fd_sc_hd__or2_1 _09134_ (.A(\adder_inst.fraction1_32neg[14] ),
    .B(_05133_),
    .X(_03160_));
 sky130_fd_sc_hd__a221oi_1 _09135_ (.A1(\adder_inst.fraction1_32neg[12] ),
    .A2(_05125_),
    .B1(_03149_),
    .B2(_05091_),
    .C1(_03147_),
    .Y(_03161_));
 sky130_fd_sc_hd__o211ai_4 _09136_ (.A1(_03146_),
    .A2(_01351_),
    .B1(_03155_),
    .C1(_03151_),
    .Y(_03162_));
 sky130_fd_sc_hd__a31oi_2 _09137_ (.A1(_03148_),
    .A2(_03151_),
    .A3(_03155_),
    .B1(_03152_),
    .Y(_03163_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(\adder_inst.fraction1_32neg[13] ),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__a21oi_1 _09139_ (.A1(_03153_),
    .A2(_03162_),
    .B1(\adder_inst.fraction1_32neg[13] ),
    .Y(_03166_));
 sky130_fd_sc_hd__o21bai_2 _09140_ (.A1(_03152_),
    .A2(_03161_),
    .B1_N(\adder_inst.fraction1_32neg[13] ),
    .Y(_03167_));
 sky130_fd_sc_hd__a31oi_4 _09141_ (.A1(_03162_),
    .A2(\adder_inst.fraction1_32neg[13] ),
    .A3(_03153_),
    .B1(_05149_),
    .Y(_03168_));
 sky130_fd_sc_hd__o21ai_2 _09142_ (.A1(\adder_inst.fraction1_32neg[13] ),
    .A2(_03163_),
    .B1(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__a32oi_4 _09143_ (.A1(\adder_inst.fraction1_32neg[13] ),
    .A2(_03153_),
    .A3(_03162_),
    .B1(_03167_),
    .B2(_03168_),
    .Y(_03170_));
 sky130_fd_sc_hd__o21ai_1 _09144_ (.A1(_05149_),
    .A2(_03166_),
    .B1(_03164_),
    .Y(_03171_));
 sky130_fd_sc_hd__a22oi_2 _09145_ (.A1(_05134_),
    .A2(_01362_),
    .B1(_03169_),
    .B2(_03164_),
    .Y(_03172_));
 sky130_fd_sc_hd__o21ai_1 _09146_ (.A1(\adder_inst.fraction1_32neg[14] ),
    .A2(_05133_),
    .B1(_03171_),
    .Y(_03173_));
 sky130_fd_sc_hd__a21oi_1 _09147_ (.A1(_03160_),
    .A2(_03171_),
    .B1(_03157_),
    .Y(_03174_));
 sky130_fd_sc_hd__a21oi_2 _09148_ (.A1(_03158_),
    .A2(_03173_),
    .B1(_01373_),
    .Y(_03175_));
 sky130_fd_sc_hd__o21ai_1 _09149_ (.A1(_03157_),
    .A2(_03172_),
    .B1(\adder_inst.fraction1_32neg[15] ),
    .Y(_03177_));
 sky130_fd_sc_hd__o211ai_2 _09150_ (.A1(_03159_),
    .A2(_03170_),
    .B1(_01373_),
    .C1(_03158_),
    .Y(_03178_));
 sky130_fd_sc_hd__o31a_1 _09151_ (.A1(\adder_inst.fraction1_32neg[15] ),
    .A2(_03157_),
    .A3(_03172_),
    .B1(_05140_),
    .X(_03179_));
 sky130_fd_sc_hd__o31ai_1 _09152_ (.A1(\adder_inst.fraction1_32neg[15] ),
    .A2(_03157_),
    .A3(_03172_),
    .B1(_05140_),
    .Y(_03180_));
 sky130_fd_sc_hd__a21oi_1 _09153_ (.A1(_05140_),
    .A2(_03178_),
    .B1(_03175_),
    .Y(_03181_));
 sky130_fd_sc_hd__and2_1 _09154_ (.A(_05187_),
    .B(\adder_inst.fraction1_32neg[16] ),
    .X(_03182_));
 sky130_fd_sc_hd__nand2_1 _09155_ (.A(_05187_),
    .B(\adder_inst.fraction1_32neg[16] ),
    .Y(_03183_));
 sky130_fd_sc_hd__a211oi_1 _09156_ (.A1(_05140_),
    .A2(_03178_),
    .B1(_03182_),
    .C1(_03175_),
    .Y(_03184_));
 sky130_fd_sc_hd__o211ai_2 _09157_ (.A1(_03174_),
    .A2(_01373_),
    .B1(_03183_),
    .C1(_03180_),
    .Y(_03185_));
 sky130_fd_sc_hd__o311a_1 _09158_ (.A1(_03175_),
    .A2(_03179_),
    .A3(_03182_),
    .B1(_03093_),
    .C1(\adder_inst.fraction1_32neg[17] ),
    .X(_03186_));
 sky130_fd_sc_hd__or3b_1 _09159_ (.A(_03092_),
    .B(_03184_),
    .C_N(\adder_inst.fraction1_32neg[17] ),
    .X(_03188_));
 sky130_fd_sc_hd__o21bai_2 _09160_ (.A1(_03092_),
    .A2(_03184_),
    .B1_N(\adder_inst.fraction1_32neg[17] ),
    .Y(_03189_));
 sky130_fd_sc_hd__a31oi_2 _09161_ (.A1(_03185_),
    .A2(\adder_inst.fraction1_32neg[17] ),
    .A3(_03093_),
    .B1(_05181_),
    .Y(_03190_));
 sky130_fd_sc_hd__a21oi_2 _09162_ (.A1(_03189_),
    .A2(_03190_),
    .B1(_03186_),
    .Y(_03191_));
 sky130_fd_sc_hd__a32o_1 _09163_ (.A1(\adder_inst.fraction1_32neg[17] ),
    .A2(_03093_),
    .A3(_03185_),
    .B1(_03189_),
    .B2(_03190_),
    .X(_03192_));
 sky130_fd_sc_hd__o21a_1 _09164_ (.A1(_03091_),
    .A2(_03191_),
    .B1(_03090_),
    .X(_03193_));
 sky130_fd_sc_hd__xor2_1 _09165_ (.A(\adder_inst.fraction1_32neg[17] ),
    .B(_05181_),
    .X(_03194_));
 sky130_fd_sc_hd__nor2_1 _09166_ (.A(_03089_),
    .B(_03091_),
    .Y(_03195_));
 sky130_fd_sc_hd__or4b_1 _09167_ (.A(_03092_),
    .B(_03182_),
    .C(_03194_),
    .D_N(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__a21boi_2 _09168_ (.A1(\adder_inst.fraction1_32neg[19] ),
    .A2(_05171_),
    .B1_N(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__o211a_1 _09169_ (.A1(_03091_),
    .A2(_03191_),
    .B1(_03197_),
    .C1(_03090_),
    .X(_03199_));
 sky130_fd_sc_hd__o211ai_4 _09170_ (.A1(_03091_),
    .A2(_03191_),
    .B1(_03197_),
    .C1(_03090_),
    .Y(_03200_));
 sky130_fd_sc_hd__xnor2_2 _09171_ (.A(\adder_inst.fraction1_32neg[19] ),
    .B(_05171_),
    .Y(_03201_));
 sky130_fd_sc_hd__nor4_1 _09172_ (.A(_03196_),
    .B(_03201_),
    .C(_03175_),
    .D(_03179_),
    .Y(_03202_));
 sky130_fd_sc_hd__inv_2 _09173_ (.A(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__o21a_2 _09174_ (.A1(\adder_inst.fraction1_32neg[19] ),
    .A2(_05171_),
    .B1(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__inv_2 _09175_ (.A(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_1 _09176_ (.A(_03200_),
    .B(_03204_),
    .Y(_03206_));
 sky130_fd_sc_hd__o2111a_1 _09177_ (.A1(\adder_inst.fraction1_32neg[19] ),
    .A2(_05171_),
    .B1(\adder_inst.fraction1_32neg[20] ),
    .C1(_03203_),
    .D1(_03200_),
    .X(_03207_));
 sky130_fd_sc_hd__o2111ai_4 _09178_ (.A1(\adder_inst.fraction1_32neg[19] ),
    .A2(_05171_),
    .B1(\adder_inst.fraction1_32neg[20] ),
    .C1(_03203_),
    .D1(_03200_),
    .Y(_03208_));
 sky130_fd_sc_hd__a21oi_4 _09179_ (.A1(_03200_),
    .A2(_03204_),
    .B1(\adder_inst.fraction1_32neg[20] ),
    .Y(_03210_));
 sky130_fd_sc_hd__a21o_1 _09180_ (.A1(_03200_),
    .A2(_03204_),
    .B1(\adder_inst.fraction1_32neg[20] ),
    .X(_03211_));
 sky130_fd_sc_hd__a22oi_1 _09181_ (.A1(_05215_),
    .A2(_05217_),
    .B1(_03206_),
    .B2(_01384_),
    .Y(_03212_));
 sky130_fd_sc_hd__o32ai_4 _09182_ (.A1(_01384_),
    .A2(_03199_),
    .A3(_03205_),
    .B1(_05219_),
    .B2(_03210_),
    .Y(_03213_));
 sky130_fd_sc_hd__o211a_1 _09183_ (.A1(_05219_),
    .A2(_03210_),
    .B1(_03208_),
    .C1(_01395_),
    .X(_03214_));
 sky130_fd_sc_hd__o211ai_2 _09184_ (.A1(_05219_),
    .A2(_03210_),
    .B1(_03208_),
    .C1(_01395_),
    .Y(_03215_));
 sky130_fd_sc_hd__o21a_1 _09185_ (.A1(_03207_),
    .A2(_03212_),
    .B1(\adder_inst.fraction1_32neg[21] ),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_1 _09186_ (.A(_03213_),
    .B(\adder_inst.fraction1_32neg[21] ),
    .Y(_03217_));
 sky130_fd_sc_hd__a22oi_2 _09187_ (.A1(_05201_),
    .A2(_05202_),
    .B1(_03213_),
    .B2(\adder_inst.fraction1_32neg[21] ),
    .Y(_03218_));
 sky130_fd_sc_hd__o21ai_1 _09188_ (.A1(\adder_inst.fraction1_32neg[21] ),
    .A2(_03213_),
    .B1(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__a2bb2oi_1 _09189_ (.A1_N(_05199_),
    .A2_N(_05200_),
    .B1(_03215_),
    .B2(_03217_),
    .Y(_03221_));
 sky130_fd_sc_hd__o22ai_1 _09190_ (.A1(_05199_),
    .A2(_05200_),
    .B1(_03214_),
    .B2(_03216_),
    .Y(_03222_));
 sky130_fd_sc_hd__a211oi_4 _09191_ (.A1(_03215_),
    .A2(_03218_),
    .B1(_05231_),
    .C1(_03221_),
    .Y(_03223_));
 sky130_fd_sc_hd__nand3_2 _09192_ (.A(_03222_),
    .B(_05230_),
    .C(_03219_),
    .Y(_03224_));
 sky130_fd_sc_hd__o211a_1 _09193_ (.A1(net11),
    .A2(_02077_),
    .B1(\adder_inst.fraction2_32neg[19] ),
    .C1(_05172_),
    .X(_03225_));
 sky130_fd_sc_hd__nand2_2 _09194_ (.A(_05174_),
    .B(\adder_inst.fraction2_32neg[19] ),
    .Y(_03226_));
 sky130_fd_sc_hd__nor2_2 _09195_ (.A(_01483_),
    .B(_05165_),
    .Y(_03227_));
 sky130_fd_sc_hd__nor2_1 _09196_ (.A(\adder_inst.fraction2_32neg[18] ),
    .B(_05164_),
    .Y(_03228_));
 sky130_fd_sc_hd__nor2_1 _09197_ (.A(_01472_),
    .B(_05186_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(_05185_),
    .B(\adder_inst.fraction2_32neg[16] ),
    .Y(_03230_));
 sky130_fd_sc_hd__nand2_1 _09199_ (.A(_05135_),
    .B(\adder_inst.fraction2_32neg[14] ),
    .Y(_03232_));
 sky130_fd_sc_hd__nor2_1 _09200_ (.A(\adder_inst.fraction2_32neg[12] ),
    .B(_05124_),
    .Y(_03233_));
 sky130_fd_sc_hd__or2_1 _09201_ (.A(\adder_inst.fraction2_32neg[6] ),
    .B(_05049_),
    .X(_03234_));
 sky130_fd_sc_hd__o21a_1 _09202_ (.A1(_03836_),
    .A2(_03869_),
    .B1(_01428_),
    .X(_03235_));
 sky130_fd_sc_hd__a221o_1 _09203_ (.A1(net27),
    .A2(_02088_),
    .B1(_04295_),
    .B2(_03902_),
    .C1(\adder_inst.fraction2_32neg[4] ),
    .X(_03236_));
 sky130_fd_sc_hd__nand2_1 _09204_ (.A(\adder_inst.fraction2_32neg[3] ),
    .B(_04634_),
    .Y(_03237_));
 sky130_fd_sc_hd__a221o_1 _09205_ (.A1(net23),
    .A2(_02088_),
    .B1(_05028_),
    .B2(_03902_),
    .C1(\adder_inst.fraction2_32neg[2] ),
    .X(_03238_));
 sky130_fd_sc_hd__a21oi_1 _09206_ (.A1(_04962_),
    .A2(_04969_),
    .B1(\adder_inst.fraction2_32neg[1] ),
    .Y(_03239_));
 sky130_fd_sc_hd__a32oi_2 _09207_ (.A1(\adder_inst.fraction2_32neg[1] ),
    .A2(_04962_),
    .A3(_04969_),
    .B1(\adder_inst.fraction1[0] ),
    .B2(\adder_inst.fraction2_32neg[0] ),
    .Y(_03240_));
 sky130_fd_sc_hd__a21oi_1 _09208_ (.A1(_01406_),
    .A2(_04979_),
    .B1(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__o2bb2ai_1 _09209_ (.A1_N(\adder_inst.fraction2_32neg[2] ),
    .A2_N(_05032_),
    .B1(_03239_),
    .B2(_03240_),
    .Y(_03243_));
 sky130_fd_sc_hd__o31a_1 _09210_ (.A1(\adder_inst.fraction2_32neg[2] ),
    .A2(_05008_),
    .A3(_05029_),
    .B1(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__nand2b_1 _09211_ (.A_N(\adder_inst.fraction2_32neg[3] ),
    .B(_04645_),
    .Y(_03245_));
 sky130_fd_sc_hd__o21bai_1 _09212_ (.A1(_05008_),
    .A2(_05029_),
    .B1_N(\adder_inst.fraction2_32neg[2] ),
    .Y(_03246_));
 sky130_fd_sc_hd__nand3_1 _09213_ (.A(_05030_),
    .B(\adder_inst.fraction2_32neg[2] ),
    .C(_05009_),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _09214_ (.A(_03246_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__a221oi_2 _09215_ (.A1(_01241_),
    .A2(_02088_),
    .B1(_04930_),
    .B2(_03847_),
    .C1(\adder_inst.fraction2_32neg[1] ),
    .Y(_03249_));
 sky130_fd_sc_hd__a21oi_1 _09216_ (.A1(_04962_),
    .A2(_04969_),
    .B1(_01406_),
    .Y(_03250_));
 sky130_fd_sc_hd__o2111ai_2 _09217_ (.A1(_03249_),
    .A2(_03250_),
    .B1(_03004_),
    .C1(_03005_),
    .D1(_03248_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand4_1 _09218_ (.A(_03238_),
    .B(_03243_),
    .C(_03245_),
    .D(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__nand2_1 _09219_ (.A(_03237_),
    .B(_03245_),
    .Y(_03254_));
 sky130_fd_sc_hd__o21a_1 _09220_ (.A1(_04634_),
    .A2(_03244_),
    .B1(\adder_inst.fraction2_32neg[3] ),
    .X(_03255_));
 sky130_fd_sc_hd__a31o_1 _09221_ (.A1(_04634_),
    .A2(_03238_),
    .A3(_03243_),
    .B1(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__nand2_1 _09222_ (.A(_04317_),
    .B(\adder_inst.fraction2_32neg[4] ),
    .Y(_03257_));
 sky130_fd_sc_hd__o211ai_1 _09223_ (.A1(_01417_),
    .A2(_04306_),
    .B1(_03237_),
    .C1(_03252_),
    .Y(_03258_));
 sky130_fd_sc_hd__o21ai_1 _09224_ (.A1(\adder_inst.fraction2_32neg[4] ),
    .A2(_04317_),
    .B1(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__a211o_1 _09225_ (.A1(_03770_),
    .A2(_03847_),
    .B1(_03836_),
    .C1(_01428_),
    .X(_03260_));
 sky130_fd_sc_hd__a2bb2oi_1 _09226_ (.A1_N(_01428_),
    .A2_N(_03891_),
    .B1(_03236_),
    .B2(_03258_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand2_1 _09227_ (.A(_05049_),
    .B(\adder_inst.fraction2_32neg[6] ),
    .Y(_03262_));
 sky130_fd_sc_hd__o22ai_2 _09228_ (.A1(_01439_),
    .A2(_05050_),
    .B1(_03235_),
    .B2(_03261_),
    .Y(_03263_));
 sky130_fd_sc_hd__and3_1 _09229_ (.A(_05069_),
    .B(_03234_),
    .C(_03263_),
    .X(_03265_));
 sky130_fd_sc_hd__o211ai_1 _09230_ (.A1(\adder_inst.fraction2_32neg[6] ),
    .A2(_05049_),
    .B1(_05069_),
    .C1(_03263_),
    .Y(_03266_));
 sky130_fd_sc_hd__a2bb2oi_1 _09231_ (.A1_N(_05066_),
    .A2_N(_05067_),
    .B1(_03234_),
    .B2(_03263_),
    .Y(_03267_));
 sky130_fd_sc_hd__nor2_1 _09232_ (.A(_03265_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_1 _09233_ (.A(_03236_),
    .B(_03257_),
    .Y(_03269_));
 sky130_fd_sc_hd__xor2_1 _09234_ (.A(_01450_),
    .B(_05069_),
    .X(_03270_));
 sky130_fd_sc_hd__nand2b_1 _09235_ (.A_N(_03235_),
    .B(_03260_),
    .Y(_03271_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(_03234_),
    .B(_03262_),
    .Y(_03272_));
 sky130_fd_sc_hd__or4_2 _09237_ (.A(_03269_),
    .B(_03270_),
    .C(_03271_),
    .D(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__o211ai_2 _09238_ (.A1(_01450_),
    .A2(_03267_),
    .B1(_03273_),
    .C1(_03266_),
    .Y(_03274_));
 sky130_fd_sc_hd__a211o_1 _09239_ (.A1(_04634_),
    .A2(_03244_),
    .B1(_03255_),
    .C1(_03273_),
    .X(_03276_));
 sky130_fd_sc_hd__o21ai_1 _09240_ (.A1(_03256_),
    .A2(_03273_),
    .B1(_03274_),
    .Y(_03277_));
 sky130_fd_sc_hd__inv_2 _09241_ (.A(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__nor2_1 _09242_ (.A(\adder_inst.fraction2_32neg[11] ),
    .B(_05089_),
    .Y(_03279_));
 sky130_fd_sc_hd__and2_1 _09243_ (.A(_05089_),
    .B(\adder_inst.fraction2_32neg[11] ),
    .X(_03280_));
 sky130_fd_sc_hd__or2_1 _09244_ (.A(_03279_),
    .B(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__xor2_1 _09245_ (.A(\adder_inst.fraction2_32neg[9] ),
    .B(_05110_),
    .X(_03282_));
 sky130_fd_sc_hd__nor2_1 _09246_ (.A(\adder_inst.fraction2_32neg[10] ),
    .B(_05077_),
    .Y(_03283_));
 sky130_fd_sc_hd__nand2_1 _09247_ (.A(_05077_),
    .B(\adder_inst.fraction2_32neg[10] ),
    .Y(_03284_));
 sky130_fd_sc_hd__inv_2 _09248_ (.A(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__or2_1 _09249_ (.A(_03283_),
    .B(_03285_),
    .X(_03287_));
 sky130_fd_sc_hd__nor2_1 _09250_ (.A(\adder_inst.fraction2_32neg[8] ),
    .B(_05097_),
    .Y(_03288_));
 sky130_fd_sc_hd__and2_1 _09251_ (.A(_05097_),
    .B(\adder_inst.fraction2_32neg[8] ),
    .X(_03289_));
 sky130_fd_sc_hd__or2_1 _09252_ (.A(_03288_),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__or4_2 _09253_ (.A(_03281_),
    .B(_03282_),
    .C(_03287_),
    .D(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__a21o_1 _09254_ (.A1(_03274_),
    .A2(_03276_),
    .B1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__a22oi_2 _09255_ (.A1(\adder_inst.fraction2_32neg[8] ),
    .A2(_05097_),
    .B1(_03274_),
    .B2(_03276_),
    .Y(_03293_));
 sky130_fd_sc_hd__nor3_1 _09256_ (.A(_05110_),
    .B(_03288_),
    .C(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__or4_1 _09257_ (.A(_05108_),
    .B(_05109_),
    .C(_03288_),
    .D(_03293_),
    .X(_03295_));
 sky130_fd_sc_hd__o22ai_2 _09258_ (.A1(_05108_),
    .A2(_05109_),
    .B1(_03288_),
    .B2(_03293_),
    .Y(_03296_));
 sky130_fd_sc_hd__o31a_1 _09259_ (.A1(_05110_),
    .A2(_03288_),
    .A3(_03293_),
    .B1(\adder_inst.fraction2_32neg[9] ),
    .X(_03298_));
 sky130_fd_sc_hd__a21oi_1 _09260_ (.A1(_03296_),
    .A2(\adder_inst.fraction2_32neg[9] ),
    .B1(_03294_),
    .Y(_03299_));
 sky130_fd_sc_hd__nor2_1 _09261_ (.A(_03283_),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__o21a_1 _09262_ (.A1(_03283_),
    .A2(_03299_),
    .B1(_03284_),
    .X(_03301_));
 sky130_fd_sc_hd__o22ai_1 _09263_ (.A1(\adder_inst.fraction2_32neg[11] ),
    .A2(_05089_),
    .B1(_03285_),
    .B2(_03300_),
    .Y(_03302_));
 sky130_fd_sc_hd__a21bo_1 _09264_ (.A1(\adder_inst.fraction2_32neg[11] ),
    .A2(_05089_),
    .B1_N(_03291_),
    .X(_03303_));
 sky130_fd_sc_hd__inv_2 _09265_ (.A(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__o21bai_1 _09266_ (.A1(_03279_),
    .A2(_03301_),
    .B1_N(_03303_),
    .Y(_03305_));
 sky130_fd_sc_hd__o2bb2ai_2 _09267_ (.A1_N(_03304_),
    .A2_N(_03302_),
    .B1(_03291_),
    .B2(_03278_),
    .Y(_03306_));
 sky130_fd_sc_hd__nand2_1 _09268_ (.A(_05124_),
    .B(\adder_inst.fraction2_32neg[12] ),
    .Y(_03307_));
 sky130_fd_sc_hd__a22oi_1 _09269_ (.A1(_05124_),
    .A2(\adder_inst.fraction2_32neg[12] ),
    .B1(_03305_),
    .B2(_03292_),
    .Y(_03309_));
 sky130_fd_sc_hd__a221oi_2 _09270_ (.A1(_05150_),
    .A2(_05151_),
    .B1(_03306_),
    .B2(_03307_),
    .C1(_03233_),
    .Y(_03310_));
 sky130_fd_sc_hd__o22ai_1 _09271_ (.A1(_05152_),
    .A2(_05153_),
    .B1(_03233_),
    .B2(_03309_),
    .Y(_03311_));
 sky130_fd_sc_hd__and2b_1 _09272_ (.A_N(_03310_),
    .B(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__nand2_1 _09273_ (.A(\adder_inst.fraction2_32neg[13] ),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__a21oi_2 _09274_ (.A1(_03311_),
    .A2(\adder_inst.fraction2_32neg[13] ),
    .B1(_03310_),
    .Y(_03314_));
 sky130_fd_sc_hd__nor2_1 _09275_ (.A(\adder_inst.fraction2_32neg[14] ),
    .B(_05135_),
    .Y(_03315_));
 sky130_fd_sc_hd__or2_1 _09276_ (.A(\adder_inst.fraction2_32neg[14] ),
    .B(_05135_),
    .X(_03316_));
 sky130_fd_sc_hd__o21a_1 _09277_ (.A1(_03314_),
    .A2(_03315_),
    .B1(_03232_),
    .X(_03317_));
 sky130_fd_sc_hd__o221ai_2 _09278_ (.A1(_05142_),
    .A2(_01461_),
    .B1(_03315_),
    .B2(_03314_),
    .C1(_03232_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2b_1 _09279_ (.A_N(_03233_),
    .B(_03307_),
    .Y(_03320_));
 sky130_fd_sc_hd__xor2_1 _09280_ (.A(\adder_inst.fraction2_32neg[15] ),
    .B(_05142_),
    .X(_03321_));
 sky130_fd_sc_hd__nand2_1 _09281_ (.A(_03232_),
    .B(_03316_),
    .Y(_03322_));
 sky130_fd_sc_hd__nor2_1 _09282_ (.A(\adder_inst.fraction2_32neg[13] ),
    .B(_05155_),
    .Y(_03323_));
 sky130_fd_sc_hd__or3_1 _09283_ (.A(_03320_),
    .B(_03323_),
    .C(_03321_),
    .X(_03324_));
 sky130_fd_sc_hd__a211oi_1 _09284_ (.A1(\adder_inst.fraction2_32neg[13] ),
    .A2(_05155_),
    .B1(_03322_),
    .C1(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__inv_2 _09285_ (.A(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__a21oi_1 _09286_ (.A1(_01461_),
    .A2(_05142_),
    .B1(_03325_),
    .Y(_03327_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_03318_),
    .B(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__or2_1 _09288_ (.A(_03306_),
    .B(_03326_),
    .X(_03329_));
 sky130_fd_sc_hd__o2bb2ai_1 _09289_ (.A1_N(_03327_),
    .A2_N(_03318_),
    .B1(_03306_),
    .B2(_03326_),
    .Y(_03331_));
 sky130_fd_sc_hd__or2_1 _09290_ (.A(\adder_inst.fraction2_32neg[16] ),
    .B(_05185_),
    .X(_03332_));
 sky130_fd_sc_hd__a22oi_1 _09291_ (.A1(_01472_),
    .A2(_05186_),
    .B1(_03328_),
    .B2(_03329_),
    .Y(_03333_));
 sky130_fd_sc_hd__o21ai_1 _09292_ (.A1(\adder_inst.fraction2_32neg[16] ),
    .A2(_05185_),
    .B1(_03331_),
    .Y(_03334_));
 sky130_fd_sc_hd__a2bb2oi_1 _09293_ (.A1_N(_05176_),
    .A2_N(_05177_),
    .B1(_03230_),
    .B2(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__o22ai_2 _09294_ (.A1(_05176_),
    .A2(_05177_),
    .B1(_03229_),
    .B2(_03333_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand3_2 _09295_ (.A(_03334_),
    .B(_05178_),
    .C(_03230_),
    .Y(_03337_));
 sky130_fd_sc_hd__and3_1 _09296_ (.A(_03336_),
    .B(_03337_),
    .C(\adder_inst.fraction2_32neg[17] ),
    .X(_03338_));
 sky130_fd_sc_hd__nand3_1 _09297_ (.A(_03336_),
    .B(_03337_),
    .C(\adder_inst.fraction2_32neg[17] ),
    .Y(_03339_));
 sky130_fd_sc_hd__a21oi_1 _09298_ (.A1(_03337_),
    .A2(\adder_inst.fraction2_32neg[17] ),
    .B1(_03335_),
    .Y(_03340_));
 sky130_fd_sc_hd__a21o_1 _09299_ (.A1(\adder_inst.fraction2_32neg[17] ),
    .A2(_03337_),
    .B1(_03335_),
    .X(_03342_));
 sky130_fd_sc_hd__a22oi_2 _09300_ (.A1(_05165_),
    .A2(_01483_),
    .B1(_03339_),
    .B2(_03336_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21bai_1 _09301_ (.A1(_03228_),
    .A2(_03340_),
    .B1_N(_03227_),
    .Y(_03344_));
 sky130_fd_sc_hd__or2_1 _09302_ (.A(\adder_inst.fraction2_32neg[19] ),
    .B(_05174_),
    .X(_03345_));
 sky130_fd_sc_hd__nor2_1 _09303_ (.A(_03227_),
    .B(_03228_),
    .Y(_03346_));
 sky130_fd_sc_hd__o22a_1 _09304_ (.A1(\adder_inst.fraction2_32neg[19] ),
    .A2(_05174_),
    .B1(_03227_),
    .B2(_03343_),
    .X(_03347_));
 sky130_fd_sc_hd__o22ai_4 _09305_ (.A1(\adder_inst.fraction2_32neg[19] ),
    .A2(_05174_),
    .B1(_03227_),
    .B2(_03343_),
    .Y(_03348_));
 sky130_fd_sc_hd__a2bb2oi_4 _09306_ (.A1_N(_05208_),
    .A2_N(_05209_),
    .B1(_03226_),
    .B2(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__o21ai_1 _09307_ (.A1(_03225_),
    .A2(_03347_),
    .B1(_05210_),
    .Y(_03350_));
 sky130_fd_sc_hd__a211oi_2 _09308_ (.A1(_03344_),
    .A2(_03345_),
    .B1(_05210_),
    .C1(_03225_),
    .Y(_03351_));
 sky130_fd_sc_hd__a31oi_2 _09309_ (.A1(_05211_),
    .A2(_03226_),
    .A3(_03348_),
    .B1(_01494_),
    .Y(_03353_));
 sky130_fd_sc_hd__a31o_1 _09310_ (.A1(_05211_),
    .A2(_03226_),
    .A3(_03348_),
    .B1(_01494_),
    .X(_03354_));
 sky130_fd_sc_hd__o22ai_4 _09311_ (.A1(_02220_),
    .A2(_05204_),
    .B1(_03349_),
    .B2(_03353_),
    .Y(_03355_));
 sky130_fd_sc_hd__o211ai_4 _09312_ (.A1(_01494_),
    .A2(_03351_),
    .B1(_03350_),
    .C1(_05205_),
    .Y(_03356_));
 sky130_fd_sc_hd__a21oi_2 _09313_ (.A1(_03355_),
    .A2(_03356_),
    .B1(\adder_inst.fraction2_32neg[21] ),
    .Y(_03357_));
 sky130_fd_sc_hd__a21o_1 _09314_ (.A1(_03355_),
    .A2(_03356_),
    .B1(\adder_inst.fraction2_32neg[21] ),
    .X(_03358_));
 sky130_fd_sc_hd__a31oi_1 _09315_ (.A1(_03355_),
    .A2(_03356_),
    .A3(\adder_inst.fraction2_32neg[21] ),
    .B1(_05230_),
    .Y(_03359_));
 sky130_fd_sc_hd__a31o_1 _09316_ (.A1(_03355_),
    .A2(_03356_),
    .A3(\adder_inst.fraction2_32neg[21] ),
    .B1(_05230_),
    .X(_03360_));
 sky130_fd_sc_hd__o21bai_4 _09317_ (.A1(_03357_),
    .A2(_03360_),
    .B1_N(net116),
    .Y(_03361_));
 sky130_fd_sc_hd__a21oi_1 _09318_ (.A1(_03358_),
    .A2(_03359_),
    .B1(net116),
    .Y(_03362_));
 sky130_fd_sc_hd__o211ai_4 _09319_ (.A1(_03357_),
    .A2(_03360_),
    .B1(net114),
    .C1(_03224_),
    .Y(_03364_));
 sky130_fd_sc_hd__a2bb2oi_4 _09320_ (.A1_N(net114),
    .A2_N(_03086_),
    .B1(_03224_),
    .B2(_03362_),
    .Y(_03365_));
 sky130_fd_sc_hd__o22ai_4 _09321_ (.A1(net114),
    .A2(_03086_),
    .B1(_03223_),
    .B2(_03361_),
    .Y(_03366_));
 sky130_fd_sc_hd__xnor2_1 _09322_ (.A(_05169_),
    .B(_03076_),
    .Y(_03367_));
 sky130_fd_sc_hd__nor2_2 _09323_ (.A(net114),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__o31a_1 _09324_ (.A1(_03089_),
    .A2(_03091_),
    .A3(_03191_),
    .B1(_05230_),
    .X(_03369_));
 sky130_fd_sc_hd__o21ai_4 _09325_ (.A1(_03192_),
    .A2(_03195_),
    .B1(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__o21ai_1 _09326_ (.A1(_03346_),
    .A2(_03342_),
    .B1(net102),
    .Y(_03371_));
 sky130_fd_sc_hd__a21o_2 _09327_ (.A1(_03342_),
    .A2(_03346_),
    .B1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__a31oi_4 _09328_ (.A1(net114),
    .A2(_03370_),
    .A3(_03372_),
    .B1(_03368_),
    .Y(_03373_));
 sky130_fd_sc_hd__a31o_4 _09329_ (.A1(net114),
    .A2(_03370_),
    .A3(_03372_),
    .B1(_03368_),
    .X(_03375_));
 sky130_fd_sc_hd__o22ai_2 _09330_ (.A1(_05212_),
    .A2(_05213_),
    .B1(_03207_),
    .B2(_03210_),
    .Y(_03376_));
 sky130_fd_sc_hd__o211ai_2 _09331_ (.A1(_05214_),
    .A2(_05216_),
    .B1(_03208_),
    .C1(_03211_),
    .Y(_03377_));
 sky130_fd_sc_hd__o21ai_1 _09332_ (.A1(_03349_),
    .A2(_03351_),
    .B1(_01494_),
    .Y(_03378_));
 sky130_fd_sc_hd__o211ai_4 _09333_ (.A1(_03354_),
    .A2(_03349_),
    .B1(_05231_),
    .C1(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__a31oi_4 _09334_ (.A1(_03376_),
    .A2(_03377_),
    .A3(_05230_),
    .B1(net116),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_4 _09335_ (.A(_03380_),
    .B(_03379_),
    .Y(_03381_));
 sky130_fd_sc_hd__inv_2 _09336_ (.A(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__o21a_1 _09337_ (.A1(_05220_),
    .A2(_05221_),
    .B1(_03081_),
    .X(_03383_));
 sky130_fd_sc_hd__o21ai_4 _09338_ (.A1(_05223_),
    .A2(_03081_),
    .B1(net116),
    .Y(_03384_));
 sky130_fd_sc_hd__a21o_4 _09339_ (.A1(_05223_),
    .A2(_03081_),
    .B1(_03384_),
    .X(_03386_));
 sky130_fd_sc_hd__inv_2 _09340_ (.A(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a2bb2oi_4 _09341_ (.A1_N(_03384_),
    .A2_N(_03383_),
    .B1(_03379_),
    .B2(_03380_),
    .Y(_03388_));
 sky130_fd_sc_hd__o2bb2ai_4 _09342_ (.A1_N(_03379_),
    .A2_N(_03380_),
    .B1(_03383_),
    .B2(_03384_),
    .Y(_03389_));
 sky130_fd_sc_hd__xor2_2 _09343_ (.A(_03193_),
    .B(_03201_),
    .X(_03390_));
 sky130_fd_sc_hd__or3_1 _09344_ (.A(_05231_),
    .B(net116),
    .C(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__o21ai_1 _09345_ (.A1(_05175_),
    .A2(_03078_),
    .B1(net116),
    .Y(_03392_));
 sky130_fd_sc_hd__a21o_2 _09346_ (.A1(_05175_),
    .A2(_03078_),
    .B1(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__and3_1 _09347_ (.A(_03226_),
    .B(_03344_),
    .C(_03345_),
    .X(_03394_));
 sky130_fd_sc_hd__a21oi_1 _09348_ (.A1(_03226_),
    .A2(_03345_),
    .B1(_03344_),
    .Y(_03395_));
 sky130_fd_sc_hd__o21ai_4 _09349_ (.A1(_03394_),
    .A2(_03395_),
    .B1(_05234_),
    .Y(_03397_));
 sky130_fd_sc_hd__o211a_2 _09350_ (.A1(_00000_),
    .A2(_03390_),
    .B1(_03393_),
    .C1(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__o211ai_4 _09351_ (.A1(_00000_),
    .A2(_03390_),
    .B1(_03393_),
    .C1(_03397_),
    .Y(_03399_));
 sky130_fd_sc_hd__a32oi_4 _09352_ (.A1(_03391_),
    .A2(_03393_),
    .A3(_03397_),
    .B1(net101),
    .B2(_03087_),
    .Y(_03400_));
 sky130_fd_sc_hd__a21oi_4 _09353_ (.A1(_03381_),
    .A2(_03386_),
    .B1(_03398_),
    .Y(_03401_));
 sky130_fd_sc_hd__a31o_2 _09354_ (.A1(_03391_),
    .A2(_03393_),
    .A3(_03397_),
    .B1(_03388_),
    .X(_03402_));
 sky130_fd_sc_hd__a21oi_4 _09355_ (.A1(_03087_),
    .A2(net101),
    .B1(_03388_),
    .Y(_03403_));
 sky130_fd_sc_hd__o2bb2ai_4 _09356_ (.A1_N(_03087_),
    .A2_N(_03364_),
    .B1(_03382_),
    .B2(_03387_),
    .Y(_03404_));
 sky130_fd_sc_hd__a21oi_4 _09357_ (.A1(_03087_),
    .A2(net101),
    .B1(_03402_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_8 _09358_ (.A(_03366_),
    .B(_03401_),
    .Y(_03406_));
 sky130_fd_sc_hd__a211oi_4 _09359_ (.A1(_03087_),
    .A2(net101),
    .B1(_03373_),
    .C1(_03402_),
    .Y(_03408_));
 sky130_fd_sc_hd__a211o_4 _09360_ (.A1(_03087_),
    .A2(net101),
    .B1(_03373_),
    .C1(_03402_),
    .X(_03409_));
 sky130_fd_sc_hd__a21oi_1 _09361_ (.A1(_03188_),
    .A2(_03189_),
    .B1(_05182_),
    .Y(_03410_));
 sky130_fd_sc_hd__a311o_1 _09362_ (.A1(_05182_),
    .A2(_03188_),
    .A3(_03189_),
    .B1(net102),
    .C1(_03410_),
    .X(_03411_));
 sky130_fd_sc_hd__a21oi_1 _09363_ (.A1(_03336_),
    .A2(_03337_),
    .B1(\adder_inst.fraction2_32neg[17] ),
    .Y(_03412_));
 sky130_fd_sc_hd__xor2_2 _09364_ (.A(_05182_),
    .B(_03075_),
    .X(_03413_));
 sky130_fd_sc_hd__o31a_1 _09365_ (.A1(_05230_),
    .A2(_03338_),
    .A3(_03412_),
    .B1(_03411_),
    .X(_03414_));
 sky130_fd_sc_hd__nor2_1 _09366_ (.A(net116),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__a21oi_4 _09367_ (.A1(net116),
    .A2(_03413_),
    .B1(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__inv_2 _09368_ (.A(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__a211o_1 _09369_ (.A1(net116),
    .A2(_03413_),
    .B1(_03415_),
    .C1(_03388_),
    .X(_03419_));
 sky130_fd_sc_hd__a21o_1 _09370_ (.A1(_03087_),
    .A2(_03364_),
    .B1(_03375_),
    .X(_03420_));
 sky130_fd_sc_hd__o211ai_4 _09371_ (.A1(_03373_),
    .A2(_03389_),
    .B1(_03419_),
    .C1(_03366_),
    .Y(_03421_));
 sky130_fd_sc_hd__a22o_1 _09372_ (.A1(net98),
    .A2(_03399_),
    .B1(_03420_),
    .B2(_03389_),
    .X(_03422_));
 sky130_fd_sc_hd__o21ai_1 _09373_ (.A1(_03406_),
    .A2(_03421_),
    .B1(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__and4_4 _09374_ (.A(net98),
    .B(_03375_),
    .C(_03401_),
    .D(_03416_),
    .X(_03424_));
 sky130_fd_sc_hd__nand4_4 _09375_ (.A(net98),
    .B(_03375_),
    .C(_03401_),
    .D(_03416_),
    .Y(_03425_));
 sky130_fd_sc_hd__a221o_1 _09376_ (.A1(_05140_),
    .A2(_03178_),
    .B1(_03183_),
    .B2(_03093_),
    .C1(_03175_),
    .X(_03426_));
 sky130_fd_sc_hd__o311a_1 _09377_ (.A1(_03092_),
    .A2(_03182_),
    .A3(_03181_),
    .B1(_05230_),
    .C1(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__nand3_1 _09378_ (.A(_03230_),
    .B(_03331_),
    .C(_03332_),
    .Y(_03428_));
 sky130_fd_sc_hd__a21o_1 _09379_ (.A1(_03230_),
    .A2(_03332_),
    .B1(_03331_),
    .X(_03430_));
 sky130_fd_sc_hd__a31o_1 _09380_ (.A1(net102),
    .A2(_03428_),
    .A3(_03430_),
    .B1(net116),
    .X(_03431_));
 sky130_fd_sc_hd__a21oi_1 _09381_ (.A1(_05188_),
    .A2(_05189_),
    .B1(_03069_),
    .Y(_03432_));
 sky130_fd_sc_hd__a311o_1 _09382_ (.A1(_05188_),
    .A2(_05189_),
    .A3(_03069_),
    .B1(net115),
    .C1(_03432_),
    .X(_03433_));
 sky130_fd_sc_hd__o21ai_4 _09383_ (.A1(_03427_),
    .A2(_03431_),
    .B1(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__inv_2 _09384_ (.A(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__a21oi_1 _09385_ (.A1(_03177_),
    .A2(_03178_),
    .B1(_05140_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21oi_1 _09386_ (.A1(_03177_),
    .A2(_03179_),
    .B1(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__xor2_1 _09387_ (.A(_05144_),
    .B(_03061_),
    .X(_03438_));
 sky130_fd_sc_hd__or2_1 _09388_ (.A(_03321_),
    .B(_03317_),
    .X(_03439_));
 sky130_fd_sc_hd__a21oi_1 _09389_ (.A1(_03317_),
    .A2(_03321_),
    .B1(_05230_),
    .Y(_03441_));
 sky130_fd_sc_hd__a221o_1 _09390_ (.A1(_03441_),
    .A2(_03439_),
    .B1(_03437_),
    .B2(_05230_),
    .C1(net116),
    .X(_03442_));
 sky130_fd_sc_hd__o21a_1 _09391_ (.A1(net115),
    .A2(_03438_),
    .B1(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__inv_2 _09392_ (.A(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__o21a_1 _09393_ (.A1(_03157_),
    .A2(_03159_),
    .B1(_03171_),
    .X(_03445_));
 sky130_fd_sc_hd__a311oi_1 _09394_ (.A1(_03158_),
    .A2(_03160_),
    .A3(_03170_),
    .B1(_03445_),
    .C1(_00000_),
    .Y(_03446_));
 sky130_fd_sc_hd__o21ai_1 _09395_ (.A1(_05138_),
    .A2(_03060_),
    .B1(net116),
    .Y(_03447_));
 sky130_fd_sc_hd__a21oi_1 _09396_ (.A1(_05138_),
    .A2(_03060_),
    .B1(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__xnor2_1 _09397_ (.A(_03314_),
    .B(_03322_),
    .Y(_03449_));
 sky130_fd_sc_hd__a311o_2 _09398_ (.A1(net102),
    .A2(net115),
    .A3(_03449_),
    .B1(_03448_),
    .C1(_03446_),
    .X(_03450_));
 sky130_fd_sc_hd__inv_2 _09399_ (.A(_03450_),
    .Y(_03452_));
 sky130_fd_sc_hd__a21o_1 _09400_ (.A1(_03164_),
    .A2(_03167_),
    .B1(_05148_),
    .X(_03453_));
 sky130_fd_sc_hd__o21a_1 _09401_ (.A1(\adder_inst.fraction2_32neg[13] ),
    .A2(_03312_),
    .B1(net102),
    .X(_03454_));
 sky130_fd_sc_hd__a32oi_4 _09402_ (.A1(_05230_),
    .A2(_03169_),
    .A3(_03453_),
    .B1(_03454_),
    .B2(_03313_),
    .Y(_03455_));
 sky130_fd_sc_hd__a21oi_1 _09403_ (.A1(_03057_),
    .A2(_03058_),
    .B1(_05148_),
    .Y(_03456_));
 sky130_fd_sc_hd__or3_1 _09404_ (.A(_03456_),
    .B(net115),
    .C(_03059_),
    .X(_03457_));
 sky130_fd_sc_hd__o21ai_1 _09405_ (.A1(net116),
    .A2(_03455_),
    .B1(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__o21ai_1 _09406_ (.A1(_03147_),
    .A2(_03150_),
    .B1(_03156_),
    .Y(_03459_));
 sky130_fd_sc_hd__o31a_1 _09407_ (.A1(_03147_),
    .A2(_03150_),
    .A3(_03156_),
    .B1(_05230_),
    .X(_03460_));
 sky130_fd_sc_hd__o21ai_1 _09408_ (.A1(_03306_),
    .A2(_03320_),
    .B1(net102),
    .Y(_03461_));
 sky130_fd_sc_hd__a21oi_1 _09409_ (.A1(_03306_),
    .A2(_03320_),
    .B1(_03461_),
    .Y(_03463_));
 sky130_fd_sc_hd__and3_1 _09410_ (.A(_03052_),
    .B(_05129_),
    .C(_03042_),
    .X(_03464_));
 sky130_fd_sc_hd__a21oi_1 _09411_ (.A1(_03042_),
    .A2(_03052_),
    .B1(_05129_),
    .Y(_03465_));
 sky130_fd_sc_hd__a211o_1 _09412_ (.A1(_03460_),
    .A2(_03459_),
    .B1(net116),
    .C1(_03463_),
    .X(_03466_));
 sky130_fd_sc_hd__o31a_2 _09413_ (.A1(net115),
    .A2(_03464_),
    .A3(_03465_),
    .B1(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__a21o_1 _09414_ (.A1(_03148_),
    .A2(_03149_),
    .B1(_05091_),
    .X(_03468_));
 sky130_fd_sc_hd__nor2_1 _09415_ (.A(_05094_),
    .B(_03049_),
    .Y(_03469_));
 sky130_fd_sc_hd__o211a_1 _09416_ (.A1(_05081_),
    .A2(_03048_),
    .B1(_05094_),
    .C1(_05082_),
    .X(_03470_));
 sky130_fd_sc_hd__o211a_1 _09417_ (.A1(_03147_),
    .A2(_03151_),
    .B1(_03468_),
    .C1(_05230_),
    .X(_03471_));
 sky130_fd_sc_hd__a21oi_1 _09418_ (.A1(_03281_),
    .A2(_03301_),
    .B1(_05230_),
    .Y(_03472_));
 sky130_fd_sc_hd__o21a_1 _09419_ (.A1(_03281_),
    .A2(_03301_),
    .B1(_03472_),
    .X(_03474_));
 sky130_fd_sc_hd__or3_1 _09420_ (.A(net116),
    .B(_03471_),
    .C(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__o31a_2 _09421_ (.A1(net115),
    .A2(_03469_),
    .A3(_03470_),
    .B1(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__a21oi_1 _09422_ (.A1(_03129_),
    .A2(_03142_),
    .B1(_00000_),
    .Y(_03477_));
 sky130_fd_sc_hd__o21a_1 _09423_ (.A1(_03129_),
    .A2(_03142_),
    .B1(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__o21ai_1 _09424_ (.A1(_05083_),
    .A2(_03048_),
    .B1(_05232_),
    .Y(_03479_));
 sky130_fd_sc_hd__a21oi_1 _09425_ (.A1(_05083_),
    .A2(_03048_),
    .B1(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__xnor2_1 _09426_ (.A(_03287_),
    .B(_03299_),
    .Y(_03481_));
 sky130_fd_sc_hd__a31o_1 _09427_ (.A1(net102),
    .A2(net115),
    .A3(_03481_),
    .B1(_03480_),
    .X(_03482_));
 sky130_fd_sc_hd__nor2_1 _09428_ (.A(_03482_),
    .B(_03478_),
    .Y(_03483_));
 sky130_fd_sc_hd__a21o_1 _09429_ (.A1(_03137_),
    .A2(_03139_),
    .B1(_05111_),
    .X(_03485_));
 sky130_fd_sc_hd__and3_1 _09430_ (.A(_05230_),
    .B(_03141_),
    .C(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__a21oi_1 _09431_ (.A1(_03295_),
    .A2(_03296_),
    .B1(\adder_inst.fraction2_32neg[9] ),
    .Y(_03487_));
 sky130_fd_sc_hd__a211o_1 _09432_ (.A1(_03296_),
    .A2(_03298_),
    .B1(_03487_),
    .C1(_05230_),
    .X(_03488_));
 sky130_fd_sc_hd__nand2_1 _09433_ (.A(_05233_),
    .B(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__xor2_1 _09434_ (.A(_05111_),
    .B(_03047_),
    .X(_03490_));
 sky130_fd_sc_hd__o22a_4 _09435_ (.A1(_05233_),
    .A2(_03490_),
    .B1(_03486_),
    .B2(_03489_),
    .X(_03491_));
 sky130_fd_sc_hd__o221a_1 _09436_ (.A1(_01252_),
    .A2(_02088_),
    .B1(_03011_),
    .B2(_03013_),
    .C1(_04936_),
    .X(_03492_));
 sky130_fd_sc_hd__or2_1 _09437_ (.A(_03014_),
    .B(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__o21ai_1 _09438_ (.A1(_04949_),
    .A2(_03100_),
    .B1(_05230_),
    .Y(_03494_));
 sky130_fd_sc_hd__a21o_1 _09439_ (.A1(_04949_),
    .A2(_03100_),
    .B1(_03494_),
    .X(_03496_));
 sky130_fd_sc_hd__o211a_1 _09440_ (.A1(_03249_),
    .A2(_03250_),
    .B1(\adder_inst.fraction2_32neg[0] ),
    .C1(\adder_inst.fraction1[0] ),
    .X(_03497_));
 sky130_fd_sc_hd__a211oi_1 _09441_ (.A1(\adder_inst.fraction2_32neg[0] ),
    .A2(\adder_inst.fraction1[0] ),
    .B1(_03249_),
    .C1(_03250_),
    .Y(_03498_));
 sky130_fd_sc_hd__o311a_1 _09442_ (.A1(_05230_),
    .A2(_03497_),
    .A3(_03498_),
    .B1(_05233_),
    .C1(_03496_),
    .X(_03499_));
 sky130_fd_sc_hd__a21oi_4 _09443_ (.A1(_05232_),
    .A2(_03493_),
    .B1(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__xnor2_1 _09444_ (.A(_03107_),
    .B(_03114_),
    .Y(_03501_));
 sky130_fd_sc_hd__and3_1 _09445_ (.A(_05230_),
    .B(_05233_),
    .C(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__o21ai_1 _09446_ (.A1(_03028_),
    .A2(_03025_),
    .B1(_05232_),
    .Y(_03503_));
 sky130_fd_sc_hd__a21oi_1 _09447_ (.A1(_03025_),
    .A2(_03028_),
    .B1(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__xor2_1 _09448_ (.A(_03256_),
    .B(_03269_),
    .X(_03505_));
 sky130_fd_sc_hd__a311oi_4 _09449_ (.A1(net102),
    .A2(_05233_),
    .A3(_03505_),
    .B1(_03504_),
    .C1(_03502_),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_1 _09450_ (.A(_03259_),
    .B(_03271_),
    .Y(_03508_));
 sky130_fd_sc_hd__xor2_1 _09451_ (.A(_03825_),
    .B(_03035_),
    .X(_03509_));
 sky130_fd_sc_hd__nor2_1 _09452_ (.A(_05233_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__nor2_1 _09453_ (.A(_03814_),
    .B(_03118_),
    .Y(_03511_));
 sky130_fd_sc_hd__o211a_1 _09454_ (.A1(_03119_),
    .A2(_03511_),
    .B1(_05233_),
    .C1(_05230_),
    .X(_03512_));
 sky130_fd_sc_hd__a311oi_4 _09455_ (.A1(net102),
    .A2(_05233_),
    .A3(_03508_),
    .B1(_03510_),
    .C1(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__xor2_1 _09456_ (.A(_03241_),
    .B(_03248_),
    .X(_03514_));
 sky130_fd_sc_hd__xnor2_1 _09457_ (.A(_03015_),
    .B(_03019_),
    .Y(_03515_));
 sky130_fd_sc_hd__or4b_1 _09458_ (.A(_03095_),
    .B(_03097_),
    .C(_03101_),
    .D_N(_03102_),
    .X(_03516_));
 sky130_fd_sc_hd__a2bb2o_1 _09459_ (.A1_N(_03097_),
    .A2_N(_03101_),
    .B1(_03102_),
    .B2(_03096_),
    .X(_03518_));
 sky130_fd_sc_hd__nand2_1 _09460_ (.A(_03516_),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__o22a_1 _09461_ (.A1(_05233_),
    .A2(_03515_),
    .B1(_03519_),
    .B2(_00000_),
    .X(_03520_));
 sky130_fd_sc_hd__o31a_2 _09462_ (.A1(_05230_),
    .A2(_05232_),
    .A3(_03514_),
    .B1(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__a21oi_1 _09463_ (.A1(_03123_),
    .A2(_03125_),
    .B1(_03134_),
    .Y(_03522_));
 sky130_fd_sc_hd__and3_1 _09464_ (.A(_03123_),
    .B(_03125_),
    .C(_03134_),
    .X(_03523_));
 sky130_fd_sc_hd__nor2_1 _09465_ (.A(_03522_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__or3_1 _09466_ (.A(_05103_),
    .B(_03038_),
    .C(_03040_),
    .X(_03525_));
 sky130_fd_sc_hd__o21ai_1 _09467_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_05103_),
    .Y(_03526_));
 sky130_fd_sc_hd__a21o_1 _09468_ (.A1(_03525_),
    .A2(_03526_),
    .B1(net115),
    .X(_03527_));
 sky130_fd_sc_hd__a21oi_1 _09469_ (.A1(_03274_),
    .A2(_03276_),
    .B1(_03290_),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_1 _09470_ (.A(_03278_),
    .B(_03290_),
    .Y(_03530_));
 sky130_fd_sc_hd__or4b_1 _09471_ (.A(_05230_),
    .B(_05232_),
    .C(_03529_),
    .D_N(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__o311a_2 _09472_ (.A1(net102),
    .A2(_05232_),
    .A3(_03524_),
    .B1(_03527_),
    .C1(_03531_),
    .X(_03532_));
 sky130_fd_sc_hd__a211oi_1 _09473_ (.A1(_01428_),
    .A2(_03891_),
    .B1(_03272_),
    .C1(_03261_),
    .Y(_03533_));
 sky130_fd_sc_hd__o21a_1 _09474_ (.A1(_03235_),
    .A2(_03261_),
    .B1(_03272_),
    .X(_03534_));
 sky130_fd_sc_hd__or2_1 _09475_ (.A(_03533_),
    .B(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__xor2_1 _09476_ (.A(_05115_),
    .B(_03036_),
    .X(_03536_));
 sky130_fd_sc_hd__o21ba_1 _09477_ (.A1(_03108_),
    .A2(_03111_),
    .B1_N(_03120_),
    .X(_03537_));
 sky130_fd_sc_hd__a2111oi_1 _09478_ (.A1(_03117_),
    .A2(_03814_),
    .B1(_03111_),
    .C1(_03116_),
    .D1(_03108_),
    .Y(_03538_));
 sky130_fd_sc_hd__o32a_1 _09479_ (.A1(_03537_),
    .A2(_03538_),
    .A3(_00000_),
    .B1(_03536_),
    .B2(_05233_),
    .X(_03540_));
 sky130_fd_sc_hd__a21boi_4 _09480_ (.A1(_05234_),
    .A2(_03535_),
    .B1_N(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(_03094_),
    .B(_03105_),
    .Y(_03542_));
 sky130_fd_sc_hd__xnor2_1 _09482_ (.A(_03104_),
    .B(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_03017_),
    .B(_03024_),
    .Y(_03544_));
 sky130_fd_sc_hd__o21a_1 _09484_ (.A1(_03017_),
    .A2(_03024_),
    .B1(_05232_),
    .X(_03545_));
 sky130_fd_sc_hd__xor2_1 _09485_ (.A(_03244_),
    .B(_03254_),
    .X(_03546_));
 sky130_fd_sc_hd__a2bb2o_1 _09486_ (.A1_N(_03543_),
    .A2_N(_00000_),
    .B1(_05234_),
    .B2(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__a21oi_4 _09487_ (.A1(_03544_),
    .A2(_03545_),
    .B1(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__o211ai_1 _09488_ (.A1(_05060_),
    .A2(_05061_),
    .B1(_03123_),
    .C1(_03124_),
    .Y(_03549_));
 sky130_fd_sc_hd__a221o_1 _09489_ (.A1(net62),
    .A2(_02077_),
    .B1(_03123_),
    .B2(_03124_),
    .C1(_05060_),
    .X(_03551_));
 sky130_fd_sc_hd__nand2_1 _09490_ (.A(_03549_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__nand2b_1 _09491_ (.A_N(_03038_),
    .B(_03039_),
    .Y(_03553_));
 sky130_fd_sc_hd__a311o_1 _09492_ (.A1(net62),
    .A2(net112),
    .A3(net109),
    .B1(_05060_),
    .C1(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__o21ai_1 _09493_ (.A1(_05060_),
    .A2(_05061_),
    .B1(_03553_),
    .Y(_03555_));
 sky130_fd_sc_hd__xor2_1 _09494_ (.A(_01450_),
    .B(_03268_),
    .X(_03556_));
 sky130_fd_sc_hd__a32o_1 _09495_ (.A1(_05232_),
    .A2(_03554_),
    .A3(_03555_),
    .B1(_05234_),
    .B2(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__a31oi_4 _09496_ (.A1(_05230_),
    .A2(net115),
    .A3(_03552_),
    .B1(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__xnor2_1 _09497_ (.A(net15),
    .B(\adder_inst.fraction2_32neg[22] ),
    .Y(_03559_));
 sky130_fd_sc_hd__a21boi_1 _09498_ (.A1(\adder_inst.fraction2_32neg[21] ),
    .A2(_03356_),
    .B1_N(_03355_),
    .Y(_03560_));
 sky130_fd_sc_hd__a21oi_1 _09499_ (.A1(_03560_),
    .A2(_03559_),
    .B1(_05230_),
    .Y(_03562_));
 sky130_fd_sc_hd__o21a_1 _09500_ (.A1(_03559_),
    .A2(_03560_),
    .B1(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__xnor2_1 _09501_ (.A(net47),
    .B(\adder_inst.fraction1_32neg[22] ),
    .Y(_03564_));
 sky130_fd_sc_hd__a21oi_1 _09502_ (.A1(_03217_),
    .A2(_03219_),
    .B1(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a31o_1 _09503_ (.A1(_03217_),
    .A2(_03219_),
    .A3(_03564_),
    .B1(_05231_),
    .X(_03566_));
 sky130_fd_sc_hd__nor2_1 _09504_ (.A(_03565_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__o21ai_1 _09505_ (.A1(_03563_),
    .A2(_03567_),
    .B1(net114),
    .Y(_03568_));
 sky130_fd_sc_hd__a22o_1 _09506_ (.A1(_05201_),
    .A2(_05202_),
    .B1(_05205_),
    .B2(_03082_),
    .X(_03569_));
 sky130_fd_sc_hd__o21ai_1 _09507_ (.A1(_05205_),
    .A2(_03082_),
    .B1(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__xnor2_1 _09508_ (.A(_05227_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__o21ai_4 _09509_ (.A1(net114),
    .A2(_03571_),
    .B1(_03568_),
    .Y(_03573_));
 sky130_fd_sc_hd__and3_1 _09510_ (.A(_03366_),
    .B(_03373_),
    .C(_03401_),
    .X(_03574_));
 sky130_fd_sc_hd__nand4_4 _09511_ (.A(net98),
    .B(_03373_),
    .C(_03389_),
    .D(_03399_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_1 _09512_ (.A(_03388_),
    .B(_03450_),
    .Y(_03576_));
 sky130_fd_sc_hd__o21ai_1 _09513_ (.A1(_03388_),
    .A2(_03458_),
    .B1(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__o211ai_2 _09514_ (.A1(_03085_),
    .A2(_03083_),
    .B1(_03444_),
    .C1(net101),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_1 _09515_ (.A(net99),
    .B(_03577_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand4_1 _09516_ (.A(net98),
    .B(_03577_),
    .C(_03401_),
    .D(_03373_),
    .Y(_03580_));
 sky130_fd_sc_hd__o211ai_1 _09517_ (.A1(net116),
    .A2(_03455_),
    .B1(_03457_),
    .C1(_03388_),
    .Y(_03581_));
 sky130_fd_sc_hd__o21ai_2 _09518_ (.A1(_03388_),
    .A2(_03467_),
    .B1(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__o211ai_1 _09519_ (.A1(net114),
    .A2(_03086_),
    .B1(_03452_),
    .C1(net101),
    .Y(_03584_));
 sky130_fd_sc_hd__nand4_1 _09520_ (.A(net98),
    .B(_03375_),
    .C(_03582_),
    .D(_03401_),
    .Y(_03585_));
 sky130_fd_sc_hd__nand2_1 _09521_ (.A(_03388_),
    .B(_03444_),
    .Y(_03586_));
 sky130_fd_sc_hd__o21ai_2 _09522_ (.A1(_03388_),
    .A2(_03452_),
    .B1(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__nand2_1 _09523_ (.A(net98),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__o221ai_4 _09524_ (.A1(net114),
    .A2(_03086_),
    .B1(_03223_),
    .B2(_03361_),
    .C1(_03434_),
    .Y(_03589_));
 sky130_fd_sc_hd__a21oi_4 _09525_ (.A1(_03588_),
    .A2(_03589_),
    .B1(_03405_),
    .Y(_03590_));
 sky130_fd_sc_hd__nand2_2 _09526_ (.A(_03580_),
    .B(_03585_),
    .Y(_03591_));
 sky130_fd_sc_hd__o21ai_2 _09527_ (.A1(_03591_),
    .A2(_03590_),
    .B1(_03425_),
    .Y(_03592_));
 sky130_fd_sc_hd__a21o_1 _09528_ (.A1(_03381_),
    .A2(_03386_),
    .B1(_03435_),
    .X(_03593_));
 sky130_fd_sc_hd__nand2_2 _09529_ (.A(_03388_),
    .B(_03416_),
    .Y(_03595_));
 sky130_fd_sc_hd__o21ai_4 _09530_ (.A1(_03388_),
    .A2(_03435_),
    .B1(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__a21oi_4 _09531_ (.A1(_03087_),
    .A2(net101),
    .B1(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__a21o_2 _09532_ (.A1(_03087_),
    .A2(net101),
    .B1(_03596_),
    .X(_03598_));
 sky130_fd_sc_hd__a31o_1 _09533_ (.A1(net98),
    .A2(_03593_),
    .A3(_03595_),
    .B1(_03409_),
    .X(_03599_));
 sky130_fd_sc_hd__nor2_8 _09534_ (.A(_03597_),
    .B(_03425_),
    .Y(_03600_));
 sky130_fd_sc_hd__a31o_4 _09535_ (.A1(net98),
    .A2(_03593_),
    .A3(_03595_),
    .B1(_03425_),
    .X(_03601_));
 sky130_fd_sc_hd__nand3b_1 _09536_ (.A_N(_03467_),
    .B(_03386_),
    .C(_03381_),
    .Y(_03602_));
 sky130_fd_sc_hd__o21ai_1 _09537_ (.A1(_03388_),
    .A2(_03476_),
    .B1(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__o211a_1 _09538_ (.A1(_03388_),
    .A2(_03476_),
    .B1(_03602_),
    .C1(_03366_),
    .X(_03604_));
 sky130_fd_sc_hd__nand4_1 _09539_ (.A(net98),
    .B(_03603_),
    .C(_03401_),
    .D(_03373_),
    .Y(_03606_));
 sky130_fd_sc_hd__o211a_1 _09540_ (.A1(_03085_),
    .A2(_03083_),
    .B1(_03467_),
    .C1(net101),
    .X(_03607_));
 sky130_fd_sc_hd__o21ai_1 _09541_ (.A1(_03478_),
    .A2(_03482_),
    .B1(_03389_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21ai_1 _09542_ (.A1(_03389_),
    .A2(_03476_),
    .B1(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__a21oi_1 _09543_ (.A1(_03087_),
    .A2(_03364_),
    .B1(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand4_1 _09544_ (.A(_03366_),
    .B(_03375_),
    .C(_03609_),
    .D(_03401_),
    .Y(_03611_));
 sky130_fd_sc_hd__o211a_1 _09545_ (.A1(_03365_),
    .A2(_03582_),
    .B1(_03584_),
    .C1(_03406_),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_1 _09546_ (.A(_03606_),
    .B(_03611_),
    .Y(_03613_));
 sky130_fd_sc_hd__o21ai_2 _09547_ (.A1(_03613_),
    .A2(_03612_),
    .B1(_03600_),
    .Y(_03614_));
 sky130_fd_sc_hd__and4_2 _09548_ (.A(_03405_),
    .B(_03597_),
    .C(_03416_),
    .D(_03375_),
    .X(_03615_));
 sky130_fd_sc_hd__nand2_4 _09549_ (.A(_03424_),
    .B(_03597_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand4_1 _09550_ (.A(net98),
    .B(_03375_),
    .C(_03603_),
    .D(_03401_),
    .Y(_03618_));
 sky130_fd_sc_hd__a22oi_4 _09551_ (.A1(_03400_),
    .A2(_03389_),
    .B1(_03579_),
    .B2(_03578_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand4_1 _09552_ (.A(net98),
    .B(_03582_),
    .C(_03401_),
    .D(_03373_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_2 _09553_ (.A(_03618_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__o21ai_2 _09554_ (.A1(_03621_),
    .A2(_03619_),
    .B1(_03615_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand3_1 _09555_ (.A(_03592_),
    .B(_03614_),
    .C(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__o211ai_1 _09556_ (.A1(net114),
    .A2(_03086_),
    .B1(_03417_),
    .C1(net101),
    .Y(_03624_));
 sky130_fd_sc_hd__nand2_1 _09557_ (.A(_03388_),
    .B(_03434_),
    .Y(_03625_));
 sky130_fd_sc_hd__o21a_1 _09558_ (.A1(_03388_),
    .A2(_03443_),
    .B1(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__o21ai_2 _09559_ (.A1(_03388_),
    .A2(_03443_),
    .B1(_03625_),
    .Y(_03628_));
 sky130_fd_sc_hd__o211ai_1 _09560_ (.A1(_03085_),
    .A2(_03083_),
    .B1(_03416_),
    .C1(net101),
    .Y(_03629_));
 sky130_fd_sc_hd__o21ai_2 _09561_ (.A1(_03365_),
    .A2(_03626_),
    .B1(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__nand4_2 _09562_ (.A(net98),
    .B(_03628_),
    .C(_03401_),
    .D(_03373_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand4_2 _09563_ (.A(net98),
    .B(_03375_),
    .C(_03587_),
    .D(_03401_),
    .Y(_03632_));
 sky130_fd_sc_hd__o211ai_2 _09564_ (.A1(net114),
    .A2(_03086_),
    .B1(_03373_),
    .C1(net101),
    .Y(_03633_));
 sky130_fd_sc_hd__o21a_1 _09565_ (.A1(_03596_),
    .A2(_03365_),
    .B1(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__o21ai_4 _09566_ (.A1(_03596_),
    .A2(_03365_),
    .B1(_03633_),
    .Y(_03635_));
 sky130_fd_sc_hd__o221a_1 _09567_ (.A1(net98),
    .A2(_03375_),
    .B1(_03398_),
    .B2(_03404_),
    .C1(_03598_),
    .X(_03636_));
 sky130_fd_sc_hd__nand2_1 _09568_ (.A(_03631_),
    .B(_03632_),
    .Y(_03637_));
 sky130_fd_sc_hd__a21oi_4 _09569_ (.A1(_03634_),
    .A2(_03406_),
    .B1(_03637_),
    .Y(_03639_));
 sky130_fd_sc_hd__o211ai_4 _09570_ (.A1(_03405_),
    .A2(_03635_),
    .B1(_03632_),
    .C1(_03631_),
    .Y(_03640_));
 sky130_fd_sc_hd__nand4_4 _09571_ (.A(net98),
    .B(_03375_),
    .C(_03628_),
    .D(_03401_),
    .Y(_03641_));
 sky130_fd_sc_hd__o211ai_4 _09572_ (.A1(net98),
    .A2(_03399_),
    .B1(_03406_),
    .C1(_03421_),
    .Y(_03642_));
 sky130_fd_sc_hd__o211a_4 _09573_ (.A1(_03575_),
    .A2(_03635_),
    .B1(_03641_),
    .C1(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__o211ai_4 _09574_ (.A1(_03575_),
    .A2(_03635_),
    .B1(_03641_),
    .C1(_03642_),
    .Y(_03644_));
 sky130_fd_sc_hd__o221a_1 _09575_ (.A1(net114),
    .A2(_03086_),
    .B1(_03223_),
    .B2(_03361_),
    .C1(_03500_),
    .X(_03645_));
 sky130_fd_sc_hd__a31o_1 _09576_ (.A1(_03007_),
    .A2(_03366_),
    .A3(_03388_),
    .B1(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__and3_4 _09577_ (.A(_03644_),
    .B(_03424_),
    .C(_03598_),
    .X(_03647_));
 sky130_fd_sc_hd__nand2_8 _09578_ (.A(_03644_),
    .B(_03600_),
    .Y(_03648_));
 sky130_fd_sc_hd__and3_1 _09579_ (.A(_03600_),
    .B(_03639_),
    .C(_03644_),
    .X(_03650_));
 sky130_fd_sc_hd__nand3_4 _09580_ (.A(_03600_),
    .B(_03639_),
    .C(_03644_),
    .Y(_03651_));
 sky130_fd_sc_hd__a31oi_1 _09581_ (.A1(_03592_),
    .A2(_03614_),
    .A3(_03622_),
    .B1(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__a31o_1 _09582_ (.A1(_03592_),
    .A2(_03614_),
    .A3(_03622_),
    .B1(_03651_),
    .X(_03653_));
 sky130_fd_sc_hd__nand4_1 _09583_ (.A(net98),
    .B(_03587_),
    .C(_03401_),
    .D(_03373_),
    .Y(_03654_));
 sky130_fd_sc_hd__nand4_1 _09584_ (.A(net98),
    .B(_03375_),
    .C(_03577_),
    .D(_03401_),
    .Y(_03655_));
 sky130_fd_sc_hd__o211a_1 _09585_ (.A1(_03365_),
    .A2(_03628_),
    .B1(_03624_),
    .C1(_03406_),
    .X(_03656_));
 sky130_fd_sc_hd__nand2_2 _09586_ (.A(_03654_),
    .B(_03655_),
    .Y(_03657_));
 sky130_fd_sc_hd__a21oi_4 _09587_ (.A1(_03406_),
    .A2(_03630_),
    .B1(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__o21ai_1 _09588_ (.A1(_03657_),
    .A2(_03656_),
    .B1(_03425_),
    .Y(_03659_));
 sky130_fd_sc_hd__o21ai_2 _09589_ (.A1(_03621_),
    .A2(_03619_),
    .B1(_03600_),
    .Y(_03661_));
 sky130_fd_sc_hd__o21ai_2 _09590_ (.A1(_03590_),
    .A2(_03591_),
    .B1(_03615_),
    .Y(_03662_));
 sky130_fd_sc_hd__o211ai_4 _09591_ (.A1(_03424_),
    .A2(_03658_),
    .B1(_03661_),
    .C1(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__o21ai_1 _09592_ (.A1(_03601_),
    .A2(_03643_),
    .B1(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__and3_1 _09593_ (.A(_03640_),
    .B(_03424_),
    .C(_03598_),
    .X(_03665_));
 sky130_fd_sc_hd__or3_1 _09594_ (.A(_03425_),
    .B(_03597_),
    .C(_03639_),
    .X(_03666_));
 sky130_fd_sc_hd__o21a_4 _09595_ (.A1(_03637_),
    .A2(_03636_),
    .B1(_03644_),
    .X(_03667_));
 sky130_fd_sc_hd__and3_4 _09596_ (.A(_03640_),
    .B(_03644_),
    .C(_03600_),
    .X(_03668_));
 sky130_fd_sc_hd__nand4_4 _09597_ (.A(_03598_),
    .B(_03640_),
    .C(_03644_),
    .D(_03424_),
    .Y(_03669_));
 sky130_fd_sc_hd__o21ai_2 _09598_ (.A1(_03621_),
    .A2(_03619_),
    .B1(_03425_),
    .Y(_03670_));
 sky130_fd_sc_hd__o21ai_2 _09599_ (.A1(_03613_),
    .A2(_03612_),
    .B1(_03615_),
    .Y(_03672_));
 sky130_fd_sc_hd__a311o_1 _09600_ (.A1(net98),
    .A2(_03593_),
    .A3(_03595_),
    .B1(_03491_),
    .C1(_03425_),
    .X(_03673_));
 sky130_fd_sc_hd__o211ai_4 _09601_ (.A1(_03491_),
    .A2(_03601_),
    .B1(_03670_),
    .C1(_03672_),
    .Y(_03674_));
 sky130_fd_sc_hd__nand3_1 _09602_ (.A(_03674_),
    .B(_03667_),
    .C(_03600_),
    .Y(_03675_));
 sky130_fd_sc_hd__a221oi_2 _09603_ (.A1(_03648_),
    .A2(_03663_),
    .B1(_03668_),
    .B2(_03674_),
    .C1(_03652_),
    .Y(_03676_));
 sky130_fd_sc_hd__nand3_2 _09604_ (.A(_03653_),
    .B(_03664_),
    .C(_03675_),
    .Y(_03677_));
 sky130_fd_sc_hd__o21ai_4 _09605_ (.A1(_03591_),
    .A2(_03590_),
    .B1(_03600_),
    .Y(_03678_));
 sky130_fd_sc_hd__o21ai_2 _09606_ (.A1(_03657_),
    .A2(_03656_),
    .B1(_03615_),
    .Y(_03679_));
 sky130_fd_sc_hd__o21ai_2 _09607_ (.A1(_03617_),
    .A2(_03658_),
    .B1(_03678_),
    .Y(_03680_));
 sky130_fd_sc_hd__a211o_2 _09608_ (.A1(_03678_),
    .A2(_03679_),
    .B1(_03640_),
    .C1(_03648_),
    .X(_03681_));
 sky130_fd_sc_hd__o21ai_1 _09609_ (.A1(_03657_),
    .A2(_03656_),
    .B1(_03600_),
    .Y(_03683_));
 sky130_fd_sc_hd__o221ai_4 _09610_ (.A1(_03424_),
    .A2(_03643_),
    .B1(_03639_),
    .B2(_03617_),
    .C1(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__o21ai_2 _09611_ (.A1(_03601_),
    .A2(_03643_),
    .B1(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__a31o_1 _09612_ (.A1(_03659_),
    .A2(_03661_),
    .A3(_03662_),
    .B1(_03669_),
    .X(_03686_));
 sky130_fd_sc_hd__a22oi_4 _09613_ (.A1(_03663_),
    .A2(_03668_),
    .B1(_03684_),
    .B2(_03648_),
    .Y(_03687_));
 sky130_fd_sc_hd__o31a_1 _09614_ (.A1(_03373_),
    .A2(_03406_),
    .A3(_03417_),
    .B1(_03640_),
    .X(_03688_));
 sky130_fd_sc_hd__o211a_4 _09615_ (.A1(_03424_),
    .A2(_03639_),
    .B1(_03678_),
    .C1(_03679_),
    .X(_03689_));
 sky130_fd_sc_hd__o211ai_4 _09616_ (.A1(_03424_),
    .A2(_03639_),
    .B1(_03678_),
    .C1(_03679_),
    .Y(_03690_));
 sky130_fd_sc_hd__o311a_2 _09617_ (.A1(_03640_),
    .A2(_03648_),
    .A3(_03689_),
    .B1(_03686_),
    .C1(_03685_),
    .X(_03691_));
 sky130_fd_sc_hd__o211ai_4 _09618_ (.A1(_03651_),
    .A2(_03689_),
    .B1(_03686_),
    .C1(_03685_),
    .Y(_03692_));
 sky130_fd_sc_hd__a22oi_2 _09619_ (.A1(_03641_),
    .A2(_03424_),
    .B1(_03423_),
    .B2(_03599_),
    .Y(_03694_));
 sky130_fd_sc_hd__nand4_4 _09620_ (.A(_03644_),
    .B(_03658_),
    .C(_03424_),
    .D(_03600_),
    .Y(_03695_));
 sky130_fd_sc_hd__o22a_1 _09621_ (.A1(_03665_),
    .A2(_03694_),
    .B1(_03684_),
    .B2(_03648_),
    .X(_03696_));
 sky130_fd_sc_hd__o21ai_2 _09622_ (.A1(_03665_),
    .A2(_03694_),
    .B1(_03695_),
    .Y(_03697_));
 sky130_fd_sc_hd__and3_4 _09623_ (.A(_03695_),
    .B(_03667_),
    .C(_03600_),
    .X(_03698_));
 sky130_fd_sc_hd__nand3_4 _09624_ (.A(_03600_),
    .B(_03667_),
    .C(_03695_),
    .Y(_03699_));
 sky130_fd_sc_hd__and3_4 _09625_ (.A(_03668_),
    .B(_03690_),
    .C(_03695_),
    .X(_03700_));
 sky130_fd_sc_hd__nand4_4 _09626_ (.A(_03690_),
    .B(_03695_),
    .C(_03600_),
    .D(_03667_),
    .Y(_03701_));
 sky130_fd_sc_hd__a31o_1 _09627_ (.A1(_03659_),
    .A2(_03661_),
    .A3(_03662_),
    .B1(_03651_),
    .X(_03702_));
 sky130_fd_sc_hd__a31o_1 _09628_ (.A1(_03592_),
    .A2(_03614_),
    .A3(_03622_),
    .B1(_03669_),
    .X(_03703_));
 sky130_fd_sc_hd__o211ai_4 _09629_ (.A1(_03647_),
    .A2(_03689_),
    .B1(_03702_),
    .C1(_03703_),
    .Y(_03705_));
 sky130_fd_sc_hd__a21oi_4 _09630_ (.A1(_03687_),
    .A2(_03681_),
    .B1(_03701_),
    .Y(_03706_));
 sky130_fd_sc_hd__a21o_2 _09631_ (.A1(_03687_),
    .A2(_03681_),
    .B1(_03701_),
    .X(_03707_));
 sky130_fd_sc_hd__a31o_1 _09632_ (.A1(_03653_),
    .A2(_03664_),
    .A3(_03675_),
    .B1(_03701_),
    .X(_03708_));
 sky130_fd_sc_hd__a211o_1 _09633_ (.A1(_03681_),
    .A2(_03687_),
    .B1(_03701_),
    .C1(_03676_),
    .X(_03709_));
 sky130_fd_sc_hd__o21ai_1 _09634_ (.A1(_03669_),
    .A2(_03689_),
    .B1(_03697_),
    .Y(_03710_));
 sky130_fd_sc_hd__o211ai_2 _09635_ (.A1(_03692_),
    .A2(_03699_),
    .B1(_03701_),
    .C1(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__and3_4 _09636_ (.A(_03692_),
    .B(_03705_),
    .C(_03700_),
    .X(_03712_));
 sky130_fd_sc_hd__nand4_4 _09637_ (.A(_03690_),
    .B(_03692_),
    .C(_03705_),
    .D(_03698_),
    .Y(_03713_));
 sky130_fd_sc_hd__a311oi_2 _09638_ (.A1(_03670_),
    .A2(_03672_),
    .A3(_03673_),
    .B1(_03648_),
    .C1(_03640_),
    .Y(_03714_));
 sky130_fd_sc_hd__a31o_1 _09639_ (.A1(_03670_),
    .A2(_03672_),
    .A3(_03673_),
    .B1(_03651_),
    .X(_03716_));
 sky130_fd_sc_hd__nand2_1 _09640_ (.A(net100),
    .B(_03483_),
    .Y(_03717_));
 sky130_fd_sc_hd__a211o_1 _09641_ (.A1(_03380_),
    .A2(_03379_),
    .B1(_03491_),
    .C1(_03387_),
    .X(_03718_));
 sky130_fd_sc_hd__o21ai_1 _09642_ (.A1(_03388_),
    .A2(_03532_),
    .B1(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__o21ai_4 _09643_ (.A1(net100),
    .A2(_03719_),
    .B1(_03717_),
    .Y(_03720_));
 sky130_fd_sc_hd__o21ai_1 _09644_ (.A1(_03601_),
    .A2(_03643_),
    .B1(_03623_),
    .Y(_03721_));
 sky130_fd_sc_hd__o2bb2ai_1 _09645_ (.A1_N(_03623_),
    .A2_N(_03648_),
    .B1(_03669_),
    .B2(_03720_),
    .Y(_03722_));
 sky130_fd_sc_hd__o211ai_1 _09646_ (.A1(_03669_),
    .A2(_03720_),
    .B1(_03721_),
    .C1(_03716_),
    .Y(_03723_));
 sky130_fd_sc_hd__o22ai_1 _09647_ (.A1(_03680_),
    .A2(_03688_),
    .B1(_03714_),
    .B2(_03722_),
    .Y(_03724_));
 sky130_fd_sc_hd__a21oi_2 _09648_ (.A1(_03724_),
    .A2(_03698_),
    .B1(_03691_),
    .Y(_03725_));
 sky130_fd_sc_hd__and3_1 _09649_ (.A(_03687_),
    .B(_03700_),
    .C(_03681_),
    .X(_03727_));
 sky130_fd_sc_hd__nand4b_2 _09650_ (.A_N(_03701_),
    .B(_03686_),
    .C(_03685_),
    .D(_03681_),
    .Y(_03728_));
 sky130_fd_sc_hd__nor2_1 _09651_ (.A(_03690_),
    .B(_03699_),
    .Y(_03729_));
 sky130_fd_sc_hd__a211o_1 _09652_ (.A1(_03425_),
    .A2(_03640_),
    .B1(_03680_),
    .C1(_03699_),
    .X(_03730_));
 sky130_fd_sc_hd__o2bb2ai_2 _09653_ (.A1_N(_03729_),
    .A2_N(_03705_),
    .B1(_03676_),
    .B2(_03728_),
    .Y(_03731_));
 sky130_fd_sc_hd__nor2_4 _09654_ (.A(_03731_),
    .B(_03725_),
    .Y(_03732_));
 sky130_fd_sc_hd__or2_2 _09655_ (.A(_03731_),
    .B(_03725_),
    .X(_03733_));
 sky130_fd_sc_hd__nor2_4 _09656_ (.A(_03713_),
    .B(_03732_),
    .Y(_03734_));
 sky130_fd_sc_hd__o2111ai_4 _09657_ (.A1(_03680_),
    .A2(_03688_),
    .B1(_03705_),
    .C1(_03698_),
    .D1(_03691_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand3_4 _09658_ (.A(_03709_),
    .B(_03711_),
    .C(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__nor3b_4 _09659_ (.A(_03691_),
    .B(_03708_),
    .C_N(_03705_),
    .Y(_03738_));
 sky130_fd_sc_hd__nand3_4 _09660_ (.A(_03706_),
    .B(_03705_),
    .C(_03677_),
    .Y(_03739_));
 sky130_fd_sc_hd__nor2_1 _09661_ (.A(_03387_),
    .B(_03548_),
    .Y(_03740_));
 sky130_fd_sc_hd__a2bb2o_1 _09662_ (.A1_N(_03388_),
    .A2_N(_03521_),
    .B1(_03381_),
    .B2(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__a21oi_1 _09663_ (.A1(_03087_),
    .A2(_03364_),
    .B1(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__a31o_1 _09664_ (.A1(_03087_),
    .A2(_03364_),
    .A3(_03507_),
    .B1(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__nand4_1 _09665_ (.A(_03401_),
    .B(_03741_),
    .C(_03366_),
    .D(_03375_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_1 _09666_ (.A(net100),
    .B(_03513_),
    .Y(_03745_));
 sky130_fd_sc_hd__nand2_1 _09667_ (.A(_03388_),
    .B(_03507_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21boi_1 _09668_ (.A1(_03389_),
    .A2(_03548_),
    .B1_N(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__o21ai_4 _09669_ (.A1(net100),
    .A2(_03747_),
    .B1(_03745_),
    .Y(_03749_));
 sky130_fd_sc_hd__a211o_1 _09670_ (.A1(_03380_),
    .A2(_03379_),
    .B1(_03513_),
    .C1(_03387_),
    .X(_03750_));
 sky130_fd_sc_hd__o21ai_2 _09671_ (.A1(_03388_),
    .A2(_03507_),
    .B1(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__nand2_1 _09672_ (.A(net100),
    .B(_03541_),
    .Y(_03752_));
 sky130_fd_sc_hd__o21ai_4 _09673_ (.A1(net100),
    .A2(_03751_),
    .B1(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__o221a_2 _09674_ (.A1(_03575_),
    .A2(_03749_),
    .B1(_03753_),
    .B2(_03405_),
    .C1(_03744_),
    .X(_03754_));
 sky130_fd_sc_hd__o221ai_1 _09675_ (.A1(_03575_),
    .A2(_03749_),
    .B1(_03405_),
    .B2(_03753_),
    .C1(_03744_),
    .Y(_03755_));
 sky130_fd_sc_hd__and3_1 _09676_ (.A(_03381_),
    .B(_03386_),
    .C(_03521_),
    .X(_03756_));
 sky130_fd_sc_hd__a21oi_1 _09677_ (.A1(_03389_),
    .A2(_03500_),
    .B1(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__a221o_1 _09678_ (.A1(_03500_),
    .A2(_03389_),
    .B1(_03364_),
    .B2(_03087_),
    .C1(_03756_),
    .X(_03758_));
 sky130_fd_sc_hd__nand4_1 _09679_ (.A(_03401_),
    .B(_03757_),
    .C(_03366_),
    .D(_03375_),
    .Y(_03760_));
 sky130_fd_sc_hd__o21ai_1 _09680_ (.A1(net100),
    .A2(_03741_),
    .B1(_03574_),
    .Y(_03761_));
 sky130_fd_sc_hd__o211ai_2 _09681_ (.A1(_03405_),
    .A2(_03749_),
    .B1(_03760_),
    .C1(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__nand4_2 _09682_ (.A(_03373_),
    .B(_03751_),
    .C(_03401_),
    .D(_03366_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand2_1 _09683_ (.A(net100),
    .B(_03558_),
    .Y(_03764_));
 sky130_fd_sc_hd__a21o_1 _09684_ (.A1(_03381_),
    .A2(_03386_),
    .B1(_03513_),
    .X(_03765_));
 sky130_fd_sc_hd__o21ai_2 _09685_ (.A1(_03389_),
    .A2(_03541_),
    .B1(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__o21a_4 _09686_ (.A1(net100),
    .A2(_03766_),
    .B1(_03764_),
    .X(_03767_));
 sky130_fd_sc_hd__o21ai_4 _09687_ (.A1(net100),
    .A2(_03766_),
    .B1(_03764_),
    .Y(_03768_));
 sky130_fd_sc_hd__o221ai_4 _09688_ (.A1(_03409_),
    .A2(_03749_),
    .B1(_03405_),
    .B2(_03768_),
    .C1(_03763_),
    .Y(_03769_));
 sky130_fd_sc_hd__a22oi_1 _09689_ (.A1(_03762_),
    .A2(_03600_),
    .B1(_03425_),
    .B2(_03769_),
    .Y(_03771_));
 sky130_fd_sc_hd__o21ai_1 _09690_ (.A1(_03617_),
    .A2(_03754_),
    .B1(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__or4b_1 _09691_ (.A(net100),
    .B(_03375_),
    .C(_03402_),
    .D_N(_03757_),
    .X(_03773_));
 sky130_fd_sc_hd__mux2_1 _09692_ (.A0(_03007_),
    .A1(_03500_),
    .S(_03388_),
    .X(_03774_));
 sky130_fd_sc_hd__mux2_1 _09693_ (.A0(_03774_),
    .A1(_03521_),
    .S(net100),
    .X(_03775_));
 sky130_fd_sc_hd__o221ai_4 _09694_ (.A1(_03743_),
    .A2(_03405_),
    .B1(_03409_),
    .B2(_03775_),
    .C1(_03773_),
    .Y(_03776_));
 sky130_fd_sc_hd__a22oi_1 _09695_ (.A1(_03615_),
    .A2(_03762_),
    .B1(_03776_),
    .B2(_03600_),
    .Y(_03777_));
 sky130_fd_sc_hd__o21ai_1 _09696_ (.A1(_03424_),
    .A2(_03754_),
    .B1(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__or4_1 _09697_ (.A(_03425_),
    .B(_03597_),
    .C(_03643_),
    .D(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__o21ai_1 _09698_ (.A1(_03647_),
    .A2(_03772_),
    .B1(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__o31a_1 _09699_ (.A1(_03601_),
    .A2(_03639_),
    .A3(_03643_),
    .B1(_03780_),
    .X(_03782_));
 sky130_fd_sc_hd__nor2_4 _09700_ (.A(_03739_),
    .B(_03732_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _09701_ (.A(_03733_),
    .B(_03738_),
    .Y(_03784_));
 sky130_fd_sc_hd__o21ai_1 _09702_ (.A1(_03714_),
    .A2(_03722_),
    .B1(_03729_),
    .Y(_03785_));
 sky130_fd_sc_hd__o21ai_1 _09703_ (.A1(_03669_),
    .A2(_03697_),
    .B1(_03677_),
    .Y(_03786_));
 sky130_fd_sc_hd__a21oi_1 _09704_ (.A1(_03381_),
    .A2(_03386_),
    .B1(_03491_),
    .Y(_03787_));
 sky130_fd_sc_hd__a221o_1 _09705_ (.A1(_03399_),
    .A2(_03403_),
    .B1(_03458_),
    .B2(_03365_),
    .C1(_03604_),
    .X(_03788_));
 sky130_fd_sc_hd__or3_1 _09706_ (.A(_03607_),
    .B(_03610_),
    .C(_03575_),
    .X(_03789_));
 sky130_fd_sc_hd__o311a_1 _09707_ (.A1(_03373_),
    .A2(_03406_),
    .A3(_03491_),
    .B1(_03788_),
    .C1(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__o211ai_1 _09708_ (.A1(net114),
    .A2(_03086_),
    .B1(_03476_),
    .C1(_03364_),
    .Y(_03791_));
 sky130_fd_sc_hd__o2bb2ai_1 _09709_ (.A1_N(_03087_),
    .A2_N(_03364_),
    .B1(_03389_),
    .B2(_03483_),
    .Y(_03793_));
 sky130_fd_sc_hd__a22oi_1 _09710_ (.A1(_03787_),
    .A2(_03366_),
    .B1(_03793_),
    .B2(_03791_),
    .Y(_03794_));
 sky130_fd_sc_hd__a31o_1 _09711_ (.A1(_03366_),
    .A2(_03389_),
    .A3(_03399_),
    .B1(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__nand2_1 _09712_ (.A(net100),
    .B(_03491_),
    .Y(_03796_));
 sky130_fd_sc_hd__a21o_1 _09713_ (.A1(_03381_),
    .A2(_03386_),
    .B1(_03558_),
    .X(_03797_));
 sky130_fd_sc_hd__o21ai_1 _09714_ (.A1(_03389_),
    .A2(_03532_),
    .B1(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__o21ai_2 _09715_ (.A1(net100),
    .A2(_03798_),
    .B1(_03796_),
    .Y(_03799_));
 sky130_fd_sc_hd__o221ai_4 _09716_ (.A1(_03575_),
    .A2(_03720_),
    .B1(_03799_),
    .B2(_03409_),
    .C1(_03795_),
    .Y(_03800_));
 sky130_fd_sc_hd__a2bb2oi_1 _09717_ (.A1_N(_03617_),
    .A2_N(_03720_),
    .B1(_03600_),
    .B2(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__o21ai_2 _09718_ (.A1(_03424_),
    .A2(_03790_),
    .B1(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _09719_ (.A(_03700_),
    .B(_03802_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand3_2 _09720_ (.A(_03785_),
    .B(_03786_),
    .C(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__a22o_1 _09721_ (.A1(_03677_),
    .A2(_03729_),
    .B1(_03705_),
    .B2(_03699_),
    .X(_03806_));
 sky130_fd_sc_hd__and4_1 _09722_ (.A(_03687_),
    .B(_03723_),
    .C(_03700_),
    .D(_03681_),
    .X(_03807_));
 sky130_fd_sc_hd__a211oi_4 _09723_ (.A1(_03805_),
    .A2(_03706_),
    .B1(_03806_),
    .C1(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__a211o_4 _09724_ (.A1(_03805_),
    .A2(_03706_),
    .B1(_03807_),
    .C1(_03806_),
    .X(_03809_));
 sky130_fd_sc_hd__and3_1 _09725_ (.A(_03733_),
    .B(_03809_),
    .C(_03738_),
    .X(_03810_));
 sky130_fd_sc_hd__nand2_2 _09726_ (.A(_03783_),
    .B(_03809_),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2_1 _09727_ (.A(net100),
    .B(_03532_),
    .Y(_03812_));
 sky130_fd_sc_hd__o21ai_1 _09728_ (.A1(_03389_),
    .A2(_03558_),
    .B1(_03366_),
    .Y(_03813_));
 sky130_fd_sc_hd__a2bb2oi_4 _09729_ (.A1_N(_03541_),
    .A2_N(_03404_),
    .B1(_03813_),
    .B2(_03812_),
    .Y(_03815_));
 sky130_fd_sc_hd__nand2_1 _09730_ (.A(_03712_),
    .B(_03808_),
    .Y(_03816_));
 sky130_fd_sc_hd__a21oi_1 _09731_ (.A1(_03736_),
    .A2(_03816_),
    .B1(_03734_),
    .Y(_03817_));
 sky130_fd_sc_hd__and3_1 _09732_ (.A(_03698_),
    .B(_03815_),
    .C(_03690_),
    .X(_03818_));
 sky130_fd_sc_hd__and3_1 _09733_ (.A(_03818_),
    .B(_03705_),
    .C(_03692_),
    .X(_03819_));
 sky130_fd_sc_hd__nand4_2 _09734_ (.A(_03692_),
    .B(_03705_),
    .C(_03815_),
    .D(_03700_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21oi_2 _09735_ (.A1(_03783_),
    .A2(_03819_),
    .B1(_03817_),
    .Y(_03821_));
 sky130_fd_sc_hd__and3_1 _09736_ (.A(_03783_),
    .B(_03809_),
    .C(_03820_),
    .X(_03822_));
 sky130_fd_sc_hd__nand3_4 _09737_ (.A(_03783_),
    .B(_03809_),
    .C(_03820_),
    .Y(_03823_));
 sky130_fd_sc_hd__or4_1 _09738_ (.A(_03732_),
    .B(_03739_),
    .C(_03767_),
    .D(_03809_),
    .X(_03824_));
 sky130_fd_sc_hd__and4_1 _09739_ (.A(_03733_),
    .B(_03736_),
    .C(_03753_),
    .D(_03712_),
    .X(_03826_));
 sky130_fd_sc_hd__nand4_1 _09740_ (.A(_03733_),
    .B(_03736_),
    .C(_03753_),
    .D(_03712_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_4 _09741_ (.A(_03826_),
    .B(_03809_),
    .Y(_03828_));
 sky130_fd_sc_hd__nand2_1 _09742_ (.A(_03738_),
    .B(_03753_),
    .Y(_03829_));
 sky130_fd_sc_hd__o211a_1 _09743_ (.A1(_03733_),
    .A2(_03712_),
    .B1(_03828_),
    .C1(_03824_),
    .X(_03830_));
 sky130_fd_sc_hd__o2bb2a_1 _09744_ (.A1_N(_03815_),
    .A2_N(_03738_),
    .B1(_03736_),
    .B2(_03816_),
    .X(_03831_));
 sky130_fd_sc_hd__o211a_1 _09745_ (.A1(_03783_),
    .A2(_03831_),
    .B1(_03823_),
    .C1(_03830_),
    .X(_03832_));
 sky130_fd_sc_hd__o211a_2 _09746_ (.A1(_03784_),
    .A2(_03820_),
    .B1(_03810_),
    .C1(_03767_),
    .X(_03833_));
 sky130_fd_sc_hd__a211o_2 _09747_ (.A1(_03783_),
    .A2(_03819_),
    .B1(_03811_),
    .C1(_03768_),
    .X(_03834_));
 sky130_fd_sc_hd__and3_2 _09748_ (.A(_03828_),
    .B(_03822_),
    .C(_03767_),
    .X(_03835_));
 sky130_fd_sc_hd__o21ai_2 _09749_ (.A1(_03808_),
    .A2(_03827_),
    .B1(_03833_),
    .Y(_03837_));
 sky130_fd_sc_hd__nand2_1 _09750_ (.A(_03772_),
    .B(_03647_),
    .Y(_03838_));
 sky130_fd_sc_hd__a2bb2o_1 _09751_ (.A1_N(_03409_),
    .A2_N(_03753_),
    .B1(_03766_),
    .B2(_03574_),
    .X(_03839_));
 sky130_fd_sc_hd__a2bb2o_1 _09752_ (.A1_N(_03405_),
    .A2_N(_03815_),
    .B1(_03416_),
    .B2(_03408_),
    .X(_03840_));
 sky130_fd_sc_hd__o22ai_4 _09753_ (.A1(_03425_),
    .A2(_03769_),
    .B1(_03839_),
    .B2(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__inv_2 _09754_ (.A(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__or4_2 _09755_ (.A(_03417_),
    .B(_03597_),
    .C(_03409_),
    .D(_03630_),
    .X(_03843_));
 sky130_fd_sc_hd__o221a_2 _09756_ (.A1(_03600_),
    .A2(_03841_),
    .B1(_03843_),
    .B2(_03754_),
    .C1(_03838_),
    .X(_03844_));
 sky130_fd_sc_hd__o221ai_4 _09757_ (.A1(_03600_),
    .A2(_03841_),
    .B1(_03843_),
    .B2(_03754_),
    .C1(_03838_),
    .Y(_03845_));
 sky130_fd_sc_hd__a32o_1 _09758_ (.A1(_03768_),
    .A2(_03822_),
    .A3(_03842_),
    .B1(_03835_),
    .B2(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__nor2_1 _09759_ (.A(_03832_),
    .B(_03846_),
    .Y(_03848_));
 sky130_fd_sc_hd__nor2_1 _09760_ (.A(_03828_),
    .B(_03834_),
    .Y(_03849_));
 sky130_fd_sc_hd__o31a_2 _09761_ (.A1(_03768_),
    .A2(_03823_),
    .A3(_03828_),
    .B1(_03848_),
    .X(_03850_));
 sky130_fd_sc_hd__o21a_1 _09762_ (.A1(_03713_),
    .A2(_03767_),
    .B1(_03736_),
    .X(_03851_));
 sky130_fd_sc_hd__a21oi_1 _09763_ (.A1(_03712_),
    .A2(_03815_),
    .B1(_03736_),
    .Y(_03852_));
 sky130_fd_sc_hd__o22a_1 _09764_ (.A1(_03809_),
    .A2(_03712_),
    .B1(_03852_),
    .B2(_03851_),
    .X(_03853_));
 sky130_fd_sc_hd__a31o_1 _09765_ (.A1(_03712_),
    .A2(_03733_),
    .A3(_03736_),
    .B1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__o211ai_1 _09766_ (.A1(_03784_),
    .A2(_03808_),
    .B1(_03827_),
    .C1(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand4_1 _09767_ (.A(_03424_),
    .B(_03643_),
    .C(_03769_),
    .D(_03598_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand4_1 _09768_ (.A(_03598_),
    .B(_03644_),
    .C(_03755_),
    .D(_03424_),
    .Y(_03857_));
 sky130_fd_sc_hd__a22oi_1 _09769_ (.A1(_03815_),
    .A2(_03574_),
    .B1(_03406_),
    .B2(_03799_),
    .Y(_03859_));
 sky130_fd_sc_hd__o211ai_1 _09770_ (.A1(_03409_),
    .A2(_03767_),
    .B1(_03425_),
    .C1(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__o2111a_1 _09771_ (.A1(_03617_),
    .A2(_03753_),
    .B1(_03856_),
    .C1(_03857_),
    .D1(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__nand4_1 _09772_ (.A(_03373_),
    .B(_03798_),
    .C(_03401_),
    .D(net98),
    .Y(_03862_));
 sky130_fd_sc_hd__o221a_1 _09773_ (.A1(_03409_),
    .A2(_03815_),
    .B1(_03720_),
    .B2(_03405_),
    .C1(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__o22ai_1 _09774_ (.A1(_03601_),
    .A2(_03753_),
    .B1(_03863_),
    .B2(_03424_),
    .Y(_03864_));
 sky130_fd_sc_hd__a31o_1 _09775_ (.A1(_03424_),
    .A2(_03597_),
    .A3(_03767_),
    .B1(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__o22ai_1 _09776_ (.A1(_03651_),
    .A2(_03841_),
    .B1(_03669_),
    .B2(_03861_),
    .Y(_03866_));
 sky130_fd_sc_hd__a21oi_1 _09777_ (.A1(_03648_),
    .A2(_03865_),
    .B1(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__nand4_1 _09778_ (.A(_03647_),
    .B(_03866_),
    .C(_03696_),
    .D(_03640_),
    .Y(_03868_));
 sky130_fd_sc_hd__o21ai_1 _09779_ (.A1(_03409_),
    .A2(_03417_),
    .B1(_03800_),
    .Y(_03870_));
 sky130_fd_sc_hd__o31a_1 _09780_ (.A1(_03409_),
    .A2(_03423_),
    .A3(_03815_),
    .B1(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__o32a_1 _09781_ (.A1(_03601_),
    .A2(_03643_),
    .A3(_03753_),
    .B1(_03768_),
    .B2(_03843_),
    .X(_03872_));
 sky130_fd_sc_hd__o21ai_1 _09782_ (.A1(_03600_),
    .A2(_03871_),
    .B1(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__nor3_1 _09783_ (.A(_03695_),
    .B(_03643_),
    .C(_03666_),
    .Y(_03874_));
 sky130_fd_sc_hd__or3_1 _09784_ (.A(_03695_),
    .B(_03643_),
    .C(_03666_),
    .X(_03875_));
 sky130_fd_sc_hd__a22oi_2 _09785_ (.A1(_03842_),
    .A2(_03874_),
    .B1(_03873_),
    .B2(_03669_),
    .Y(_03876_));
 sky130_fd_sc_hd__o21ai_2 _09786_ (.A1(_03699_),
    .A2(_03867_),
    .B1(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__a2bb2o_1 _09787_ (.A1_N(_03612_),
    .A2_N(_03613_),
    .B1(_03408_),
    .B2(_03416_),
    .X(_03878_));
 sky130_fd_sc_hd__o221a_1 _09788_ (.A1(_03491_),
    .A2(_03617_),
    .B1(_03720_),
    .B2(_03601_),
    .C1(_03648_),
    .X(_03879_));
 sky130_fd_sc_hd__a21oi_1 _09789_ (.A1(_03879_),
    .A2(_03878_),
    .B1(_03668_),
    .Y(_03881_));
 sky130_fd_sc_hd__o21ai_1 _09790_ (.A1(_03648_),
    .A2(_03802_),
    .B1(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__o311a_1 _09791_ (.A1(_03639_),
    .A2(_03648_),
    .A3(_03815_),
    .B1(_03882_),
    .C1(_03699_),
    .X(_03883_));
 sky130_fd_sc_hd__a211o_1 _09792_ (.A1(_03768_),
    .A2(_03698_),
    .B1(_03700_),
    .C1(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__or4b_1 _09793_ (.A(_03639_),
    .B(_03648_),
    .C(_03697_),
    .D_N(_03753_),
    .X(_03885_));
 sky130_fd_sc_hd__o2bb2a_1 _09794_ (.A1_N(_03650_),
    .A2_N(_03815_),
    .B1(_03647_),
    .B2(_03802_),
    .X(_03886_));
 sky130_fd_sc_hd__o211a_1 _09795_ (.A1(_03767_),
    .A2(_03875_),
    .B1(_03886_),
    .C1(_03885_),
    .X(_03887_));
 sky130_fd_sc_hd__o22a_1 _09796_ (.A1(_03707_),
    .A2(_03877_),
    .B1(_03887_),
    .B2(_03700_),
    .X(_03888_));
 sky130_fd_sc_hd__o21ai_1 _09797_ (.A1(_03707_),
    .A2(_03877_),
    .B1(_03712_),
    .Y(_03889_));
 sky130_fd_sc_hd__o32a_1 _09798_ (.A1(_03705_),
    .A2(_03707_),
    .A3(_03841_),
    .B1(_03753_),
    .B2(_03728_),
    .X(_03890_));
 sky130_fd_sc_hd__nand3_1 _09799_ (.A(_03889_),
    .B(_03890_),
    .C(_03884_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _09800_ (.A(_03732_),
    .B(_03738_),
    .Y(_03893_));
 sky130_fd_sc_hd__o2bb2a_1 _09801_ (.A1_N(_03700_),
    .A2_N(_03815_),
    .B1(_03802_),
    .B2(_03730_),
    .X(_03894_));
 sky130_fd_sc_hd__o221ai_1 _09802_ (.A1(_03691_),
    .A2(_03701_),
    .B1(_03723_),
    .B2(_03698_),
    .C1(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__o211a_1 _09803_ (.A1(_03707_),
    .A2(_03768_),
    .B1(_03895_),
    .C1(_03713_),
    .X(_03896_));
 sky130_fd_sc_hd__a31o_1 _09804_ (.A1(_03705_),
    .A2(_03706_),
    .A3(_03753_),
    .B1(_03738_),
    .X(_03897_));
 sky130_fd_sc_hd__o22ai_1 _09805_ (.A1(_03841_),
    .A2(_03893_),
    .B1(_03897_),
    .B2(_03896_),
    .Y(_03898_));
 sky130_fd_sc_hd__a31o_1 _09806_ (.A1(_03734_),
    .A2(_03736_),
    .A3(_03892_),
    .B1(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__nand2_1 _09807_ (.A(_03899_),
    .B(_03822_),
    .Y(_03900_));
 sky130_fd_sc_hd__nor2_1 _09808_ (.A(_03811_),
    .B(_03821_),
    .Y(_03901_));
 sky130_fd_sc_hd__o311a_4 _09809_ (.A1(_03811_),
    .A2(_03821_),
    .A3(_03841_),
    .B1(_03855_),
    .C1(_03900_),
    .X(_03903_));
 sky130_fd_sc_hd__o22a_1 _09810_ (.A1(_03844_),
    .A2(_03730_),
    .B1(_03698_),
    .B2(_03867_),
    .X(_03904_));
 sky130_fd_sc_hd__nand4_1 _09811_ (.A(_03647_),
    .B(_03778_),
    .C(_03696_),
    .D(_03640_),
    .Y(_03905_));
 sky130_fd_sc_hd__o221a_1 _09812_ (.A1(_03668_),
    .A2(_03861_),
    .B1(_03875_),
    .B2(_03844_),
    .C1(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__a21oi_1 _09813_ (.A1(_03904_),
    .A2(_03906_),
    .B1(_03707_),
    .Y(_03907_));
 sky130_fd_sc_hd__a221oi_2 _09814_ (.A1(_03727_),
    .A2(_03845_),
    .B1(_03877_),
    .B2(_03701_),
    .C1(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__and2_1 _09815_ (.A(_03908_),
    .B(_03713_),
    .X(_03909_));
 sky130_fd_sc_hd__and3_1 _09816_ (.A(_03833_),
    .B(_03842_),
    .C(_03828_),
    .X(_03910_));
 sky130_fd_sc_hd__or3b_2 _09817_ (.A(_03834_),
    .B(_03841_),
    .C_N(_03828_),
    .X(_03911_));
 sky130_fd_sc_hd__or3_2 _09818_ (.A(_03837_),
    .B(_03841_),
    .C(_03903_),
    .X(_03912_));
 sky130_fd_sc_hd__o31a_1 _09819_ (.A1(_03828_),
    .A2(_03834_),
    .A3(_03903_),
    .B1(_03848_),
    .X(_03914_));
 sky130_fd_sc_hd__nor2_4 _09820_ (.A(_03912_),
    .B(_03850_),
    .Y(_03915_));
 sky130_fd_sc_hd__or4_4 _09821_ (.A(_03837_),
    .B(_03903_),
    .C(_03841_),
    .D(_03850_),
    .X(_03916_));
 sky130_fd_sc_hd__and3_1 _09822_ (.A(_03868_),
    .B(_03876_),
    .C(_03727_),
    .X(_03917_));
 sky130_fd_sc_hd__o211a_1 _09823_ (.A1(_03705_),
    .A2(_03844_),
    .B1(_03692_),
    .C1(_03700_),
    .X(_03918_));
 sky130_fd_sc_hd__o32ai_1 _09824_ (.A1(_03405_),
    .A2(_03607_),
    .A3(_03610_),
    .B1(_03720_),
    .B2(_03409_),
    .Y(_03919_));
 sky130_fd_sc_hd__o21bai_1 _09825_ (.A1(_03491_),
    .A2(_03575_),
    .B1_N(_03919_),
    .Y(_03920_));
 sky130_fd_sc_hd__a2bb2o_1 _09826_ (.A1_N(_03601_),
    .A2_N(_03815_),
    .B1(_03920_),
    .B2(_03425_),
    .X(_03921_));
 sky130_fd_sc_hd__a211o_1 _09827_ (.A1(_03615_),
    .A2(_03800_),
    .B1(_03647_),
    .C1(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__or4b_1 _09828_ (.A(_03643_),
    .B(_03666_),
    .C(_03695_),
    .D_N(_03753_),
    .X(_03923_));
 sky130_fd_sc_hd__o221a_1 _09829_ (.A1(_03651_),
    .A2(_03767_),
    .B1(_03842_),
    .B2(_03699_),
    .C1(_03922_),
    .X(_03925_));
 sky130_fd_sc_hd__a21oi_1 _09830_ (.A1(_03925_),
    .A2(_03923_),
    .B1(_03700_),
    .Y(_03926_));
 sky130_fd_sc_hd__or3_1 _09831_ (.A(_03917_),
    .B(_03918_),
    .C(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__o21ai_2 _09832_ (.A1(_03713_),
    .A2(_03908_),
    .B1(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__a21oi_1 _09833_ (.A1(_03705_),
    .A2(_03706_),
    .B1(_03888_),
    .Y(_03929_));
 sky130_fd_sc_hd__a221o_1 _09834_ (.A1(_03727_),
    .A2(_03841_),
    .B1(_03844_),
    .B2(_03712_),
    .C1(_03738_),
    .X(_03930_));
 sky130_fd_sc_hd__o2bb2a_1 _09835_ (.A1_N(_03738_),
    .A2_N(_03928_),
    .B1(_03930_),
    .B2(_03929_),
    .X(_03931_));
 sky130_fd_sc_hd__a31o_1 _09836_ (.A1(_03712_),
    .A2(_03808_),
    .A3(_03845_),
    .B1(_03784_),
    .X(_03932_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(_03753_),
    .A1(_03841_),
    .S(_03705_),
    .X(_03933_));
 sky130_fd_sc_hd__a211o_1 _09838_ (.A1(_03815_),
    .A2(_03689_),
    .B1(_03669_),
    .C1(_03697_),
    .X(_03934_));
 sky130_fd_sc_hd__a2bb2o_1 _09839_ (.A1_N(_03651_),
    .A2_N(_03720_),
    .B1(_03674_),
    .B2(_03648_),
    .X(_03936_));
 sky130_fd_sc_hd__a21oi_1 _09840_ (.A1(_03874_),
    .A2(_03802_),
    .B1(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__a221o_1 _09841_ (.A1(_03700_),
    .A2(_03768_),
    .B1(_03937_),
    .B2(_03934_),
    .C1(_03706_),
    .X(_03938_));
 sky130_fd_sc_hd__o211ai_1 _09842_ (.A1(_03933_),
    .A2(_03707_),
    .B1(_03739_),
    .C1(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__o211a_1 _09843_ (.A1(_03892_),
    .A2(_03893_),
    .B1(_03932_),
    .C1(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__a41oi_2 _09844_ (.A1(_03733_),
    .A2(_03928_),
    .A3(_03738_),
    .A4(_03809_),
    .B1(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__nor2_1 _09845_ (.A(_03823_),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__a221o_1 _09846_ (.A1(_03811_),
    .A2(_03899_),
    .B1(_03901_),
    .B2(_03845_),
    .C1(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__a22oi_4 _09847_ (.A1(_03845_),
    .A2(_03849_),
    .B1(_03943_),
    .B2(_03835_),
    .Y(_03944_));
 sky130_fd_sc_hd__o21ai_4 _09848_ (.A1(_03833_),
    .A2(_03903_),
    .B1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__nand2_8 _09849_ (.A(_03945_),
    .B(_03915_),
    .Y(_03947_));
 sky130_fd_sc_hd__or4b_4 _09850_ (.A(_03573_),
    .B(_03850_),
    .C(_03912_),
    .D_N(_03945_),
    .X(_03948_));
 sky130_fd_sc_hd__o21a_4 _09851_ (.A1(_03573_),
    .A2(_03947_),
    .B1(net65),
    .X(_03949_));
 sky130_fd_sc_hd__o21ai_2 _09852_ (.A1(_03573_),
    .A2(_03947_),
    .B1(net65),
    .Y(_03950_));
 sky130_fd_sc_hd__and3_1 _09853_ (.A(_03007_),
    .B(net100),
    .C(_03949_),
    .X(_03951_));
 sky130_fd_sc_hd__a31o_1 _09854_ (.A1(_02981_),
    .A2(_02983_),
    .A3(_02997_),
    .B1(_03951_),
    .X(net66));
 sky130_fd_sc_hd__o211a_1 _09855_ (.A1(_01788_),
    .A2(_01789_),
    .B1(_01913_),
    .C1(_02929_),
    .X(_03952_));
 sky130_fd_sc_hd__or2_1 _09856_ (.A(_02930_),
    .B(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__nand2_1 _09857_ (.A(_02977_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__o211a_1 _09858_ (.A1(_02977_),
    .A2(_02982_),
    .B1(_02997_),
    .C1(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__a21oi_2 _09859_ (.A1(_03915_),
    .A2(_03945_),
    .B1(_03950_),
    .Y(_03957_));
 sky130_fd_sc_hd__a31o_1 _09860_ (.A1(net65),
    .A2(_03646_),
    .A3(_03948_),
    .B1(_03955_),
    .X(net77));
 sky130_fd_sc_hd__or3_1 _09861_ (.A(_01667_),
    .B(_01788_),
    .C(_02930_),
    .X(_03958_));
 sky130_fd_sc_hd__and2_1 _09862_ (.A(_02931_),
    .B(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__or4b_1 _09863_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_03953_),
    .X(_03960_));
 sky130_fd_sc_hd__o21a_1 _09864_ (.A1(_02976_),
    .A2(_03959_),
    .B1(_02997_),
    .X(_03961_));
 sky130_fd_sc_hd__and3_1 _09865_ (.A(_03775_),
    .B(net65),
    .C(_03406_),
    .X(_03962_));
 sky130_fd_sc_hd__a21o_1 _09866_ (.A1(_03960_),
    .A2(_03961_),
    .B1(_03962_),
    .X(net88));
 sky130_fd_sc_hd__and3_1 _09867_ (.A(_01665_),
    .B(_02931_),
    .C(_02933_),
    .X(_03963_));
 sky130_fd_sc_hd__or2_1 _09868_ (.A(_02934_),
    .B(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__nand2_1 _09869_ (.A(_02977_),
    .B(_03964_),
    .Y(_03966_));
 sky130_fd_sc_hd__or4_1 _09870_ (.A(_02972_),
    .B(_03959_),
    .C(_02973_),
    .D(_02971_),
    .X(_03967_));
 sky130_fd_sc_hd__o221a_1 _09871_ (.A1(_03398_),
    .A2(_03404_),
    .B1(_03548_),
    .B2(_03366_),
    .C1(_03758_),
    .X(_03968_));
 sky130_fd_sc_hd__a211o_1 _09872_ (.A1(_03775_),
    .A2(_03574_),
    .B1(_03968_),
    .C1(_03915_),
    .X(_03969_));
 sky130_fd_sc_hd__and3_1 _09873_ (.A(_03916_),
    .B(_03969_),
    .C(net65),
    .X(_03970_));
 sky130_fd_sc_hd__a31o_1 _09874_ (.A1(_03966_),
    .A2(_03967_),
    .A3(_02997_),
    .B1(_03970_),
    .X(net91));
 sky130_fd_sc_hd__and2_1 _09875_ (.A(_02936_),
    .B(_01419_),
    .X(_03971_));
 sky130_fd_sc_hd__or2_1 _09876_ (.A(_02937_),
    .B(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__o31a_1 _09877_ (.A1(_02971_),
    .A2(_02972_),
    .A3(_02973_),
    .B1(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__a2111oi_1 _09878_ (.A1(_02976_),
    .A2(_03964_),
    .B1(_02996_),
    .C1(_02989_),
    .D1(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__a21oi_1 _09879_ (.A1(_03408_),
    .A2(_03416_),
    .B1(_03776_),
    .Y(_03976_));
 sky130_fd_sc_hd__a31o_1 _09880_ (.A1(net65),
    .A2(_03947_),
    .A3(_03976_),
    .B1(_03974_),
    .X(net92));
 sky130_fd_sc_hd__or4b_1 _09881_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_03972_),
    .X(_03977_));
 sky130_fd_sc_hd__a211oi_1 _09882_ (.A1(_01416_),
    .A2(_01414_),
    .B1(_01293_),
    .C1(_02937_),
    .Y(_03978_));
 sky130_fd_sc_hd__nor2_1 _09883_ (.A(_02938_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__a21o_1 _09884_ (.A1(_02970_),
    .A2(_02974_),
    .B1(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__o221a_1 _09885_ (.A1(_03424_),
    .A2(_03762_),
    .B1(_03776_),
    .B2(_03617_),
    .C1(_03916_),
    .X(_03981_));
 sky130_fd_sc_hd__nor2_1 _09886_ (.A(_03981_),
    .B(_03950_),
    .Y(_03982_));
 sky130_fd_sc_hd__a32o_1 _09887_ (.A1(_03977_),
    .A2(_03980_),
    .A3(_02997_),
    .B1(_03982_),
    .B2(_03916_),
    .X(net93));
 sky130_fd_sc_hd__o211a_1 _09888_ (.A1(_03424_),
    .A2(_03754_),
    .B1(_03648_),
    .C1(_03777_),
    .X(_03983_));
 sky130_fd_sc_hd__and3_1 _09889_ (.A(_03835_),
    .B(_03842_),
    .C(_03903_),
    .X(_03985_));
 sky130_fd_sc_hd__nor3_1 _09890_ (.A(_01156_),
    .B(_01291_),
    .C(_02938_),
    .Y(_03986_));
 sky130_fd_sc_hd__nor2_1 _09891_ (.A(_02939_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__mux2_1 _09892_ (.A0(_03987_),
    .A1(_03979_),
    .S(_02976_),
    .X(_03988_));
 sky130_fd_sc_hd__a22o_1 _09893_ (.A1(_03957_),
    .A2(_03983_),
    .B1(_03988_),
    .B2(_02997_),
    .X(net94));
 sky130_fd_sc_hd__a211oi_1 _09894_ (.A1(_01150_),
    .A2(_01152_),
    .B1(_02939_),
    .C1(_01023_),
    .Y(_03989_));
 sky130_fd_sc_hd__nor2_1 _09895_ (.A(_02940_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__mux2_1 _09896_ (.A0(_03990_),
    .A1(_03987_),
    .S(_02976_),
    .X(_03991_));
 sky130_fd_sc_hd__and3_1 _09897_ (.A(_03916_),
    .B(_03782_),
    .C(net65),
    .X(_03992_));
 sky130_fd_sc_hd__a21o_1 _09898_ (.A1(_02997_),
    .A2(_03991_),
    .B1(_03992_),
    .X(net95));
 sky130_fd_sc_hd__a22o_1 _09899_ (.A1(_03669_),
    .A2(_03844_),
    .B1(_03780_),
    .B2(_03874_),
    .X(_03994_));
 sky130_fd_sc_hd__or4_1 _09900_ (.A(_02972_),
    .B(_03990_),
    .C(_02973_),
    .D(_02971_),
    .X(_03995_));
 sky130_fd_sc_hd__nor3_1 _09901_ (.A(_00903_),
    .B(_01022_),
    .C(_02940_),
    .Y(_03996_));
 sky130_fd_sc_hd__nor2_1 _09902_ (.A(_02941_),
    .B(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__a2bb2o_1 _09903_ (.A1_N(_02941_),
    .A2_N(_03996_),
    .B1(_02974_),
    .B2(_02970_),
    .X(_03998_));
 sky130_fd_sc_hd__a32o_1 _09904_ (.A1(_03995_),
    .A2(_03998_),
    .A3(_02997_),
    .B1(_03957_),
    .B2(_03994_),
    .X(net96));
 sky130_fd_sc_hd__nor3_1 _09905_ (.A(_00901_),
    .B(_02941_),
    .C(_02942_),
    .Y(_03999_));
 sky130_fd_sc_hd__nor2_1 _09906_ (.A(_02943_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__mux2_1 _09907_ (.A0(_04000_),
    .A1(_03997_),
    .S(_02976_),
    .X(_04001_));
 sky130_fd_sc_hd__o31a_1 _09908_ (.A1(_03669_),
    .A2(_03689_),
    .A3(_03697_),
    .B1(_03906_),
    .X(_04002_));
 sky130_fd_sc_hd__and3_1 _09909_ (.A(_03916_),
    .B(_04002_),
    .C(net65),
    .X(_04004_));
 sky130_fd_sc_hd__a21o_1 _09910_ (.A1(_02997_),
    .A2(_04001_),
    .B1(_04004_),
    .X(net97));
 sky130_fd_sc_hd__xnor2_1 _09911_ (.A(_00692_),
    .B(_02944_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand2_1 _09912_ (.A(_02977_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__or4_1 _09913_ (.A(_02972_),
    .B(_04000_),
    .C(_02973_),
    .D(_02971_),
    .X(_04007_));
 sky130_fd_sc_hd__o211a_1 _09914_ (.A1(_03701_),
    .A2(_03906_),
    .B1(_03904_),
    .C1(_03707_),
    .X(_04008_));
 sky130_fd_sc_hd__and3_1 _09915_ (.A(_03949_),
    .B(_04008_),
    .C(_03916_),
    .X(_04009_));
 sky130_fd_sc_hd__a31o_1 _09916_ (.A1(_04006_),
    .A2(_04007_),
    .A3(_02997_),
    .B1(_04009_),
    .X(net67));
 sky130_fd_sc_hd__xnor2_1 _09917_ (.A(_00601_),
    .B(_02945_),
    .Y(_04010_));
 sky130_fd_sc_hd__mux2_1 _09918_ (.A0(_04010_),
    .A1(_04005_),
    .S(_02976_),
    .X(_04011_));
 sky130_fd_sc_hd__nor3_1 _09919_ (.A(_02989_),
    .B(_02996_),
    .C(_04011_),
    .Y(_04013_));
 sky130_fd_sc_hd__a31o_1 _09920_ (.A1(net65),
    .A2(_03909_),
    .A3(_03947_),
    .B1(_04013_),
    .X(net68));
 sky130_fd_sc_hd__and3_1 _09921_ (.A(_00509_),
    .B(_00599_),
    .C(_02947_),
    .X(_04014_));
 sky130_fd_sc_hd__nor2_1 _09922_ (.A(_02948_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__or4b_1 _09923_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_04010_),
    .X(_04016_));
 sky130_fd_sc_hd__o211a_1 _09924_ (.A1(_02976_),
    .A2(_04015_),
    .B1(_02997_),
    .C1(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__a2bb2o_1 _09925_ (.A1_N(_03738_),
    .A2_N(_03928_),
    .B1(_03828_),
    .B2(_03833_),
    .X(_04018_));
 sky130_fd_sc_hd__a31o_1 _09926_ (.A1(_03837_),
    .A2(_03949_),
    .A3(_04018_),
    .B1(_04017_),
    .X(net69));
 sky130_fd_sc_hd__and4_1 _09927_ (.A(_03784_),
    .B(_03916_),
    .C(_03931_),
    .D(net65),
    .X(_04019_));
 sky130_fd_sc_hd__and2_1 _09928_ (.A(_02949_),
    .B(_00424_),
    .X(_04020_));
 sky130_fd_sc_hd__or2_1 _09929_ (.A(_02950_),
    .B(_04020_),
    .X(_04022_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(_02977_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__or4_1 _09931_ (.A(_02972_),
    .B(_04015_),
    .C(_02973_),
    .D(_02971_),
    .X(_04024_));
 sky130_fd_sc_hd__a31o_1 _09932_ (.A1(_04023_),
    .A2(_04024_),
    .A3(_02997_),
    .B1(_04019_),
    .X(net70));
 sky130_fd_sc_hd__xnor2_1 _09933_ (.A(_02951_),
    .B(_02953_),
    .Y(_04025_));
 sky130_fd_sc_hd__nand2_1 _09934_ (.A(_02977_),
    .B(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__or4b_1 _09935_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_04022_),
    .X(_04027_));
 sky130_fd_sc_hd__a31o_1 _09936_ (.A1(_03705_),
    .A2(_03706_),
    .A3(_03736_),
    .B1(_03892_),
    .X(_04028_));
 sky130_fd_sc_hd__or3b_1 _09937_ (.A(_03713_),
    .B(_03845_),
    .C_N(_03736_),
    .X(_04029_));
 sky130_fd_sc_hd__a22o_1 _09938_ (.A1(_03734_),
    .A2(_03736_),
    .B1(_04028_),
    .B2(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__or4_1 _09939_ (.A(_03732_),
    .B(_03739_),
    .C(_03809_),
    .D(_03928_),
    .X(_04032_));
 sky130_fd_sc_hd__a31oi_1 _09940_ (.A1(_03916_),
    .A2(_04030_),
    .A3(_04032_),
    .B1(_03950_),
    .Y(_04033_));
 sky130_fd_sc_hd__a32o_1 _09941_ (.A1(_04026_),
    .A2(_04027_),
    .A3(_02997_),
    .B1(_04033_),
    .B2(_03916_),
    .X(net71));
 sky130_fd_sc_hd__a2bb2o_1 _09942_ (.A1_N(_03912_),
    .A2_N(_03850_),
    .B1(_03823_),
    .B2(_03941_),
    .X(_04034_));
 sky130_fd_sc_hd__and3_1 _09943_ (.A(_03916_),
    .B(_04034_),
    .C(net65),
    .X(_04035_));
 sky130_fd_sc_hd__xnor2_1 _09944_ (.A(_02954_),
    .B(_02955_),
    .Y(_04036_));
 sky130_fd_sc_hd__or4b_1 _09945_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_04025_),
    .X(_04037_));
 sky130_fd_sc_hd__o21a_1 _09946_ (.A1(_02976_),
    .A2(_04036_),
    .B1(_02997_),
    .X(_04038_));
 sky130_fd_sc_hd__a21o_1 _09947_ (.A1(_04037_),
    .A2(_04038_),
    .B1(_04035_),
    .X(net72));
 sky130_fd_sc_hd__and4b_1 _09948_ (.A_N(_03943_),
    .B(_03949_),
    .C(_03834_),
    .D(_03916_),
    .X(_04039_));
 sky130_fd_sc_hd__or4_1 _09949_ (.A(_02972_),
    .B(_04036_),
    .C(_02973_),
    .D(_02971_),
    .X(_04041_));
 sky130_fd_sc_hd__nand2_1 _09950_ (.A(_02956_),
    .B(_00197_),
    .Y(_04042_));
 sky130_fd_sc_hd__nand2_1 _09951_ (.A(_02958_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand2_1 _09952_ (.A(_02977_),
    .B(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__a31o_1 _09953_ (.A1(_04044_),
    .A2(_02997_),
    .A3(_04041_),
    .B1(_04039_),
    .X(net73));
 sky130_fd_sc_hd__and3_1 _09954_ (.A(_00136_),
    .B(_00195_),
    .C(_02958_),
    .X(_04045_));
 sky130_fd_sc_hd__nor2_1 _09955_ (.A(_02959_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__a21o_1 _09956_ (.A1(_02970_),
    .A2(_02974_),
    .B1(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__or4b_1 _09957_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_04043_),
    .X(_04048_));
 sky130_fd_sc_hd__a2bb2o_1 _09958_ (.A1_N(_03706_),
    .A2_N(_03805_),
    .B1(_03818_),
    .B2(_03692_),
    .X(_04049_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(_04049_),
    .A1(_03768_),
    .S(_03712_),
    .X(_04051_));
 sky130_fd_sc_hd__a21oi_1 _09960_ (.A1(_03739_),
    .A2(_04051_),
    .B1(_03783_),
    .Y(_04052_));
 sky130_fd_sc_hd__a32o_1 _09961_ (.A1(_03734_),
    .A2(_03736_),
    .A3(_03842_),
    .B1(_04052_),
    .B2(_03829_),
    .X(_04053_));
 sky130_fd_sc_hd__o31a_1 _09962_ (.A1(_03732_),
    .A2(_03739_),
    .A3(_03808_),
    .B1(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__o211a_1 _09963_ (.A1(_03767_),
    .A2(_03845_),
    .B1(_03810_),
    .C1(_03821_),
    .X(_04055_));
 sky130_fd_sc_hd__a211o_1 _09964_ (.A1(_03901_),
    .A2(_03899_),
    .B1(_04055_),
    .C1(_04054_),
    .X(_04056_));
 sky130_fd_sc_hd__o31ai_1 _09965_ (.A1(_03828_),
    .A2(_03834_),
    .A3(_03943_),
    .B1(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__and3_1 _09966_ (.A(_03916_),
    .B(_04057_),
    .C(net65),
    .X(_04058_));
 sky130_fd_sc_hd__a31o_1 _09967_ (.A1(_04048_),
    .A2(_02997_),
    .A3(_04047_),
    .B1(_04058_),
    .X(net74));
 sky130_fd_sc_hd__or4_1 _09968_ (.A(_02972_),
    .B(_04046_),
    .C(_02973_),
    .D(_02971_),
    .X(_04059_));
 sky130_fd_sc_hd__a211oi_1 _09969_ (.A1(_00133_),
    .A2(_00131_),
    .B1(_00083_),
    .C1(_02959_),
    .Y(_04061_));
 sky130_fd_sc_hd__nor2_1 _09970_ (.A(_02960_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__o211ai_1 _09971_ (.A1(_02976_),
    .A2(_04062_),
    .B1(_02997_),
    .C1(_04059_),
    .Y(_04063_));
 sky130_fd_sc_hd__o31ai_1 _09972_ (.A1(_03910_),
    .A2(_03945_),
    .A3(_03950_),
    .B1(_04063_),
    .Y(net75));
 sky130_fd_sc_hd__or3_1 _09973_ (.A(_05392_),
    .B(_00081_),
    .C(_02960_),
    .X(_04064_));
 sky130_fd_sc_hd__nand2_1 _09974_ (.A(_02961_),
    .B(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand2_1 _09975_ (.A(_02977_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__or4_1 _09976_ (.A(_02972_),
    .B(_04062_),
    .C(_02973_),
    .D(_02971_),
    .X(_04067_));
 sky130_fd_sc_hd__a22o_1 _09977_ (.A1(_03911_),
    .A2(_03914_),
    .B1(_03944_),
    .B2(_03985_),
    .X(_04068_));
 sky130_fd_sc_hd__a32o_1 _09978_ (.A1(_04066_),
    .A2(_04067_),
    .A3(_02997_),
    .B1(_04068_),
    .B2(_03957_),
    .X(net76));
 sky130_fd_sc_hd__o211a_1 _09979_ (.A1(_03833_),
    .A2(_03903_),
    .B1(_03910_),
    .C1(_03944_),
    .X(_04070_));
 sky130_fd_sc_hd__a2111oi_1 _09980_ (.A1(_03821_),
    .A2(_03841_),
    .B1(_03768_),
    .C1(_03784_),
    .D1(_03808_),
    .Y(_04071_));
 sky130_fd_sc_hd__a21oi_1 _09981_ (.A1(_03821_),
    .A2(_03828_),
    .B1(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__a211o_1 _09982_ (.A1(_03835_),
    .A2(_03903_),
    .B1(_04070_),
    .C1(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__o211a_1 _09983_ (.A1(_03850_),
    .A2(_03911_),
    .B1(_04073_),
    .C1(_03957_),
    .X(_04074_));
 sky130_fd_sc_hd__xor2_1 _09984_ (.A(_05349_),
    .B(_02963_),
    .X(_04075_));
 sky130_fd_sc_hd__a21o_1 _09985_ (.A1(_02970_),
    .A2(_02974_),
    .B1(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__or4b_1 _09986_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_04065_),
    .X(_04077_));
 sky130_fd_sc_hd__a31o_1 _09987_ (.A1(_04077_),
    .A2(_02997_),
    .A3(_04076_),
    .B1(_04074_),
    .X(net78));
 sky130_fd_sc_hd__or4_1 _09988_ (.A(_02972_),
    .B(_04075_),
    .C(_02973_),
    .D(_02971_),
    .X(_04078_));
 sky130_fd_sc_hd__xnor2_1 _09989_ (.A(_02964_),
    .B(_02967_),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _09990_ (.A(_02977_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a31o_1 _09991_ (.A1(_04081_),
    .A2(_02997_),
    .A3(_04078_),
    .B1(_03957_),
    .X(net79));
 sky130_fd_sc_hd__o22a_1 _09992_ (.A1(_02972_),
    .A2(_02970_),
    .B1(_05305_),
    .B2(_02975_),
    .X(_04082_));
 sky130_fd_sc_hd__a21o_1 _09993_ (.A1(_02972_),
    .A2(_02973_),
    .B1(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__or4b_1 _09994_ (.A(_02971_),
    .B(_02972_),
    .C(_02973_),
    .D_N(_04080_),
    .X(_04084_));
 sky130_fd_sc_hd__a32o_1 _09995_ (.A1(_04083_),
    .A2(_04084_),
    .A3(_02997_),
    .B1(_03573_),
    .B2(net65),
    .X(net80));
 sky130_fd_sc_hd__or4_1 _09996_ (.A(_02143_),
    .B(_02971_),
    .C(_02972_),
    .D(_02973_),
    .X(_04085_));
 sky130_fd_sc_hd__a2bb2o_2 _09997_ (.A1_N(_02110_),
    .A2_N(_02121_),
    .B1(_02970_),
    .B2(_02974_),
    .X(_04086_));
 sky130_fd_sc_hd__a21oi_1 _09998_ (.A1(_04085_),
    .A2(_04086_),
    .B1(_02996_),
    .Y(_04087_));
 sky130_fd_sc_hd__and3_2 _09999_ (.A(_01010_),
    .B(_02000_),
    .C(_02022_),
    .X(_04089_));
 sky130_fd_sc_hd__and3_2 _10000_ (.A(_01021_),
    .B(_02044_),
    .C(_02066_),
    .X(_04090_));
 sky130_fd_sc_hd__a31o_4 _10001_ (.A1(_01010_),
    .A2(_02000_),
    .A3(_02022_),
    .B1(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__a21oi_1 _10002_ (.A1(_01010_),
    .A2(_02077_),
    .B1(_04090_),
    .Y(_04092_));
 sky130_fd_sc_hd__o2bb2a_2 _10003_ (.A1_N(_03381_),
    .A2_N(_03386_),
    .B1(_03398_),
    .B2(_03375_),
    .X(_04093_));
 sky130_fd_sc_hd__o22ai_4 _10004_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_04093_),
    .B2(_03365_),
    .Y(_04094_));
 sky130_fd_sc_hd__or4_2 _10005_ (.A(_03402_),
    .B(_04091_),
    .C(_03365_),
    .D(_03373_),
    .X(_04095_));
 sky130_fd_sc_hd__o31a_4 _10006_ (.A1(_03365_),
    .A2(_04091_),
    .A3(_04093_),
    .B1(_04094_),
    .X(_04096_));
 sky130_fd_sc_hd__o31ai_4 _10007_ (.A1(_03365_),
    .A2(_04091_),
    .A3(_04093_),
    .B1(_04094_),
    .Y(_04097_));
 sky130_fd_sc_hd__and4_2 _10008_ (.A(_03640_),
    .B(_03644_),
    .C(_04096_),
    .D(_03600_),
    .X(_04098_));
 sky130_fd_sc_hd__nand4_1 _10009_ (.A(_03640_),
    .B(_03644_),
    .C(_04096_),
    .D(_03600_),
    .Y(_04100_));
 sky130_fd_sc_hd__a211o_1 _10010_ (.A1(_03087_),
    .A2(net101),
    .B1(_03596_),
    .C1(net103),
    .X(_04101_));
 sky130_fd_sc_hd__o32a_1 _10011_ (.A1(_03409_),
    .A2(_03417_),
    .A3(_04101_),
    .B1(_04097_),
    .B2(_03615_),
    .X(_04102_));
 sky130_fd_sc_hd__a2bb2o_1 _10012_ (.A1_N(_03425_),
    .A2_N(_04101_),
    .B1(_03617_),
    .B2(_04096_),
    .X(_04103_));
 sky130_fd_sc_hd__o21ai_1 _10013_ (.A1(_03601_),
    .A2(_03643_),
    .B1(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__and3_1 _10014_ (.A(_03644_),
    .B(_04097_),
    .C(_03600_),
    .X(_04105_));
 sky130_fd_sc_hd__nand3_1 _10015_ (.A(_03644_),
    .B(_04097_),
    .C(_03600_),
    .Y(_04106_));
 sky130_fd_sc_hd__o22a_1 _10016_ (.A1(_03640_),
    .A2(_04106_),
    .B1(_04102_),
    .B2(_03647_),
    .X(_04107_));
 sky130_fd_sc_hd__o311a_4 _10017_ (.A1(_03640_),
    .A2(_03648_),
    .A3(_04096_),
    .B1(_04100_),
    .C1(_04104_),
    .X(_04108_));
 sky130_fd_sc_hd__a221o_1 _10018_ (.A1(_03648_),
    .A2(_04103_),
    .B1(_04105_),
    .B2(_03639_),
    .C1(_04098_),
    .X(_04109_));
 sky130_fd_sc_hd__and3_2 _10019_ (.A(_03706_),
    .B(_04109_),
    .C(_03705_),
    .X(_04111_));
 sky130_fd_sc_hd__a21o_1 _10020_ (.A1(_04100_),
    .A2(_04107_),
    .B1(_03713_),
    .X(_04112_));
 sky130_fd_sc_hd__nor3b_2 _10021_ (.A(_04096_),
    .B(_03669_),
    .C_N(_03695_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand4_4 _10022_ (.A(_03647_),
    .B(_03695_),
    .C(_04097_),
    .D(_03640_),
    .Y(_04114_));
 sky130_fd_sc_hd__o21ai_2 _10023_ (.A1(_03698_),
    .A2(_04108_),
    .B1(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__o21ai_2 _10024_ (.A1(_03689_),
    .A2(_03699_),
    .B1(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__or3_1 _10025_ (.A(_04108_),
    .B(_03701_),
    .C(_03692_),
    .X(_04117_));
 sky130_fd_sc_hd__nand4_4 _10026_ (.A(_03690_),
    .B(_03692_),
    .C(_03698_),
    .D(_04108_),
    .Y(_04118_));
 sky130_fd_sc_hd__or4bb_2 _10027_ (.A(_03701_),
    .B(_03705_),
    .C_N(_04108_),
    .D_N(_03692_),
    .X(_04119_));
 sky130_fd_sc_hd__and4_4 _10028_ (.A(_04112_),
    .B(_04116_),
    .C(_04117_),
    .D(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__nand4_4 _10029_ (.A(_04112_),
    .B(_04116_),
    .C(_04117_),
    .D(_04119_),
    .Y(_04122_));
 sky130_fd_sc_hd__or3_1 _10030_ (.A(_03768_),
    .B(_03823_),
    .C(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__a31o_1 _10031_ (.A1(_03712_),
    .A2(_03732_),
    .A3(_03736_),
    .B1(_04122_),
    .X(_04124_));
 sky130_fd_sc_hd__nand4_1 _10032_ (.A(_04122_),
    .B(_03732_),
    .C(_03712_),
    .D(_03736_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_04124_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__and3_2 _10034_ (.A(_03783_),
    .B(_04120_),
    .C(_03809_),
    .X(_04127_));
 sky130_fd_sc_hd__and3_1 _10035_ (.A(_03811_),
    .B(_04124_),
    .C(_04125_),
    .X(_04128_));
 sky130_fd_sc_hd__o21ai_1 _10036_ (.A1(_04127_),
    .A2(_04128_),
    .B1(_03823_),
    .Y(_04129_));
 sky130_fd_sc_hd__a211o_4 _10037_ (.A1(_03783_),
    .A2(_03819_),
    .B1(_04120_),
    .C1(_03811_),
    .X(_04130_));
 sky130_fd_sc_hd__o221ai_4 _10038_ (.A1(_03834_),
    .A2(_04122_),
    .B1(_04130_),
    .B2(_03767_),
    .C1(_04129_),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _10039_ (.A(_03837_),
    .B(_04131_),
    .Y(_04133_));
 sky130_fd_sc_hd__or4b_4 _10040_ (.A(_03768_),
    .B(_04120_),
    .C(_03823_),
    .D_N(_03828_),
    .X(_04134_));
 sky130_fd_sc_hd__or3_1 _10041_ (.A(_03837_),
    .B(_03841_),
    .C(_04122_),
    .X(_04135_));
 sky130_fd_sc_hd__nor2_1 _10042_ (.A(_03912_),
    .B(_04131_),
    .Y(_04136_));
 sky130_fd_sc_hd__o2bb2a_1 _10043_ (.A1_N(_04133_),
    .A2_N(_04134_),
    .B1(_03837_),
    .B2(_03841_),
    .X(_04137_));
 sky130_fd_sc_hd__a31o_1 _10044_ (.A1(_03903_),
    .A2(_03910_),
    .A3(_04120_),
    .B1(_04136_),
    .X(_04138_));
 sky130_fd_sc_hd__or4_1 _10045_ (.A(_03837_),
    .B(_03841_),
    .C(_04131_),
    .D(_03903_),
    .X(_04139_));
 sky130_fd_sc_hd__o21ai_1 _10046_ (.A1(_04137_),
    .A2(_04138_),
    .B1(_03916_),
    .Y(_04140_));
 sky130_fd_sc_hd__nand2_1 _10047_ (.A(_03915_),
    .B(_04131_),
    .Y(_04141_));
 sky130_fd_sc_hd__o221a_1 _10048_ (.A1(_03947_),
    .A2(_04131_),
    .B1(_04141_),
    .B2(_03945_),
    .C1(_03948_),
    .X(_04142_));
 sky130_fd_sc_hd__o2bb2a_1 _10049_ (.A1_N(_04140_),
    .A2_N(_04142_),
    .B1(_03948_),
    .B2(net103),
    .X(_04144_));
 sky130_fd_sc_hd__a2bb2o_1 _10050_ (.A1_N(_02989_),
    .A2_N(_04087_),
    .B1(_04144_),
    .B2(net65),
    .X(net81));
 sky130_fd_sc_hd__o21a_1 _10051_ (.A1(net48),
    .A2(net16),
    .B1(_01604_),
    .X(_04145_));
 sky130_fd_sc_hd__or3_1 _10052_ (.A(_01582_),
    .B(_01593_),
    .C(_02110_),
    .X(_04146_));
 sky130_fd_sc_hd__or3_1 _10053_ (.A(net48),
    .B(net16),
    .C(_01604_),
    .X(_04147_));
 sky130_fd_sc_hd__nand2_1 _10054_ (.A(_04146_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__a22o_1 _10055_ (.A1(_02143_),
    .A2(_02977_),
    .B1(_04146_),
    .B2(_04147_),
    .X(_04149_));
 sky130_fd_sc_hd__or3_1 _10056_ (.A(_02132_),
    .B(_04148_),
    .C(_02976_),
    .X(_04150_));
 sky130_fd_sc_hd__a21oi_1 _10057_ (.A1(_04149_),
    .A2(_04150_),
    .B1(_02996_),
    .Y(_04151_));
 sky130_fd_sc_hd__o211a_1 _10058_ (.A1(_03677_),
    .A2(_04109_),
    .B1(_03705_),
    .C1(_03706_),
    .X(_04152_));
 sky130_fd_sc_hd__a311o_1 _10059_ (.A1(net114),
    .A2(_03370_),
    .A3(_03372_),
    .B1(_04091_),
    .C1(_03368_),
    .X(_04154_));
 sky130_fd_sc_hd__nand4_2 _10060_ (.A(net99),
    .B(_03389_),
    .C(_03399_),
    .D(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__and4_1 _10061_ (.A(net99),
    .B(_03389_),
    .C(_03399_),
    .D(_04154_),
    .X(_04156_));
 sky130_fd_sc_hd__a211o_1 _10062_ (.A1(_03380_),
    .A2(_03379_),
    .B1(_04091_),
    .C1(_03387_),
    .X(_04157_));
 sky130_fd_sc_hd__a22oi_4 _10063_ (.A1(net103),
    .A2(_03388_),
    .B1(net101),
    .B2(_03087_),
    .Y(_04158_));
 sky130_fd_sc_hd__a21oi_2 _10064_ (.A1(_02000_),
    .A2(_02022_),
    .B1(net17),
    .Y(_04159_));
 sky130_fd_sc_hd__and3_1 _10065_ (.A(_00999_),
    .B(_02000_),
    .C(_02022_),
    .X(_04160_));
 sky130_fd_sc_hd__and3_1 _10066_ (.A(_02066_),
    .B(net17),
    .C(_02044_),
    .X(_04161_));
 sky130_fd_sc_hd__and3_1 _10067_ (.A(_02022_),
    .B(net49),
    .C(_02000_),
    .X(_04162_));
 sky130_fd_sc_hd__a31o_4 _10068_ (.A1(net49),
    .A2(_02000_),
    .A3(_02022_),
    .B1(_04161_),
    .X(_04163_));
 sky130_fd_sc_hd__a31o_2 _10069_ (.A1(_00999_),
    .A2(_02000_),
    .A3(_02022_),
    .B1(_04159_),
    .X(_04165_));
 sky130_fd_sc_hd__o22a_1 _10070_ (.A1(_04159_),
    .A2(_04160_),
    .B1(_04091_),
    .B2(_03389_),
    .X(_04166_));
 sky130_fd_sc_hd__a31o_1 _10071_ (.A1(_03381_),
    .A2(_03386_),
    .A3(net103),
    .B1(_04163_),
    .X(_04167_));
 sky130_fd_sc_hd__a21o_1 _10072_ (.A1(_03087_),
    .A2(net101),
    .B1(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__o2bb2ai_1 _10073_ (.A1_N(net99),
    .A2_N(_04157_),
    .B1(_04161_),
    .B2(_04162_),
    .Y(_04169_));
 sky130_fd_sc_hd__o211a_4 _10074_ (.A1(_03389_),
    .A2(_04091_),
    .B1(_04163_),
    .C1(net99),
    .X(_04170_));
 sky130_fd_sc_hd__o211ai_1 _10075_ (.A1(_03389_),
    .A2(_04091_),
    .B1(_04163_),
    .C1(net99),
    .Y(_04171_));
 sky130_fd_sc_hd__a21oi_2 _10076_ (.A1(net99),
    .A2(_04157_),
    .B1(_04163_),
    .Y(_04172_));
 sky130_fd_sc_hd__o2bb2ai_1 _10077_ (.A1_N(net99),
    .A2_N(_04157_),
    .B1(_04159_),
    .B2(_04160_),
    .Y(_04173_));
 sky130_fd_sc_hd__o21ai_4 _10078_ (.A1(_04163_),
    .A2(_04158_),
    .B1(_04155_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand3_1 _10079_ (.A(_04173_),
    .B(_04155_),
    .C(_04171_),
    .Y(_04176_));
 sky130_fd_sc_hd__o2111a_2 _10080_ (.A1(_03375_),
    .A2(_04091_),
    .B1(_04163_),
    .C1(_03399_),
    .D1(_03403_),
    .X(_04177_));
 sky130_fd_sc_hd__o2111ai_4 _10081_ (.A1(_03375_),
    .A2(_04091_),
    .B1(_04163_),
    .C1(_03399_),
    .D1(_03403_),
    .Y(_04178_));
 sky130_fd_sc_hd__o21a_1 _10082_ (.A1(_04170_),
    .A2(_04174_),
    .B1(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__o21ai_1 _10083_ (.A1(_04170_),
    .A2(_04174_),
    .B1(_04178_),
    .Y(_04180_));
 sky130_fd_sc_hd__or4_1 _10084_ (.A(_03417_),
    .B(_03597_),
    .C(_04091_),
    .D(_03409_),
    .X(_04181_));
 sky130_fd_sc_hd__o2111a_1 _10085_ (.A1(_04170_),
    .A2(_04174_),
    .B1(_03600_),
    .C1(_04178_),
    .D1(_04096_),
    .X(_04182_));
 sky130_fd_sc_hd__o2111ai_4 _10086_ (.A1(_04170_),
    .A2(_04174_),
    .B1(_03600_),
    .C1(_04178_),
    .D1(_04096_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand4_2 _10087_ (.A(_03405_),
    .B(_03416_),
    .C(_04091_),
    .D(_03375_),
    .Y(_04184_));
 sky130_fd_sc_hd__a22oi_2 _10088_ (.A1(_03424_),
    .A2(_04091_),
    .B1(_04176_),
    .B2(_04178_),
    .Y(_04185_));
 sky130_fd_sc_hd__nor2_2 _10089_ (.A(_04184_),
    .B(_04177_),
    .Y(_04187_));
 sky130_fd_sc_hd__o22ai_4 _10090_ (.A1(_04091_),
    .A2(_03601_),
    .B1(_04187_),
    .B2(_04185_),
    .Y(_04188_));
 sky130_fd_sc_hd__o31a_2 _10091_ (.A1(_03601_),
    .A2(_04097_),
    .A3(_04180_),
    .B1(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__o21ai_1 _10092_ (.A1(_04180_),
    .A2(_04181_),
    .B1(_04188_),
    .Y(_04190_));
 sky130_fd_sc_hd__a2bb2oi_2 _10093_ (.A1_N(_03648_),
    .A2_N(_04096_),
    .B1(_04183_),
    .B2(_04188_),
    .Y(_04191_));
 sky130_fd_sc_hd__o2bb2ai_4 _10094_ (.A1_N(_04183_),
    .A2_N(_04188_),
    .B1(_03648_),
    .B2(_04096_),
    .Y(_04192_));
 sky130_fd_sc_hd__and3_2 _10095_ (.A(_04188_),
    .B(_03647_),
    .C(_04097_),
    .X(_04193_));
 sky130_fd_sc_hd__nand3_4 _10096_ (.A(_04188_),
    .B(_03647_),
    .C(_04097_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand3_1 _10097_ (.A(_04188_),
    .B(_04102_),
    .C(_04183_),
    .Y(_04195_));
 sky130_fd_sc_hd__a22oi_4 _10098_ (.A1(_03668_),
    .A2(_04096_),
    .B1(_04192_),
    .B2(_04194_),
    .Y(_04196_));
 sky130_fd_sc_hd__o22ai_4 _10099_ (.A1(_03669_),
    .A2(_04097_),
    .B1(_04191_),
    .B2(_04193_),
    .Y(_04198_));
 sky130_fd_sc_hd__and3_2 _10100_ (.A(_04188_),
    .B(_04098_),
    .C(_04183_),
    .X(_04199_));
 sky130_fd_sc_hd__nand3_1 _10101_ (.A(_04098_),
    .B(_04183_),
    .C(_04188_),
    .Y(_04200_));
 sky130_fd_sc_hd__and4_1 _10102_ (.A(_03640_),
    .B(_03644_),
    .C(_04096_),
    .D(_03600_),
    .X(_04201_));
 sky130_fd_sc_hd__nand4_4 _10103_ (.A(_04192_),
    .B(_04096_),
    .C(_03667_),
    .D(_03600_),
    .Y(_04202_));
 sky130_fd_sc_hd__a31o_1 _10104_ (.A1(_03668_),
    .A2(_04096_),
    .A3(_04189_),
    .B1(_04196_),
    .X(_04203_));
 sky130_fd_sc_hd__a31o_1 _10105_ (.A1(_03668_),
    .A2(_03690_),
    .A3(_03695_),
    .B1(_04113_),
    .X(_04204_));
 sky130_fd_sc_hd__a211oi_1 _10106_ (.A1(_04098_),
    .A2(_04189_),
    .B1(_04204_),
    .C1(_04196_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand4_2 _10107_ (.A(_03701_),
    .B(_04114_),
    .C(_04198_),
    .D(_04202_),
    .Y(_04206_));
 sky130_fd_sc_hd__o221a_1 _10108_ (.A1(_03690_),
    .A2(_04097_),
    .B1(_04196_),
    .B2(_04199_),
    .C1(_03698_),
    .X(_04207_));
 sky130_fd_sc_hd__o22ai_4 _10109_ (.A1(_03700_),
    .A2(_04113_),
    .B1(_04196_),
    .B2(_04199_),
    .Y(_04209_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(_04205_),
    .B(_04207_),
    .Y(_04210_));
 sky130_fd_sc_hd__and4_2 _10111_ (.A(_03700_),
    .B(_04203_),
    .C(_04108_),
    .D(_03692_),
    .X(_04211_));
 sky130_fd_sc_hd__o2111ai_4 _10112_ (.A1(_04196_),
    .A2(_04199_),
    .B1(_03692_),
    .C1(_03700_),
    .D1(_04108_),
    .Y(_04212_));
 sky130_fd_sc_hd__nand3_4 _10113_ (.A(_04118_),
    .B(_04206_),
    .C(_04209_),
    .Y(_04213_));
 sky130_fd_sc_hd__nand2_1 _10114_ (.A(_04212_),
    .B(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__o21ai_4 _10115_ (.A1(_03738_),
    .A2(_04111_),
    .B1(_04213_),
    .Y(_04215_));
 sky130_fd_sc_hd__o211a_1 _10116_ (.A1(_03738_),
    .A2(_04111_),
    .B1(_04212_),
    .C1(_04213_),
    .X(_04216_));
 sky130_fd_sc_hd__a21oi_2 _10117_ (.A1(_04212_),
    .A2(_04213_),
    .B1(_04152_),
    .Y(_04217_));
 sky130_fd_sc_hd__a21o_1 _10118_ (.A1(_04212_),
    .A2(_04213_),
    .B1(_04152_),
    .X(_04218_));
 sky130_fd_sc_hd__o21ai_1 _10119_ (.A1(_04211_),
    .A2(_04215_),
    .B1(_04218_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand2_2 _10120_ (.A(_03783_),
    .B(_04122_),
    .Y(_04221_));
 sky130_fd_sc_hd__o21ai_1 _10121_ (.A1(_03809_),
    .A2(_04122_),
    .B1(_03783_),
    .Y(_04222_));
 sky130_fd_sc_hd__o21ai_1 _10122_ (.A1(_04216_),
    .A2(_04217_),
    .B1(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__o2111ai_1 _10123_ (.A1(_03809_),
    .A2(_04122_),
    .B1(_04214_),
    .C1(_03738_),
    .D1(_03733_),
    .Y(_04224_));
 sky130_fd_sc_hd__and2_1 _10124_ (.A(_03736_),
    .B(_04122_),
    .X(_04225_));
 sky130_fd_sc_hd__o21ai_4 _10125_ (.A1(_04216_),
    .A2(_04217_),
    .B1(_04221_),
    .Y(_04226_));
 sky130_fd_sc_hd__or3_1 _10126_ (.A(_04216_),
    .B(_04217_),
    .C(_04221_),
    .X(_04227_));
 sky130_fd_sc_hd__o2111ai_4 _10127_ (.A1(_04215_),
    .A2(_04211_),
    .B1(_03736_),
    .C1(_03734_),
    .D1(_04122_),
    .Y(_04228_));
 sky130_fd_sc_hd__a21oi_4 _10128_ (.A1(_04226_),
    .A2(_04228_),
    .B1(_04127_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand4_2 _10129_ (.A(_03810_),
    .B(_04126_),
    .C(_04226_),
    .D(_04228_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(_04127_),
    .B(_04226_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_2 _10131_ (.A(_04223_),
    .B(_04224_),
    .Y(_04233_));
 sky130_fd_sc_hd__o21ai_2 _10132_ (.A1(_03823_),
    .A2(_04120_),
    .B1(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__nor2_1 _10133_ (.A(_04130_),
    .B(_04233_),
    .Y(_04235_));
 sky130_fd_sc_hd__o21ai_4 _10134_ (.A1(_04130_),
    .A2(_04229_),
    .B1(_04234_),
    .Y(_04236_));
 sky130_fd_sc_hd__a311oi_2 _10135_ (.A1(_03767_),
    .A2(_03822_),
    .A3(_04120_),
    .B1(_03835_),
    .C1(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__o211a_1 _10136_ (.A1(_03828_),
    .A2(_04120_),
    .B1(_03833_),
    .C1(_04236_),
    .X(_04238_));
 sky130_fd_sc_hd__nor2_2 _10137_ (.A(_04237_),
    .B(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__inv_2 _10138_ (.A(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__a211o_2 _10139_ (.A1(_03903_),
    .A2(_04122_),
    .B1(_03911_),
    .C1(_04239_),
    .X(_04242_));
 sky130_fd_sc_hd__o211ai_2 _10140_ (.A1(_03903_),
    .A2(_03911_),
    .B1(_04135_),
    .C1(_04239_),
    .Y(_04243_));
 sky130_fd_sc_hd__and4_1 _10141_ (.A(_04236_),
    .B(_04120_),
    .C(_03842_),
    .D(_03835_),
    .X(_04244_));
 sky130_fd_sc_hd__and2_1 _10142_ (.A(_04242_),
    .B(_04243_),
    .X(_04245_));
 sky130_fd_sc_hd__nand4_2 _10143_ (.A(_03915_),
    .B(_04131_),
    .C(_04242_),
    .D(_04243_),
    .Y(_04246_));
 sky130_fd_sc_hd__a21oi_1 _10144_ (.A1(_03915_),
    .A2(_04131_),
    .B1(_04245_),
    .Y(_04247_));
 sky130_fd_sc_hd__a22o_1 _10145_ (.A1(_04242_),
    .A2(_04243_),
    .B1(_03915_),
    .B2(_04131_),
    .X(_04248_));
 sky130_fd_sc_hd__or3b_1 _10146_ (.A(_03947_),
    .B(_04131_),
    .C_N(_04245_),
    .X(_04249_));
 sky130_fd_sc_hd__a2bb2o_1 _10147_ (.A1_N(_03947_),
    .A2_N(_04131_),
    .B1(_04246_),
    .B2(_04248_),
    .X(_04250_));
 sky130_fd_sc_hd__or4bb_1 _10148_ (.A(_03916_),
    .B(_04131_),
    .C_N(_04245_),
    .D_N(_03945_),
    .X(_04251_));
 sky130_fd_sc_hd__a21oi_2 _10149_ (.A1(net65),
    .A2(_04163_),
    .B1(_03949_),
    .Y(_04253_));
 sky130_fd_sc_hd__a31o_1 _10150_ (.A1(_03948_),
    .A2(_04250_),
    .A3(_04251_),
    .B1(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__o21ai_1 _10151_ (.A1(_02989_),
    .A2(_04151_),
    .B1(_04254_),
    .Y(net82));
 sky130_fd_sc_hd__o2bb2a_1 _10152_ (.A1_N(net49),
    .A2_N(net17),
    .B1(_01681_),
    .B2(_01692_),
    .X(_04255_));
 sky130_fd_sc_hd__and3_1 _10153_ (.A(net49),
    .B(net17),
    .C(_01703_),
    .X(_04256_));
 sky130_fd_sc_hd__or3_1 _10154_ (.A(_04145_),
    .B(_04255_),
    .C(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__o41a_1 _10155_ (.A1(_01582_),
    .A2(_01593_),
    .A3(_01703_),
    .A4(_02110_),
    .B1(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__o31a_1 _10156_ (.A1(_02132_),
    .A2(_04148_),
    .A3(_02976_),
    .B1(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__nor2_1 _10157_ (.A(_04150_),
    .B(_04258_),
    .Y(_04260_));
 sky130_fd_sc_hd__o21ba_1 _10158_ (.A1(_04259_),
    .A2(_04260_),
    .B1_N(_02996_),
    .X(_04261_));
 sky130_fd_sc_hd__nor2_1 _10159_ (.A(_04123_),
    .B(_04233_),
    .Y(_04263_));
 sky130_fd_sc_hd__or4_2 _10160_ (.A(_03768_),
    .B(_03823_),
    .C(_04122_),
    .D(_04233_),
    .X(_04264_));
 sky130_fd_sc_hd__or4b_2 _10161_ (.A(_04109_),
    .B(_03691_),
    .C(_03708_),
    .D_N(_03705_),
    .X(_04265_));
 sky130_fd_sc_hd__or3_2 _10162_ (.A(_03739_),
    .B(_04109_),
    .C(_04211_),
    .X(_04266_));
 sky130_fd_sc_hd__nor3_1 _10163_ (.A(_04114_),
    .B(_04191_),
    .C(_04193_),
    .Y(_04267_));
 sky130_fd_sc_hd__nand3_4 _10164_ (.A(_04192_),
    .B(_04194_),
    .C(_04113_),
    .Y(_04268_));
 sky130_fd_sc_hd__or3_1 _10165_ (.A(net18),
    .B(_02033_),
    .C(_02055_),
    .X(_04269_));
 sky130_fd_sc_hd__o31a_2 _10166_ (.A1(net50),
    .A2(_01989_),
    .A3(_02011_),
    .B1(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__o21ai_4 _10167_ (.A1(net50),
    .A2(_02088_),
    .B1(_04269_),
    .Y(_04271_));
 sky130_fd_sc_hd__a21oi_4 _10168_ (.A1(net99),
    .A2(_04166_),
    .B1(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__o21ai_4 _10169_ (.A1(_04167_),
    .A2(_03365_),
    .B1(_04270_),
    .Y(_04274_));
 sky130_fd_sc_hd__a221oi_2 _10170_ (.A1(net103),
    .A2(_03388_),
    .B1(net101),
    .B2(_03087_),
    .C1(_04270_),
    .Y(_04275_));
 sky130_fd_sc_hd__o2111a_2 _10171_ (.A1(_03389_),
    .A2(_04091_),
    .B1(_04165_),
    .C1(_04271_),
    .D1(net99),
    .X(_04276_));
 sky130_fd_sc_hd__o2111ai_4 _10172_ (.A1(_03389_),
    .A2(_04091_),
    .B1(_04165_),
    .C1(_04271_),
    .D1(net99),
    .Y(_04277_));
 sky130_fd_sc_hd__a21oi_4 _10173_ (.A1(_04275_),
    .A2(_04165_),
    .B1(_04272_),
    .Y(_04278_));
 sky130_fd_sc_hd__nand2_1 _10174_ (.A(_04274_),
    .B(_04277_),
    .Y(_04279_));
 sky130_fd_sc_hd__o21ai_2 _10175_ (.A1(_03425_),
    .A2(net103),
    .B1(_04178_),
    .Y(_04280_));
 sky130_fd_sc_hd__o221a_1 _10176_ (.A1(_03425_),
    .A2(net103),
    .B1(_04272_),
    .B2(_04276_),
    .C1(_04178_),
    .X(_04281_));
 sky130_fd_sc_hd__o221ai_4 _10177_ (.A1(_03425_),
    .A2(net103),
    .B1(_04272_),
    .B2(_04276_),
    .C1(_04178_),
    .Y(_04282_));
 sky130_fd_sc_hd__a21oi_1 _10178_ (.A1(_04178_),
    .A2(_04184_),
    .B1(_04279_),
    .Y(_04283_));
 sky130_fd_sc_hd__nand2_1 _10179_ (.A(_04280_),
    .B(_04278_),
    .Y(_04285_));
 sky130_fd_sc_hd__o21ai_4 _10180_ (.A1(_04272_),
    .A2(_04276_),
    .B1(_04280_),
    .Y(_04286_));
 sky130_fd_sc_hd__o211ai_4 _10181_ (.A1(_03425_),
    .A2(net103),
    .B1(_04274_),
    .C1(_04277_),
    .Y(_04287_));
 sky130_fd_sc_hd__o2111ai_4 _10182_ (.A1(_03425_),
    .A2(net103),
    .B1(_04178_),
    .C1(_04274_),
    .D1(_04277_),
    .Y(_04288_));
 sky130_fd_sc_hd__o21ai_4 _10183_ (.A1(_04177_),
    .A2(_04287_),
    .B1(_04286_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_1 _10184_ (.A(_04282_),
    .B(_04285_),
    .Y(_04290_));
 sky130_fd_sc_hd__o211a_1 _10185_ (.A1(_04177_),
    .A2(_04287_),
    .B1(_04286_),
    .C1(_04183_),
    .X(_04291_));
 sky130_fd_sc_hd__o211ai_4 _10186_ (.A1(_04177_),
    .A2(_04287_),
    .B1(_04286_),
    .C1(_04183_),
    .Y(_04292_));
 sky130_fd_sc_hd__a21oi_2 _10187_ (.A1(_04286_),
    .A2(_04288_),
    .B1(_04183_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21o_1 _10188_ (.A1(_04286_),
    .A2(_04288_),
    .B1(_04183_),
    .X(_04294_));
 sky130_fd_sc_hd__nand4_2 _10189_ (.A(_03600_),
    .B(_04096_),
    .C(_04179_),
    .D(_04289_),
    .Y(_04296_));
 sky130_fd_sc_hd__o31a_1 _10190_ (.A1(_04281_),
    .A2(_04283_),
    .A3(_04183_),
    .B1(_04292_),
    .X(_04297_));
 sky130_fd_sc_hd__nand2_1 _10191_ (.A(_04292_),
    .B(_04294_),
    .Y(_04298_));
 sky130_fd_sc_hd__o211ai_4 _10192_ (.A1(_04291_),
    .A2(_04293_),
    .B1(_04194_),
    .C1(_04200_),
    .Y(_04299_));
 sky130_fd_sc_hd__nor4b_2 _10193_ (.A(_03648_),
    .B(_04096_),
    .C(_04290_),
    .D_N(_04188_),
    .Y(_04300_));
 sky130_fd_sc_hd__nand4_4 _10194_ (.A(_04097_),
    .B(_04188_),
    .C(_04289_),
    .D(_03647_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand4_4 _10195_ (.A(_04188_),
    .B(_04098_),
    .C(_04183_),
    .D(_04292_),
    .Y(_04302_));
 sky130_fd_sc_hd__o21a_1 _10196_ (.A1(_04194_),
    .A2(_04290_),
    .B1(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__o2111ai_1 _10197_ (.A1(_04098_),
    .A2(_04105_),
    .B1(_04183_),
    .C1(_04188_),
    .D1(_04301_),
    .Y(_04304_));
 sky130_fd_sc_hd__a21oi_1 _10198_ (.A1(_04286_),
    .A2(_04288_),
    .B1(_04106_),
    .Y(_04305_));
 sky130_fd_sc_hd__o211a_1 _10199_ (.A1(_04180_),
    .A2(_04181_),
    .B1(_04188_),
    .C1(_04305_),
    .X(_04307_));
 sky130_fd_sc_hd__o21ai_2 _10200_ (.A1(_04298_),
    .A2(_04193_),
    .B1(_04304_),
    .Y(_04308_));
 sky130_fd_sc_hd__o2111a_1 _10201_ (.A1(_03648_),
    .A2(_04195_),
    .B1(_04201_),
    .C1(_04297_),
    .D1(_04192_),
    .X(_04309_));
 sky130_fd_sc_hd__nand4_4 _10202_ (.A(_04192_),
    .B(_04201_),
    .C(_04297_),
    .D(_04194_),
    .Y(_04310_));
 sky130_fd_sc_hd__and3_1 _10203_ (.A(_04297_),
    .B(_04194_),
    .C(_04201_),
    .X(_04311_));
 sky130_fd_sc_hd__nand3_4 _10204_ (.A(_04299_),
    .B(_04301_),
    .C(_04302_),
    .Y(_04312_));
 sky130_fd_sc_hd__o31ai_2 _10205_ (.A1(_04114_),
    .A2(_04191_),
    .A3(_04193_),
    .B1(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand3b_4 _10206_ (.A_N(_04268_),
    .B(_04303_),
    .C(_04299_),
    .Y(_04314_));
 sky130_fd_sc_hd__nand2_1 _10207_ (.A(_04313_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__nor3_1 _10208_ (.A(_04199_),
    .B(_03701_),
    .C(_04196_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand3_2 _10209_ (.A(_04198_),
    .B(_04202_),
    .C(_03700_),
    .Y(_04318_));
 sky130_fd_sc_hd__nand4_1 _10210_ (.A(_04198_),
    .B(_03700_),
    .C(_04109_),
    .D(_04202_),
    .Y(_04319_));
 sky130_fd_sc_hd__o2bb2ai_4 _10211_ (.A1_N(_04313_),
    .A2_N(_04314_),
    .B1(_04318_),
    .B2(_04108_),
    .Y(_04320_));
 sky130_fd_sc_hd__nor3_2 _10212_ (.A(_04115_),
    .B(_04312_),
    .C(_04318_),
    .Y(_04321_));
 sky130_fd_sc_hd__nand4b_4 _10213_ (.A_N(_04115_),
    .B(_04316_),
    .C(_04310_),
    .D(_04308_),
    .Y(_04322_));
 sky130_fd_sc_hd__o31a_1 _10214_ (.A1(_04115_),
    .A2(_04312_),
    .A3(_04318_),
    .B1(_04320_),
    .X(_04323_));
 sky130_fd_sc_hd__nand2_1 _10215_ (.A(_04320_),
    .B(_04322_),
    .Y(_04324_));
 sky130_fd_sc_hd__o2111ai_2 _10216_ (.A1(_04108_),
    .A2(_03705_),
    .B1(_03700_),
    .C1(_03692_),
    .D1(_04203_),
    .Y(_04325_));
 sky130_fd_sc_hd__a31oi_4 _10217_ (.A1(_04198_),
    .A2(_04202_),
    .A3(_04204_),
    .B1(_04118_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand3_1 _10218_ (.A(_04320_),
    .B(_04322_),
    .C(_04325_),
    .Y(_04327_));
 sky130_fd_sc_hd__a21o_1 _10219_ (.A1(_04320_),
    .A2(_04322_),
    .B1(_04325_),
    .X(_04329_));
 sky130_fd_sc_hd__and2_1 _10220_ (.A(_04327_),
    .B(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__o211ai_4 _10221_ (.A1(_04214_),
    .A2(_04265_),
    .B1(_04327_),
    .C1(_04329_),
    .Y(_04331_));
 sky130_fd_sc_hd__inv_2 _10222_ (.A(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__o2111a_1 _10223_ (.A1(_04210_),
    .A2(_03707_),
    .B1(_03738_),
    .C1(_04323_),
    .D1(_04108_),
    .X(_04333_));
 sky130_fd_sc_hd__o2111ai_4 _10224_ (.A1(_04210_),
    .A2(_03707_),
    .B1(_03738_),
    .C1(_04323_),
    .D1(_04108_),
    .Y(_04334_));
 sky130_fd_sc_hd__nand2_2 _10225_ (.A(_04331_),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__o2bb2ai_2 _10226_ (.A1_N(_04331_),
    .A2_N(_04334_),
    .B1(_04220_),
    .B2(_04221_),
    .Y(_04336_));
 sky130_fd_sc_hd__or4bb_1 _10227_ (.A(_04220_),
    .B(_04221_),
    .C_N(_04331_),
    .D_N(_04334_),
    .X(_04337_));
 sky130_fd_sc_hd__o2111a_4 _10228_ (.A1(_04211_),
    .A2(_04215_),
    .B1(_04225_),
    .C1(_03734_),
    .D1(_04331_),
    .X(_04338_));
 sky130_fd_sc_hd__o2111ai_4 _10229_ (.A1(_04211_),
    .A2(_04215_),
    .B1(_04225_),
    .C1(_03734_),
    .D1(_04331_),
    .Y(_04340_));
 sky130_fd_sc_hd__a21oi_2 _10230_ (.A1(_04228_),
    .A2(_04335_),
    .B1(_04338_),
    .Y(_04341_));
 sky130_fd_sc_hd__nand2_2 _10231_ (.A(_04336_),
    .B(_04340_),
    .Y(_04342_));
 sky130_fd_sc_hd__o31a_1 _10232_ (.A1(_03823_),
    .A2(_04120_),
    .A3(_04233_),
    .B1(_04231_),
    .X(_04343_));
 sky130_fd_sc_hd__o21ai_1 _10233_ (.A1(_04130_),
    .A2(_04233_),
    .B1(_04231_),
    .Y(_04344_));
 sky130_fd_sc_hd__o211ai_2 _10234_ (.A1(_04130_),
    .A2(_04229_),
    .B1(_04231_),
    .C1(_04341_),
    .Y(_04345_));
 sky130_fd_sc_hd__nand2_1 _10235_ (.A(_04342_),
    .B(_04344_),
    .Y(_04346_));
 sky130_fd_sc_hd__a22oi_2 _10236_ (.A1(_04127_),
    .A2(_04226_),
    .B1(_04336_),
    .B2(_04340_),
    .Y(_04347_));
 sky130_fd_sc_hd__nor4_2 _10237_ (.A(_03823_),
    .B(_04120_),
    .C(_04229_),
    .D(_04342_),
    .Y(_04348_));
 sky130_fd_sc_hd__or4_1 _10238_ (.A(_03823_),
    .B(_04120_),
    .C(_04229_),
    .D(_04342_),
    .X(_04349_));
 sky130_fd_sc_hd__a21oi_4 _10239_ (.A1(_04228_),
    .A2(_04335_),
    .B1(_04232_),
    .Y(_04351_));
 sky130_fd_sc_hd__a21o_2 _10240_ (.A1(_04228_),
    .A2(_04335_),
    .B1(_04232_),
    .X(_04352_));
 sky130_fd_sc_hd__o22a_2 _10241_ (.A1(_04229_),
    .A2(_04130_),
    .B1(_04351_),
    .B2(_04347_),
    .X(_04353_));
 sky130_fd_sc_hd__o22ai_2 _10242_ (.A1(_04229_),
    .A2(_04130_),
    .B1(_04351_),
    .B2(_04347_),
    .Y(_04354_));
 sky130_fd_sc_hd__nand3b_4 _10243_ (.A_N(_04263_),
    .B(_04345_),
    .C(_04346_),
    .Y(_04355_));
 sky130_fd_sc_hd__nand2_4 _10244_ (.A(_04354_),
    .B(_04263_),
    .Y(_04356_));
 sky130_fd_sc_hd__o21ai_2 _10245_ (.A1(_04264_),
    .A2(_04353_),
    .B1(_04355_),
    .Y(_04357_));
 sky130_fd_sc_hd__o2111a_2 _10246_ (.A1(_03823_),
    .A2(_04229_),
    .B1(_04234_),
    .C1(_04122_),
    .D1(_03835_),
    .X(_04358_));
 sky130_fd_sc_hd__a2bb2oi_2 _10247_ (.A1_N(_04134_),
    .A2_N(_04236_),
    .B1(_04355_),
    .B2(_04356_),
    .Y(_04359_));
 sky130_fd_sc_hd__o311a_2 _10248_ (.A1(_04123_),
    .A2(_04236_),
    .A3(_04353_),
    .B1(_04355_),
    .C1(_04358_),
    .X(_04360_));
 sky130_fd_sc_hd__nand2_2 _10249_ (.A(_04355_),
    .B(_04358_),
    .Y(_04362_));
 sky130_fd_sc_hd__a21oi_4 _10250_ (.A1(_04355_),
    .A2(_04358_),
    .B1(_04359_),
    .Y(_04363_));
 sky130_fd_sc_hd__xor2_2 _10251_ (.A(_04242_),
    .B(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__and4b_1 _10252_ (.A_N(_04141_),
    .B(_04242_),
    .C(_04243_),
    .D(_04363_),
    .X(_04365_));
 sky130_fd_sc_hd__o311a_1 _10253_ (.A1(_03947_),
    .A2(_04131_),
    .A3(_04247_),
    .B1(_04364_),
    .C1(_04246_),
    .X(_04366_));
 sky130_fd_sc_hd__a21oi_1 _10254_ (.A1(_04246_),
    .A2(_04249_),
    .B1(_04364_),
    .Y(_04367_));
 sky130_fd_sc_hd__or2_1 _10255_ (.A(_04366_),
    .B(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__mux2_1 _10256_ (.A0(_04270_),
    .A1(_04368_),
    .S(_03948_),
    .X(_04369_));
 sky130_fd_sc_hd__a2bb2o_1 _10257_ (.A1_N(_04261_),
    .A2_N(_02989_),
    .B1(net65),
    .B2(_04369_),
    .X(net83));
 sky130_fd_sc_hd__or3b_1 _10258_ (.A(_01648_),
    .B(_01659_),
    .C_N(_01692_),
    .X(_04370_));
 sky130_fd_sc_hd__a2bb2o_1 _10259_ (.A1_N(_01648_),
    .A2_N(_01659_),
    .B1(net50),
    .B2(net18),
    .X(_04372_));
 sky130_fd_sc_hd__nand2_1 _10260_ (.A(_04370_),
    .B(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__o21bai_1 _10261_ (.A1(_04146_),
    .A2(_04255_),
    .B1_N(_04256_),
    .Y(_04374_));
 sky130_fd_sc_hd__xor2_1 _10262_ (.A(_04373_),
    .B(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__a21oi_1 _10263_ (.A1(_04260_),
    .A2(_04375_),
    .B1(_02996_),
    .Y(_04376_));
 sky130_fd_sc_hd__o21a_1 _10264_ (.A1(_04260_),
    .A2(_04375_),
    .B1(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__nand2_4 _10265_ (.A(_04244_),
    .B(_04363_),
    .Y(_04378_));
 sky130_fd_sc_hd__and3_1 _10266_ (.A(_04168_),
    .B(_04169_),
    .C(_04271_),
    .X(_04379_));
 sky130_fd_sc_hd__o21ai_4 _10267_ (.A1(_04170_),
    .A2(_04172_),
    .B1(_04271_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand4_1 _10268_ (.A(net99),
    .B(_03401_),
    .C(_04091_),
    .D(_04163_),
    .Y(_04381_));
 sky130_fd_sc_hd__nor2_2 _10269_ (.A(_04270_),
    .B(_04381_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21a_2 _10270_ (.A1(_04159_),
    .A2(_04160_),
    .B1(_04271_),
    .X(_04384_));
 sky130_fd_sc_hd__a311o_1 _10271_ (.A1(net49),
    .A2(_02000_),
    .A3(_02022_),
    .B1(_04161_),
    .C1(_04270_),
    .X(_04385_));
 sky130_fd_sc_hd__and3_1 _10272_ (.A(net103),
    .B(_04165_),
    .C(_04271_),
    .X(_04386_));
 sky130_fd_sc_hd__nand4_4 _10273_ (.A(net99),
    .B(_03389_),
    .C(net103),
    .D(_04384_),
    .Y(_04387_));
 sky130_fd_sc_hd__and3_1 _10274_ (.A(_00988_),
    .B(_02044_),
    .C(_02066_),
    .X(_04388_));
 sky130_fd_sc_hd__a21oi_1 _10275_ (.A1(_02044_),
    .A2(_02066_),
    .B1(net51),
    .Y(_04389_));
 sky130_fd_sc_hd__and3_1 _10276_ (.A(_02066_),
    .B(net19),
    .C(_02044_),
    .X(_04390_));
 sky130_fd_sc_hd__and3_1 _10277_ (.A(_02022_),
    .B(net51),
    .C(_02000_),
    .X(_04391_));
 sky130_fd_sc_hd__a31o_1 _10278_ (.A1(net51),
    .A2(_02000_),
    .A3(_02022_),
    .B1(_04390_),
    .X(_04392_));
 sky130_fd_sc_hd__a31o_2 _10279_ (.A1(_00988_),
    .A2(_02044_),
    .A3(_02066_),
    .B1(_04389_),
    .X(_04394_));
 sky130_fd_sc_hd__and3_1 _10280_ (.A(_04271_),
    .B(_04091_),
    .C(_04165_),
    .X(_04395_));
 sky130_fd_sc_hd__or4_1 _10281_ (.A(_04092_),
    .B(_04161_),
    .C(_04162_),
    .D(_04270_),
    .X(_04396_));
 sky130_fd_sc_hd__o22a_2 _10282_ (.A1(_04390_),
    .A2(_04391_),
    .B1(_04396_),
    .B2(_03365_),
    .X(_04397_));
 sky130_fd_sc_hd__o22ai_1 _10283_ (.A1(_04390_),
    .A2(_04391_),
    .B1(_04396_),
    .B2(_03365_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand4_1 _10284_ (.A(net99),
    .B(_04091_),
    .C(_04384_),
    .D(_04394_),
    .Y(_04399_));
 sky130_fd_sc_hd__o22ai_2 _10285_ (.A1(_04388_),
    .A2(_04389_),
    .B1(_04396_),
    .B2(_03365_),
    .Y(_04400_));
 sky130_fd_sc_hd__o211ai_2 _10286_ (.A1(_04390_),
    .A2(_04391_),
    .B1(_04395_),
    .C1(net99),
    .Y(_04401_));
 sky130_fd_sc_hd__nor4_2 _10287_ (.A(_04091_),
    .B(_04385_),
    .C(_04392_),
    .D(_03404_),
    .Y(_04402_));
 sky130_fd_sc_hd__nand4_2 _10288_ (.A(_03403_),
    .B(net103),
    .C(_04384_),
    .D(_04394_),
    .Y(_04403_));
 sky130_fd_sc_hd__a22oi_1 _10289_ (.A1(_03403_),
    .A2(_04386_),
    .B1(_04398_),
    .B2(_04399_),
    .Y(_04405_));
 sky130_fd_sc_hd__nand3_4 _10290_ (.A(_04387_),
    .B(_04400_),
    .C(_04401_),
    .Y(_04406_));
 sky130_fd_sc_hd__o41a_2 _10291_ (.A1(_04091_),
    .A2(_04385_),
    .A3(_04392_),
    .A4(_03404_),
    .B1(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__o21ai_4 _10292_ (.A1(_04387_),
    .A2(_04397_),
    .B1(_04406_),
    .Y(_04408_));
 sky130_fd_sc_hd__o211a_1 _10293_ (.A1(_04387_),
    .A2(_04397_),
    .B1(_04383_),
    .C1(_04406_),
    .X(_04409_));
 sky130_fd_sc_hd__o211ai_4 _10294_ (.A1(_04387_),
    .A2(_04397_),
    .B1(_04383_),
    .C1(_04406_),
    .Y(_04410_));
 sky130_fd_sc_hd__a21oi_2 _10295_ (.A1(_04403_),
    .A2(_04406_),
    .B1(_04383_),
    .Y(_04411_));
 sky130_fd_sc_hd__o21bai_1 _10296_ (.A1(_04402_),
    .A2(_04405_),
    .B1_N(_04383_),
    .Y(_04412_));
 sky130_fd_sc_hd__and4_1 _10297_ (.A(_04169_),
    .B(_03408_),
    .C(_04168_),
    .D(_04271_),
    .X(_04413_));
 sky130_fd_sc_hd__a22oi_4 _10298_ (.A1(net103),
    .A2(_04413_),
    .B1(_04412_),
    .B2(_04410_),
    .Y(_04414_));
 sky130_fd_sc_hd__o22ai_4 _10299_ (.A1(_04095_),
    .A2(_04380_),
    .B1(_04409_),
    .B2(_04411_),
    .Y(_04416_));
 sky130_fd_sc_hd__nor4_4 _10300_ (.A(_03409_),
    .B(_04091_),
    .C(_04380_),
    .D(_04408_),
    .Y(_04417_));
 sky130_fd_sc_hd__nand4_4 _10301_ (.A(_03408_),
    .B(_04407_),
    .C(net103),
    .D(_04379_),
    .Y(_04418_));
 sky130_fd_sc_hd__o31a_1 _10302_ (.A1(_04095_),
    .A2(_04380_),
    .A3(_04411_),
    .B1(_04416_),
    .X(_04419_));
 sky130_fd_sc_hd__nand2_4 _10303_ (.A(_04416_),
    .B(_04418_),
    .Y(_04420_));
 sky130_fd_sc_hd__and3_2 _10304_ (.A(_04187_),
    .B(_04274_),
    .C(_04277_),
    .X(_04421_));
 sky130_fd_sc_hd__a22oi_4 _10305_ (.A1(_04187_),
    .A2(_04278_),
    .B1(_04289_),
    .B2(_04182_),
    .Y(_04422_));
 sky130_fd_sc_hd__and4b_2 _10306_ (.A_N(_04184_),
    .B(_04278_),
    .C(_04176_),
    .D(_04178_),
    .X(_04423_));
 sky130_fd_sc_hd__o2111ai_4 _10307_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_04179_),
    .C1(_04278_),
    .D1(_03424_),
    .Y(_04424_));
 sky130_fd_sc_hd__o21ai_4 _10308_ (.A1(_04414_),
    .A2(_04417_),
    .B1(_04422_),
    .Y(_04425_));
 sky130_fd_sc_hd__o211ai_1 _10309_ (.A1(_04293_),
    .A2(_04421_),
    .B1(_04418_),
    .C1(_04416_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand3_2 _10310_ (.A(_04422_),
    .B(_04418_),
    .C(_04416_),
    .Y(_04428_));
 sky130_fd_sc_hd__o2bb2ai_2 _10311_ (.A1_N(_04416_),
    .A2_N(_04418_),
    .B1(_04421_),
    .B2(_04293_),
    .Y(_04429_));
 sky130_fd_sc_hd__a31oi_2 _10312_ (.A1(_04182_),
    .A2(_04282_),
    .A3(_04285_),
    .B1(_04423_),
    .Y(_04430_));
 sky130_fd_sc_hd__a21oi_1 _10313_ (.A1(_04427_),
    .A2(_04425_),
    .B1(_04300_),
    .Y(_04431_));
 sky130_fd_sc_hd__nand3_4 _10314_ (.A(_04301_),
    .B(_04428_),
    .C(_04429_),
    .Y(_04432_));
 sky130_fd_sc_hd__o211ai_4 _10315_ (.A1(_04430_),
    .A2(_04420_),
    .B1(_04300_),
    .C1(_04425_),
    .Y(_04433_));
 sky130_fd_sc_hd__and3_2 _10316_ (.A(_04425_),
    .B(_04305_),
    .C(_04189_),
    .X(_04434_));
 sky130_fd_sc_hd__nand2_1 _10317_ (.A(_04425_),
    .B(_04307_),
    .Y(_04435_));
 sky130_fd_sc_hd__o2bb2ai_2 _10318_ (.A1_N(_04302_),
    .A2_N(_04314_),
    .B1(_04431_),
    .B2(_04434_),
    .Y(_04436_));
 sky130_fd_sc_hd__o2111ai_4 _10319_ (.A1(_04268_),
    .A2(_04312_),
    .B1(_04432_),
    .C1(_04433_),
    .D1(_04302_),
    .Y(_04438_));
 sky130_fd_sc_hd__nand3b_1 _10320_ (.A_N(_04314_),
    .B(_04432_),
    .C(_04433_),
    .Y(_04439_));
 sky130_fd_sc_hd__a21oi_1 _10321_ (.A1(_04432_),
    .A2(_04435_),
    .B1(_04309_),
    .Y(_04440_));
 sky130_fd_sc_hd__o211a_1 _10322_ (.A1(_04105_),
    .A2(_04189_),
    .B1(_04311_),
    .C1(_04432_),
    .X(_04441_));
 sky130_fd_sc_hd__o211ai_2 _10323_ (.A1(_04105_),
    .A2(_04189_),
    .B1(_04311_),
    .C1(_04432_),
    .Y(_04442_));
 sky130_fd_sc_hd__o22ai_4 _10324_ (.A1(_04268_),
    .A2(_04312_),
    .B1(_04440_),
    .B2(_04441_),
    .Y(_04443_));
 sky130_fd_sc_hd__and4_2 _10325_ (.A(_04308_),
    .B(_04432_),
    .C(_04267_),
    .D(_04433_),
    .X(_04444_));
 sky130_fd_sc_hd__nand4_2 _10326_ (.A(_04308_),
    .B(_04432_),
    .C(_04267_),
    .D(_04433_),
    .Y(_04445_));
 sky130_fd_sc_hd__nand2_1 _10327_ (.A(_04436_),
    .B(_04438_),
    .Y(_04446_));
 sky130_fd_sc_hd__inv_2 _10328_ (.A(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__nand3_4 _10329_ (.A(_04322_),
    .B(_04436_),
    .C(_04438_),
    .Y(_04449_));
 sky130_fd_sc_hd__a21oi_2 _10330_ (.A1(_04436_),
    .A2(_04438_),
    .B1(_04322_),
    .Y(_04450_));
 sky130_fd_sc_hd__nand3_4 _10331_ (.A(_04443_),
    .B(_04445_),
    .C(_04321_),
    .Y(_04451_));
 sky130_fd_sc_hd__a21boi_2 _10332_ (.A1(_04315_),
    .A2(_04319_),
    .B1_N(_04326_),
    .Y(_04452_));
 sky130_fd_sc_hd__a22oi_4 _10333_ (.A1(_04326_),
    .A2(_04320_),
    .B1(_04451_),
    .B2(_04449_),
    .Y(_04453_));
 sky130_fd_sc_hd__o2bb2ai_2 _10334_ (.A1_N(_04449_),
    .A2_N(_04451_),
    .B1(_04212_),
    .B2(_04324_),
    .Y(_04454_));
 sky130_fd_sc_hd__and3_1 _10335_ (.A(_04320_),
    .B(_04449_),
    .C(_04326_),
    .X(_04455_));
 sky130_fd_sc_hd__nand2_2 _10336_ (.A(_04449_),
    .B(_04452_),
    .Y(_04456_));
 sky130_fd_sc_hd__a211o_1 _10337_ (.A1(_04206_),
    .A2(_04209_),
    .B1(_04324_),
    .C1(_04112_),
    .X(_04457_));
 sky130_fd_sc_hd__o2111a_1 _10338_ (.A1(_04205_),
    .A2(_04207_),
    .B1(_04322_),
    .C1(_04111_),
    .D1(_04320_),
    .X(_04458_));
 sky130_fd_sc_hd__and4_1 _10339_ (.A(_04213_),
    .B(_04320_),
    .C(_04322_),
    .D(_04111_),
    .X(_04460_));
 sky130_fd_sc_hd__nand4_2 _10340_ (.A(_04320_),
    .B(_04111_),
    .C(_04213_),
    .D(_04322_),
    .Y(_04461_));
 sky130_fd_sc_hd__a21oi_4 _10341_ (.A1(_04454_),
    .A2(_04456_),
    .B1(_04460_),
    .Y(_04462_));
 sky130_fd_sc_hd__o21ai_2 _10342_ (.A1(_04453_),
    .A2(_04455_),
    .B1(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__a311oi_2 _10343_ (.A1(_04320_),
    .A2(_04326_),
    .A3(_04449_),
    .B1(_04453_),
    .C1(_04457_),
    .Y(_04464_));
 sky130_fd_sc_hd__nor2_1 _10344_ (.A(_04461_),
    .B(_04453_),
    .Y(_04465_));
 sky130_fd_sc_hd__a2111o_2 _10345_ (.A1(_04118_),
    .A2(_04210_),
    .B1(_04324_),
    .C1(_04112_),
    .D1(_04453_),
    .X(_04466_));
 sky130_fd_sc_hd__o21ai_1 _10346_ (.A1(_04453_),
    .A2(_04461_),
    .B1(_04463_),
    .Y(_04467_));
 sky130_fd_sc_hd__o22a_2 _10347_ (.A1(_04330_),
    .A2(_04266_),
    .B1(_04465_),
    .B2(_04462_),
    .X(_04468_));
 sky130_fd_sc_hd__o22ai_4 _10348_ (.A1(_04330_),
    .A2(_04266_),
    .B1(_04465_),
    .B2(_04462_),
    .Y(_04469_));
 sky130_fd_sc_hd__nor2_2 _10349_ (.A(_04334_),
    .B(_04462_),
    .Y(_04471_));
 sky130_fd_sc_hd__nand2_1 _10350_ (.A(_04463_),
    .B(_04333_),
    .Y(_04472_));
 sky130_fd_sc_hd__o31a_1 _10351_ (.A1(_04266_),
    .A2(_04330_),
    .A3(_04462_),
    .B1(_04469_),
    .X(_04473_));
 sky130_fd_sc_hd__o21ai_1 _10352_ (.A1(_04334_),
    .A2(_04462_),
    .B1(_04469_),
    .Y(_04474_));
 sky130_fd_sc_hd__a21oi_1 _10353_ (.A1(_04469_),
    .A2(_04472_),
    .B1(_04338_),
    .Y(_04475_));
 sky130_fd_sc_hd__o22ai_4 _10354_ (.A1(_04332_),
    .A2(_04228_),
    .B1(_04471_),
    .B2(_04468_),
    .Y(_04476_));
 sky130_fd_sc_hd__nor4_1 _10355_ (.A(_04227_),
    .B(_04332_),
    .C(_04333_),
    .D(_04467_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_4 _10356_ (.A(_04469_),
    .B(_04338_),
    .Y(_04478_));
 sky130_fd_sc_hd__o31a_1 _10357_ (.A1(_04228_),
    .A2(_04332_),
    .A3(_04468_),
    .B1(_04476_),
    .X(_04479_));
 sky130_fd_sc_hd__o21ai_1 _10358_ (.A1(_04340_),
    .A2(_04468_),
    .B1(_04476_),
    .Y(_04480_));
 sky130_fd_sc_hd__o211ai_4 _10359_ (.A1(_04342_),
    .A2(_04343_),
    .B1(_04476_),
    .C1(_04478_),
    .Y(_04482_));
 sky130_fd_sc_hd__nand4_2 _10360_ (.A(_04336_),
    .B(_04340_),
    .C(_04344_),
    .D(_04474_),
    .Y(_04483_));
 sky130_fd_sc_hd__o41ai_2 _10361_ (.A1(_03823_),
    .A2(_04120_),
    .A3(_04229_),
    .A4(_04342_),
    .B1(_04352_),
    .Y(_04484_));
 sky130_fd_sc_hd__a21oi_4 _10362_ (.A1(_04476_),
    .A2(_04478_),
    .B1(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__and3_2 _10363_ (.A(_04356_),
    .B(_04482_),
    .C(_04483_),
    .X(_04486_));
 sky130_fd_sc_hd__o211ai_2 _10364_ (.A1(_04353_),
    .A2(_04264_),
    .B1(_04483_),
    .C1(_04482_),
    .Y(_04487_));
 sky130_fd_sc_hd__a21oi_2 _10365_ (.A1(_04482_),
    .A2(_04483_),
    .B1(_04356_),
    .Y(_04488_));
 sky130_fd_sc_hd__a31o_2 _10366_ (.A1(_04349_),
    .A2(_04352_),
    .A3(_04480_),
    .B1(_04356_),
    .X(_04489_));
 sky130_fd_sc_hd__o31a_2 _10367_ (.A1(_04264_),
    .A2(_04353_),
    .A3(_04485_),
    .B1(_04487_),
    .X(_04490_));
 sky130_fd_sc_hd__o21ai_1 _10368_ (.A1(_04356_),
    .A2(_04485_),
    .B1(_04487_),
    .Y(_04491_));
 sky130_fd_sc_hd__o32a_1 _10369_ (.A1(_04134_),
    .A2(_04236_),
    .A3(_04357_),
    .B1(_04486_),
    .B2(_04488_),
    .X(_04493_));
 sky130_fd_sc_hd__o31ai_4 _10370_ (.A1(_04134_),
    .A2(_04236_),
    .A3(_04357_),
    .B1(_04491_),
    .Y(_04494_));
 sky130_fd_sc_hd__o311a_1 _10371_ (.A1(_04264_),
    .A2(_04353_),
    .A3(_04485_),
    .B1(_04487_),
    .C1(_04360_),
    .X(_04495_));
 sky130_fd_sc_hd__a31o_2 _10372_ (.A1(_04356_),
    .A2(_04482_),
    .A3(_04483_),
    .B1(_04362_),
    .X(_04496_));
 sky130_fd_sc_hd__inv_2 _10373_ (.A(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__o21a_1 _10374_ (.A1(_04362_),
    .A2(_04486_),
    .B1(_04494_),
    .X(_04498_));
 sky130_fd_sc_hd__o21ai_4 _10375_ (.A1(_04362_),
    .A2(_04486_),
    .B1(_04494_),
    .Y(_04499_));
 sky130_fd_sc_hd__nor4_2 _10376_ (.A(_03911_),
    .B(_04122_),
    .C(_04357_),
    .D(_04239_),
    .Y(_04500_));
 sky130_fd_sc_hd__nand3_1 _10377_ (.A(_04378_),
    .B(_04494_),
    .C(_04496_),
    .Y(_04501_));
 sky130_fd_sc_hd__o21ai_1 _10378_ (.A1(_04486_),
    .A2(_04488_),
    .B1(_04500_),
    .Y(_04502_));
 sky130_fd_sc_hd__a22oi_2 _10379_ (.A1(_04244_),
    .A2(_04363_),
    .B1(_04494_),
    .B2(_04496_),
    .Y(_04504_));
 sky130_fd_sc_hd__o21ai_1 _10380_ (.A1(_04500_),
    .A2(_04499_),
    .B1(_04502_),
    .Y(_04505_));
 sky130_fd_sc_hd__o211ai_1 _10381_ (.A1(_04237_),
    .A2(_04238_),
    .B1(_04363_),
    .C1(_04136_),
    .Y(_04506_));
 sky130_fd_sc_hd__or3_2 _10382_ (.A(_04239_),
    .B(_04359_),
    .C(_04139_),
    .X(_04507_));
 sky130_fd_sc_hd__o211ai_2 _10383_ (.A1(_04378_),
    .A2(_04490_),
    .B1(_04501_),
    .C1(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__a21oi_1 _10384_ (.A1(_04501_),
    .A2(_04502_),
    .B1(_04506_),
    .Y(_04509_));
 sky130_fd_sc_hd__a21o_1 _10385_ (.A1(_04501_),
    .A2(_04502_),
    .B1(_04506_),
    .X(_04510_));
 sky130_fd_sc_hd__and4_1 _10386_ (.A(_04240_),
    .B(_04505_),
    .C(_04363_),
    .D(_04136_),
    .X(_04511_));
 sky130_fd_sc_hd__a21oi_2 _10387_ (.A1(_04378_),
    .A2(_04499_),
    .B1(_04507_),
    .Y(_04512_));
 sky130_fd_sc_hd__o41a_2 _10388_ (.A1(_04139_),
    .A2(_04239_),
    .A3(_04359_),
    .A4(_04504_),
    .B1(_04508_),
    .X(_04513_));
 sky130_fd_sc_hd__o21ai_1 _10389_ (.A1(_04504_),
    .A2(_04507_),
    .B1(_04508_),
    .Y(_04515_));
 sky130_fd_sc_hd__o21ai_1 _10390_ (.A1(_04367_),
    .A2(_04513_),
    .B1(_03948_),
    .Y(_04516_));
 sky130_fd_sc_hd__a21o_1 _10391_ (.A1(_04367_),
    .A2(_04513_),
    .B1(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__o31a_1 _10392_ (.A1(_03573_),
    .A2(_03947_),
    .A3(_04392_),
    .B1(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__a2bb2o_1 _10393_ (.A1_N(_02989_),
    .A2_N(_04377_),
    .B1(_04518_),
    .B2(net65),
    .X(net84));
 sky130_fd_sc_hd__or4_1 _10394_ (.A(_04255_),
    .B(_04256_),
    .C(_04373_),
    .D(_04148_),
    .X(_04519_));
 sky130_fd_sc_hd__a21boi_1 _10395_ (.A1(_04372_),
    .A2(_04374_),
    .B1_N(_04370_),
    .Y(_04520_));
 sky130_fd_sc_hd__and3_1 _10396_ (.A(_01791_),
    .B(_01802_),
    .C(_01659_),
    .X(_04521_));
 sky130_fd_sc_hd__a21oi_1 _10397_ (.A1(_01791_),
    .A2(_01802_),
    .B1(_01659_),
    .Y(_04522_));
 sky130_fd_sc_hd__nor3_1 _10398_ (.A(_04520_),
    .B(_04521_),
    .C(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__o21a_1 _10399_ (.A1(_04521_),
    .A2(_04522_),
    .B1(_04520_),
    .X(_04525_));
 sky130_fd_sc_hd__or2_1 _10400_ (.A(_04523_),
    .B(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__o21ai_1 _10401_ (.A1(_04086_),
    .A2(_04519_),
    .B1(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__or4_1 _10402_ (.A(_02132_),
    .B(_04519_),
    .C(_04526_),
    .D(_02976_),
    .X(_04528_));
 sky130_fd_sc_hd__a21oi_1 _10403_ (.A1(_04527_),
    .A2(_04528_),
    .B1(_02996_),
    .Y(_04529_));
 sky130_fd_sc_hd__o211ai_4 _10404_ (.A1(_04170_),
    .A2(_04172_),
    .B1(_04271_),
    .C1(_04156_),
    .Y(_04530_));
 sky130_fd_sc_hd__or3_1 _10405_ (.A(net20),
    .B(_02033_),
    .C(_02055_),
    .X(_04531_));
 sky130_fd_sc_hd__o31a_1 _10406_ (.A1(net52),
    .A2(_01989_),
    .A3(_02011_),
    .B1(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__o21ai_4 _10407_ (.A1(net52),
    .A2(_02088_),
    .B1(_04531_),
    .Y(_04533_));
 sky130_fd_sc_hd__a31oi_4 _10408_ (.A1(_04158_),
    .A2(_04384_),
    .A3(_04394_),
    .B1(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__a31o_1 _10409_ (.A1(_04158_),
    .A2(_04384_),
    .A3(_04394_),
    .B1(_04533_),
    .X(_04536_));
 sky130_fd_sc_hd__and4_1 _10410_ (.A(_04158_),
    .B(_04384_),
    .C(_04394_),
    .D(_04533_),
    .X(_04537_));
 sky130_fd_sc_hd__nand4_1 _10411_ (.A(_04158_),
    .B(_04384_),
    .C(_04394_),
    .D(_04533_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_2 _10412_ (.A(_04536_),
    .B(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_2 _10413_ (.A(_04534_),
    .B(_04537_),
    .Y(_04540_));
 sky130_fd_sc_hd__o21ai_1 _10414_ (.A1(_04408_),
    .A2(_04530_),
    .B1(_04539_),
    .Y(_04541_));
 sky130_fd_sc_hd__o21ai_1 _10415_ (.A1(_04408_),
    .A2(_04530_),
    .B1(_04540_),
    .Y(_04542_));
 sky130_fd_sc_hd__nand4_1 _10416_ (.A(_04407_),
    .B(_04156_),
    .C(_04379_),
    .D(_04539_),
    .Y(_04543_));
 sky130_fd_sc_hd__nand2_2 _10417_ (.A(_04542_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__o41ai_4 _10418_ (.A1(_04534_),
    .A2(_04537_),
    .A3(_04408_),
    .A4(_04530_),
    .B1(_04541_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand3_1 _10419_ (.A(_04416_),
    .B(_04418_),
    .C(_04423_),
    .Y(_04547_));
 sky130_fd_sc_hd__a21oi_4 _10420_ (.A1(_04416_),
    .A2(_04423_),
    .B1(_04544_),
    .Y(_04548_));
 sky130_fd_sc_hd__o21ai_4 _10421_ (.A1(_04424_),
    .A2(_04414_),
    .B1(_04545_),
    .Y(_04549_));
 sky130_fd_sc_hd__nand4_4 _10422_ (.A(_04544_),
    .B(_04418_),
    .C(_04416_),
    .D(_04421_),
    .Y(_04550_));
 sky130_fd_sc_hd__nor2_1 _10423_ (.A(_04296_),
    .B(_04420_),
    .Y(_04551_));
 sky130_fd_sc_hd__nand3b_4 _10424_ (.A_N(_04296_),
    .B(_04416_),
    .C(_04418_),
    .Y(_04552_));
 sky130_fd_sc_hd__o2bb2ai_4 _10425_ (.A1_N(_04549_),
    .A2_N(_04550_),
    .B1(_04294_),
    .B2(_04420_),
    .Y(_04553_));
 sky130_fd_sc_hd__and4_1 _10426_ (.A(_04550_),
    .B(_04293_),
    .C(_04549_),
    .D(_04419_),
    .X(_04554_));
 sky130_fd_sc_hd__a211o_2 _10427_ (.A1(_04424_),
    .A2(_04545_),
    .B1(_04296_),
    .C1(_04420_),
    .X(_04555_));
 sky130_fd_sc_hd__o31a_2 _10428_ (.A1(_04296_),
    .A2(_04420_),
    .A3(_04548_),
    .B1(_04553_),
    .X(_04556_));
 sky130_fd_sc_hd__o21ai_4 _10429_ (.A1(_04548_),
    .A2(_04552_),
    .B1(_04553_),
    .Y(_04558_));
 sky130_fd_sc_hd__o41ai_2 _10430_ (.A1(_03669_),
    .A2(_04097_),
    .A3(_04190_),
    .A4(_04298_),
    .B1(_04433_),
    .Y(_04559_));
 sky130_fd_sc_hd__o211ai_2 _10431_ (.A1(_04302_),
    .A2(_04431_),
    .B1(_04433_),
    .C1(_04558_),
    .Y(_04560_));
 sky130_fd_sc_hd__o2111ai_4 _10432_ (.A1(_04548_),
    .A2(_04552_),
    .B1(_04553_),
    .C1(_04559_),
    .D1(_04432_),
    .Y(_04561_));
 sky130_fd_sc_hd__a31oi_4 _10433_ (.A1(_04301_),
    .A2(_04428_),
    .A3(_04429_),
    .B1(_04310_),
    .Y(_04562_));
 sky130_fd_sc_hd__nand4_4 _10434_ (.A(_04435_),
    .B(_04442_),
    .C(_04553_),
    .D(_04555_),
    .Y(_04563_));
 sky130_fd_sc_hd__o21ai_2 _10435_ (.A1(_04434_),
    .A2(_04562_),
    .B1(_04558_),
    .Y(_04564_));
 sky130_fd_sc_hd__nand2_2 _10436_ (.A(_04563_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__inv_2 _10437_ (.A(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__a21oi_1 _10438_ (.A1(_04560_),
    .A2(_04561_),
    .B1(_04444_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand3_1 _10439_ (.A(_04445_),
    .B(_04563_),
    .C(_04564_),
    .Y(_04569_));
 sky130_fd_sc_hd__a21oi_2 _10440_ (.A1(_04563_),
    .A2(_04564_),
    .B1(_04439_),
    .Y(_04570_));
 sky130_fd_sc_hd__a21o_1 _10441_ (.A1(_04563_),
    .A2(_04564_),
    .B1(_04439_),
    .X(_04571_));
 sky130_fd_sc_hd__nand3_2 _10442_ (.A(_04561_),
    .B(_04444_),
    .C(_04560_),
    .Y(_04572_));
 sky130_fd_sc_hd__a31o_1 _10443_ (.A1(_04445_),
    .A2(_04563_),
    .A3(_04564_),
    .B1(_04570_),
    .X(_04573_));
 sky130_fd_sc_hd__a22oi_1 _10444_ (.A1(_04569_),
    .A2(_04572_),
    .B1(_04449_),
    .B2(_04452_),
    .Y(_04574_));
 sky130_fd_sc_hd__o2bb2ai_1 _10445_ (.A1_N(_04449_),
    .A2_N(_04452_),
    .B1(_04567_),
    .B2(_04570_),
    .Y(_04575_));
 sky130_fd_sc_hd__and4_2 _10446_ (.A(_04449_),
    .B(_04452_),
    .C(_04569_),
    .D(_04572_),
    .X(_04576_));
 sky130_fd_sc_hd__nand4_1 _10447_ (.A(_04449_),
    .B(_04452_),
    .C(_04569_),
    .D(_04572_),
    .Y(_04577_));
 sky130_fd_sc_hd__nand2_1 _10448_ (.A(_04575_),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__a21oi_1 _10449_ (.A1(_04575_),
    .A2(_04577_),
    .B1(_04450_),
    .Y(_04580_));
 sky130_fd_sc_hd__o22ai_2 _10450_ (.A1(_04322_),
    .A2(_04447_),
    .B1(_04574_),
    .B2(_04576_),
    .Y(_04581_));
 sky130_fd_sc_hd__and3_1 _10451_ (.A(_04446_),
    .B(_04565_),
    .C(_04321_),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_1 _10452_ (.A(_04450_),
    .B(_04565_),
    .Y(_04583_));
 sky130_fd_sc_hd__and3_1 _10453_ (.A(_04321_),
    .B(_04560_),
    .C(_04561_),
    .X(_04584_));
 sky130_fd_sc_hd__a22oi_4 _10454_ (.A1(_04443_),
    .A2(_04584_),
    .B1(_04578_),
    .B2(_04451_),
    .Y(_04585_));
 sky130_fd_sc_hd__o21ai_2 _10455_ (.A1(_04451_),
    .A2(_04566_),
    .B1(_04581_),
    .Y(_04586_));
 sky130_fd_sc_hd__o32a_1 _10456_ (.A1(_04453_),
    .A2(_04455_),
    .A3(_04457_),
    .B1(_04334_),
    .B2(_04462_),
    .X(_04587_));
 sky130_fd_sc_hd__o32ai_4 _10457_ (.A1(_04453_),
    .A2(_04455_),
    .A3(_04457_),
    .B1(_04334_),
    .B2(_04462_),
    .Y(_04588_));
 sky130_fd_sc_hd__o22ai_1 _10458_ (.A1(_04453_),
    .A2(_04461_),
    .B1(_04334_),
    .B2(_04462_),
    .Y(_04589_));
 sky130_fd_sc_hd__and3_1 _10459_ (.A(_04466_),
    .B(_04472_),
    .C(_04586_),
    .X(_04591_));
 sky130_fd_sc_hd__o211ai_4 _10460_ (.A1(_04334_),
    .A2(_04462_),
    .B1(_04466_),
    .C1(_04586_),
    .Y(_04592_));
 sky130_fd_sc_hd__nand2_2 _10461_ (.A(_04588_),
    .B(_04585_),
    .Y(_04593_));
 sky130_fd_sc_hd__a31oi_1 _10462_ (.A1(_04454_),
    .A2(_04458_),
    .A3(_04456_),
    .B1(_04333_),
    .Y(_04594_));
 sky130_fd_sc_hd__a31o_1 _10463_ (.A1(_04454_),
    .A2(_04458_),
    .A3(_04456_),
    .B1(_04333_),
    .X(_04595_));
 sky130_fd_sc_hd__o211ai_1 _10464_ (.A1(_04580_),
    .A2(_04582_),
    .B1(_04595_),
    .C1(_04463_),
    .Y(_04596_));
 sky130_fd_sc_hd__o21ai_1 _10465_ (.A1(_04462_),
    .A2(_04594_),
    .B1(_04585_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _10466_ (.A(_04589_),
    .B(_04585_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_1 _10467_ (.A(_04596_),
    .B(_04597_),
    .Y(_04599_));
 sky130_fd_sc_hd__a22oi_4 _10468_ (.A1(_04469_),
    .A2(_04338_),
    .B1(_04593_),
    .B2(_04592_),
    .Y(_04600_));
 sky130_fd_sc_hd__o2bb2ai_1 _10469_ (.A1_N(_04592_),
    .A2_N(_04598_),
    .B1(_04337_),
    .B2(_04474_),
    .Y(_04602_));
 sky130_fd_sc_hd__o211a_2 _10470_ (.A1(_04585_),
    .A2(_04589_),
    .B1(_04338_),
    .C1(_04469_),
    .X(_04603_));
 sky130_fd_sc_hd__a31o_1 _10471_ (.A1(_04466_),
    .A2(_04472_),
    .A3(_04586_),
    .B1(_04478_),
    .X(_04604_));
 sky130_fd_sc_hd__o21ai_1 _10472_ (.A1(_04478_),
    .A2(_04591_),
    .B1(_04602_),
    .Y(_04605_));
 sky130_fd_sc_hd__o21ai_2 _10473_ (.A1(_04338_),
    .A2(_04473_),
    .B1(_04351_),
    .Y(_04606_));
 sky130_fd_sc_hd__o22ai_4 _10474_ (.A1(_04475_),
    .A2(_04352_),
    .B1(_04603_),
    .B2(_04600_),
    .Y(_04607_));
 sky130_fd_sc_hd__and4_1 _10475_ (.A(_04476_),
    .B(_04592_),
    .C(_04593_),
    .D(_04351_),
    .X(_04608_));
 sky130_fd_sc_hd__nand4_4 _10476_ (.A(_04476_),
    .B(_04592_),
    .C(_04593_),
    .D(_04351_),
    .Y(_04609_));
 sky130_fd_sc_hd__o21ai_1 _10477_ (.A1(_04600_),
    .A2(_04606_),
    .B1(_04607_),
    .Y(_04610_));
 sky130_fd_sc_hd__o2111ai_4 _10478_ (.A1(_04340_),
    .A2(_04468_),
    .B1(_04341_),
    .C1(_04235_),
    .D1(_04476_),
    .Y(_04611_));
 sky130_fd_sc_hd__a22oi_4 _10479_ (.A1(_04348_),
    .A2(_04479_),
    .B1(_04607_),
    .B2(_04609_),
    .Y(_04613_));
 sky130_fd_sc_hd__o2bb2ai_1 _10480_ (.A1_N(_04607_),
    .A2_N(_04609_),
    .B1(_04349_),
    .B2(_04480_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand4_2 _10481_ (.A(_04607_),
    .B(_04473_),
    .C(_04341_),
    .D(_04235_),
    .Y(_04615_));
 sky130_fd_sc_hd__a21oi_4 _10482_ (.A1(_04605_),
    .A2(_04606_),
    .B1(_04611_),
    .Y(_04616_));
 sky130_fd_sc_hd__o22ai_4 _10483_ (.A1(_04485_),
    .A2(_04356_),
    .B1(_04616_),
    .B2(_04613_),
    .Y(_04617_));
 sky130_fd_sc_hd__nand3_2 _10484_ (.A(_04614_),
    .B(_04615_),
    .C(_04488_),
    .Y(_04618_));
 sky130_fd_sc_hd__a21oi_1 _10485_ (.A1(_04610_),
    .A2(_04611_),
    .B1(_04489_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_2 _10486_ (.A(_04614_),
    .B(_04488_),
    .Y(_04620_));
 sky130_fd_sc_hd__o21ai_2 _10487_ (.A1(_04489_),
    .A2(_04613_),
    .B1(_04617_),
    .Y(_04621_));
 sky130_fd_sc_hd__a22oi_4 _10488_ (.A1(_04360_),
    .A2(_04490_),
    .B1(_04617_),
    .B2(_04620_),
    .Y(_04622_));
 sky130_fd_sc_hd__o2bb2ai_4 _10489_ (.A1_N(_04617_),
    .A2_N(_04618_),
    .B1(_04362_),
    .B2(_04486_),
    .Y(_04624_));
 sky130_fd_sc_hd__o311a_2 _10490_ (.A1(_04356_),
    .A2(_04485_),
    .A3(_04613_),
    .B1(_04495_),
    .C1(_04617_),
    .X(_04625_));
 sky130_fd_sc_hd__o2111ai_4 _10491_ (.A1(_04489_),
    .A2(_04613_),
    .B1(_04490_),
    .C1(_04360_),
    .D1(_04617_),
    .Y(_04626_));
 sky130_fd_sc_hd__and4_1 _10492_ (.A(_04355_),
    .B(_04617_),
    .C(_04358_),
    .D(_04487_),
    .X(_04627_));
 sky130_fd_sc_hd__and4_1 _10493_ (.A(_04494_),
    .B(_04496_),
    .C(_04244_),
    .D(_04363_),
    .X(_04628_));
 sky130_fd_sc_hd__nand2_1 _10494_ (.A(_04498_),
    .B(_04500_),
    .Y(_04629_));
 sky130_fd_sc_hd__a22oi_4 _10495_ (.A1(_04498_),
    .A2(_04500_),
    .B1(_04624_),
    .B2(_04626_),
    .Y(_04630_));
 sky130_fd_sc_hd__o22ai_4 _10496_ (.A1(_04378_),
    .A2(_04499_),
    .B1(_04622_),
    .B2(_04625_),
    .Y(_04631_));
 sky130_fd_sc_hd__nor4_2 _10497_ (.A(_04378_),
    .B(_04493_),
    .C(_04497_),
    .D(_04621_),
    .Y(_04632_));
 sky130_fd_sc_hd__or4bb_1 _10498_ (.A(_04378_),
    .B(_04621_),
    .C_N(_04496_),
    .D_N(_04494_),
    .X(_04633_));
 sky130_fd_sc_hd__nand2_2 _10499_ (.A(_04624_),
    .B(_04628_),
    .Y(_04635_));
 sky130_fd_sc_hd__nand2_1 _10500_ (.A(_04631_),
    .B(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__o311a_1 _10501_ (.A1(_04378_),
    .A2(_04499_),
    .A3(_04622_),
    .B1(_04509_),
    .C1(_04631_),
    .X(_04637_));
 sky130_fd_sc_hd__nand3_1 _10502_ (.A(_04631_),
    .B(_04635_),
    .C(_04509_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand4_1 _10503_ (.A(_04365_),
    .B(_04513_),
    .C(_04631_),
    .D(_04635_),
    .Y(_04639_));
 sky130_fd_sc_hd__and4_1 _10504_ (.A(_04365_),
    .B(_04508_),
    .C(_04631_),
    .D(_04635_),
    .X(_04640_));
 sky130_fd_sc_hd__nand4_1 _10505_ (.A(_04365_),
    .B(_04508_),
    .C(_04631_),
    .D(_04635_),
    .Y(_04641_));
 sky130_fd_sc_hd__o22ai_1 _10506_ (.A1(_04507_),
    .A2(_04504_),
    .B1(_04632_),
    .B2(_04630_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand2_1 _10507_ (.A(_04631_),
    .B(_04512_),
    .Y(_04643_));
 sky130_fd_sc_hd__a22oi_2 _10508_ (.A1(_04365_),
    .A2(_04513_),
    .B1(_04642_),
    .B2(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__nor2_1 _10509_ (.A(_04640_),
    .B(_04644_),
    .Y(_04646_));
 sky130_fd_sc_hd__nor3b_1 _10510_ (.A(_04251_),
    .B(_04364_),
    .C_N(_04508_),
    .Y(_04647_));
 sky130_fd_sc_hd__and4bb_1 _10511_ (.A_N(_04249_),
    .B_N(_04364_),
    .C(_04513_),
    .D(_04646_),
    .X(_04648_));
 sky130_fd_sc_hd__or4bb_1 _10512_ (.A(_04249_),
    .B(_04364_),
    .C_N(_04513_),
    .D_N(_04646_),
    .X(_04649_));
 sky130_fd_sc_hd__o211a_1 _10513_ (.A1(_04646_),
    .A2(_04647_),
    .B1(_04649_),
    .C1(_03948_),
    .X(_04650_));
 sky130_fd_sc_hd__a21oi_1 _10514_ (.A1(net65),
    .A2(_04532_),
    .B1(_03949_),
    .Y(_04651_));
 sky130_fd_sc_hd__o22ai_1 _10515_ (.A1(_04529_),
    .A2(_02989_),
    .B1(_04651_),
    .B2(_04650_),
    .Y(net85));
 sky130_fd_sc_hd__a21oi_1 _10516_ (.A1(net52),
    .A2(net20),
    .B1(_01857_),
    .Y(_04652_));
 sky130_fd_sc_hd__a22o_1 _10517_ (.A1(net52),
    .A2(net20),
    .B1(_01835_),
    .B2(_01846_),
    .X(_04653_));
 sky130_fd_sc_hd__and3_1 _10518_ (.A(net52),
    .B(net20),
    .C(_01857_),
    .X(_04654_));
 sky130_fd_sc_hd__or2_1 _10519_ (.A(_04652_),
    .B(_04654_),
    .X(_04656_));
 sky130_fd_sc_hd__or4_1 _10520_ (.A(_04521_),
    .B(_04523_),
    .C(_04652_),
    .D(_04654_),
    .X(_04657_));
 sky130_fd_sc_hd__o21ai_1 _10521_ (.A1(_04521_),
    .A2(_04523_),
    .B1(_04656_),
    .Y(_04658_));
 sky130_fd_sc_hd__nand2_1 _10522_ (.A(_04657_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__o21bai_1 _10523_ (.A1(_04528_),
    .A2(_04659_),
    .B1_N(_02996_),
    .Y(_04660_));
 sky130_fd_sc_hd__a21oi_1 _10524_ (.A1(_04528_),
    .A2(_04659_),
    .B1(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__or3_1 _10525_ (.A(net21),
    .B(_02033_),
    .C(_02055_),
    .X(_04662_));
 sky130_fd_sc_hd__o31a_1 _10526_ (.A1(net53),
    .A2(_01989_),
    .A3(_02011_),
    .B1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__o21ai_2 _10527_ (.A1(net53),
    .A2(_02088_),
    .B1(_04662_),
    .Y(_04664_));
 sky130_fd_sc_hd__o21a_1 _10528_ (.A1(_04388_),
    .A2(_04389_),
    .B1(_04533_),
    .X(_04665_));
 sky130_fd_sc_hd__a31o_1 _10529_ (.A1(net99),
    .A2(_04395_),
    .A3(_04665_),
    .B1(_04664_),
    .X(_04667_));
 sky130_fd_sc_hd__nand4_4 _10530_ (.A(net99),
    .B(_04395_),
    .C(_04664_),
    .D(_04665_),
    .Y(_04668_));
 sky130_fd_sc_hd__o2bb2ai_2 _10531_ (.A1_N(_04667_),
    .A2_N(_04668_),
    .B1(_04532_),
    .B2(_04403_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand4_4 _10532_ (.A(_04402_),
    .B(_04533_),
    .C(_04667_),
    .D(_04668_),
    .Y(_04670_));
 sky130_fd_sc_hd__nand4_4 _10533_ (.A(_04383_),
    .B(_04407_),
    .C(_04540_),
    .D(_04669_),
    .Y(_04671_));
 sky130_fd_sc_hd__o2bb2ai_4 _10534_ (.A1_N(_04669_),
    .A2_N(_04670_),
    .B1(_04539_),
    .B2(_04410_),
    .Y(_04672_));
 sky130_fd_sc_hd__nand2_1 _10535_ (.A(_04671_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__a22oi_4 _10536_ (.A1(_04671_),
    .A2(_04672_),
    .B1(_04417_),
    .B2(_04540_),
    .Y(_04674_));
 sky130_fd_sc_hd__o2bb2ai_2 _10537_ (.A1_N(_04671_),
    .A2_N(_04672_),
    .B1(_04418_),
    .B2(_04539_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand4_4 _10538_ (.A(_04417_),
    .B(_04540_),
    .C(_04671_),
    .D(_04672_),
    .Y(_04676_));
 sky130_fd_sc_hd__nand2_1 _10539_ (.A(_04675_),
    .B(_04676_),
    .Y(_04678_));
 sky130_fd_sc_hd__o31a_1 _10540_ (.A1(_04420_),
    .A2(_04424_),
    .A3(_04545_),
    .B1(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__o2bb2ai_2 _10541_ (.A1_N(_04675_),
    .A2_N(_04676_),
    .B1(_04545_),
    .B2(_04547_),
    .Y(_04680_));
 sky130_fd_sc_hd__nand4_2 _10542_ (.A(_04419_),
    .B(_04423_),
    .C(_04675_),
    .D(_04544_),
    .Y(_04681_));
 sky130_fd_sc_hd__o31a_1 _10543_ (.A1(_04545_),
    .A2(_04547_),
    .A3(_04674_),
    .B1(_04680_),
    .X(_04682_));
 sky130_fd_sc_hd__a22oi_4 _10544_ (.A1(_04549_),
    .A2(_04551_),
    .B1(_04680_),
    .B2(_04681_),
    .Y(_04683_));
 sky130_fd_sc_hd__nand3_1 _10545_ (.A(_04554_),
    .B(_04675_),
    .C(_04676_),
    .Y(_04684_));
 sky130_fd_sc_hd__a21oi_2 _10546_ (.A1(_04550_),
    .A2(_04678_),
    .B1(_04555_),
    .Y(_04685_));
 sky130_fd_sc_hd__and4_1 _10547_ (.A(_04551_),
    .B(_04675_),
    .C(_04676_),
    .D(_04549_),
    .X(_04686_));
 sky130_fd_sc_hd__o2111ai_4 _10548_ (.A1(_04548_),
    .A2(_04552_),
    .B1(_04307_),
    .C1(_04553_),
    .D1(_04425_),
    .Y(_04687_));
 sky130_fd_sc_hd__o22ai_4 _10549_ (.A1(_04433_),
    .A2(_04558_),
    .B1(_04683_),
    .B2(_04685_),
    .Y(_04689_));
 sky130_fd_sc_hd__or4bb_1 _10550_ (.A(_04554_),
    .B(_04433_),
    .C_N(_04553_),
    .D_N(_04682_),
    .X(_04690_));
 sky130_fd_sc_hd__nand4_2 _10551_ (.A(_04434_),
    .B(_04553_),
    .C(_04680_),
    .D(_04681_),
    .Y(_04691_));
 sky130_fd_sc_hd__and3_1 _10552_ (.A(_04553_),
    .B(_04309_),
    .C(_04432_),
    .X(_04692_));
 sky130_fd_sc_hd__a22oi_4 _10553_ (.A1(_04556_),
    .A2(_04562_),
    .B1(_04689_),
    .B2(_04691_),
    .Y(_04693_));
 sky130_fd_sc_hd__a22o_1 _10554_ (.A1(_04556_),
    .A2(_04562_),
    .B1(_04689_),
    .B2(_04691_),
    .X(_04694_));
 sky130_fd_sc_hd__o211a_1 _10555_ (.A1(_04683_),
    .A2(_04687_),
    .B1(_04692_),
    .C1(_04689_),
    .X(_04695_));
 sky130_fd_sc_hd__o211ai_1 _10556_ (.A1(_04683_),
    .A2(_04687_),
    .B1(_04692_),
    .C1(_04689_),
    .Y(_04696_));
 sky130_fd_sc_hd__a21oi_2 _10557_ (.A1(_04689_),
    .A2(_04692_),
    .B1(_04693_),
    .Y(_04697_));
 sky130_fd_sc_hd__inv_2 _10558_ (.A(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__o211ai_4 _10559_ (.A1(_04693_),
    .A2(_04695_),
    .B1(_04571_),
    .C1(_04583_),
    .Y(_04700_));
 sky130_fd_sc_hd__o221ai_4 _10560_ (.A1(_04444_),
    .A2(_04565_),
    .B1(_04570_),
    .B2(_04450_),
    .C1(_04694_),
    .Y(_04701_));
 sky130_fd_sc_hd__o2bb2ai_4 _10561_ (.A1_N(_04700_),
    .A2_N(_04701_),
    .B1(_04456_),
    .B2(_04573_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand3_1 _10562_ (.A(_04700_),
    .B(_04701_),
    .C(_04576_),
    .Y(_04703_));
 sky130_fd_sc_hd__nand2_2 _10563_ (.A(_04700_),
    .B(_04576_),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2_1 _10564_ (.A(_04702_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__nand3_2 _10565_ (.A(_04585_),
    .B(_04702_),
    .C(_04704_),
    .Y(_04706_));
 sky130_fd_sc_hd__inv_2 _10566_ (.A(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__nand4_1 _10567_ (.A(_04588_),
    .B(_04702_),
    .C(_04704_),
    .D(_04585_),
    .Y(_04708_));
 sky130_fd_sc_hd__a22o_1 _10568_ (.A1(_04702_),
    .A2(_04704_),
    .B1(_04588_),
    .B2(_04585_),
    .X(_04709_));
 sky130_fd_sc_hd__a32o_1 _10569_ (.A1(_04454_),
    .A2(_04460_),
    .A3(_04581_),
    .B1(_04702_),
    .B2(_04704_),
    .X(_04711_));
 sky130_fd_sc_hd__nand4_1 _10570_ (.A(_04465_),
    .B(_04585_),
    .C(_04702_),
    .D(_04704_),
    .Y(_04712_));
 sky130_fd_sc_hd__a22oi_2 _10571_ (.A1(_04471_),
    .A2(_04585_),
    .B1(_04711_),
    .B2(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__a2bb2oi_2 _10572_ (.A1_N(_04587_),
    .A2_N(_04706_),
    .B1(_04705_),
    .B2(_04593_),
    .Y(_04714_));
 sky130_fd_sc_hd__o2bb2ai_1 _10573_ (.A1_N(_04593_),
    .A2_N(_04705_),
    .B1(_04706_),
    .B2(_04587_),
    .Y(_04715_));
 sky130_fd_sc_hd__o21ai_1 _10574_ (.A1(_04478_),
    .A2(_04591_),
    .B1(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand4_2 _10575_ (.A(_04709_),
    .B(_04599_),
    .C(_04477_),
    .D(_04708_),
    .Y(_04717_));
 sky130_fd_sc_hd__nor2_1 _10576_ (.A(_04604_),
    .B(_04713_),
    .Y(_04718_));
 sky130_fd_sc_hd__o21ai_4 _10577_ (.A1(_04603_),
    .A2(_04714_),
    .B1(_04717_),
    .Y(_04719_));
 sky130_fd_sc_hd__o21ai_2 _10578_ (.A1(_04600_),
    .A2(_04606_),
    .B1(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__a21oi_2 _10579_ (.A1(_04604_),
    .A2(_04715_),
    .B1(_04609_),
    .Y(_04722_));
 sky130_fd_sc_hd__o21ai_4 _10580_ (.A1(_04603_),
    .A2(_04714_),
    .B1(_04608_),
    .Y(_04723_));
 sky130_fd_sc_hd__a21oi_4 _10581_ (.A1(_04609_),
    .A2(_04719_),
    .B1(_04722_),
    .Y(_04724_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_04720_),
    .B(_04723_),
    .Y(_04725_));
 sky130_fd_sc_hd__o2111ai_4 _10583_ (.A1(_04600_),
    .A2(_04352_),
    .B1(_04348_),
    .C1(_04476_),
    .D1(_04607_),
    .Y(_04726_));
 sky130_fd_sc_hd__a21oi_4 _10584_ (.A1(_04720_),
    .A2(_04723_),
    .B1(_04616_),
    .Y(_04727_));
 sky130_fd_sc_hd__a21o_1 _10585_ (.A1(_04720_),
    .A2(_04723_),
    .B1(_04616_),
    .X(_04728_));
 sky130_fd_sc_hd__nand3_1 _10586_ (.A(_04616_),
    .B(_04720_),
    .C(_04723_),
    .Y(_04729_));
 sky130_fd_sc_hd__a21oi_2 _10587_ (.A1(_04609_),
    .A2(_04719_),
    .B1(_04726_),
    .Y(_04730_));
 sky130_fd_sc_hd__a21o_1 _10588_ (.A1(_04609_),
    .A2(_04719_),
    .B1(_04726_),
    .X(_04731_));
 sky130_fd_sc_hd__a21o_2 _10589_ (.A1(_04725_),
    .A2(_04726_),
    .B1(_04730_),
    .X(_04733_));
 sky130_fd_sc_hd__o21ai_2 _10590_ (.A1(_04615_),
    .A2(_04725_),
    .B1(_04618_),
    .Y(_04734_));
 sky130_fd_sc_hd__o22ai_4 _10591_ (.A1(_04613_),
    .A2(_04489_),
    .B1(_04730_),
    .B2(_04727_),
    .Y(_04735_));
 sky130_fd_sc_hd__o21ai_4 _10592_ (.A1(_04616_),
    .A2(_04724_),
    .B1(_04619_),
    .Y(_04736_));
 sky130_fd_sc_hd__o21ai_1 _10593_ (.A1(_04620_),
    .A2(_04727_),
    .B1(_04735_),
    .Y(_04737_));
 sky130_fd_sc_hd__a21oi_2 _10594_ (.A1(_04735_),
    .A2(_04736_),
    .B1(_04625_),
    .Y(_04738_));
 sky130_fd_sc_hd__o2bb2ai_4 _10595_ (.A1_N(_04735_),
    .A2_N(_04736_),
    .B1(_04496_),
    .B2(_04621_),
    .Y(_04739_));
 sky130_fd_sc_hd__and3_1 _10596_ (.A(_04625_),
    .B(_04728_),
    .C(_04731_),
    .X(_04740_));
 sky130_fd_sc_hd__and3_1 _10597_ (.A(_04735_),
    .B(_04497_),
    .C(_04617_),
    .X(_04741_));
 sky130_fd_sc_hd__nand2_1 _10598_ (.A(_04627_),
    .B(_04735_),
    .Y(_04742_));
 sky130_fd_sc_hd__o21ai_4 _10599_ (.A1(_04626_),
    .A2(_04733_),
    .B1(_04739_),
    .Y(_04744_));
 sky130_fd_sc_hd__o31a_1 _10600_ (.A1(_04626_),
    .A2(_04727_),
    .A3(_04730_),
    .B1(_04739_),
    .X(_04745_));
 sky130_fd_sc_hd__a221oi_1 _10601_ (.A1(_04631_),
    .A2(_04509_),
    .B1(_04742_),
    .B2(_04739_),
    .C1(_04632_),
    .Y(_04746_));
 sky130_fd_sc_hd__o221ai_4 _10602_ (.A1(_04510_),
    .A2(_04630_),
    .B1(_04738_),
    .B2(_04741_),
    .C1(_04633_),
    .Y(_04747_));
 sky130_fd_sc_hd__o211ai_2 _10603_ (.A1(_04626_),
    .A2(_04733_),
    .B1(_04632_),
    .C1(_04739_),
    .Y(_04748_));
 sky130_fd_sc_hd__o21ai_1 _10604_ (.A1(_04744_),
    .A2(_04638_),
    .B1(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__a22oi_1 _10605_ (.A1(_04631_),
    .A2(_04512_),
    .B1(_04742_),
    .B2(_04739_),
    .Y(_04750_));
 sky130_fd_sc_hd__nor3b_1 _10606_ (.A(_04744_),
    .B(_04636_),
    .C_N(_04512_),
    .Y(_04751_));
 sky130_fd_sc_hd__o2111a_1 _10607_ (.A1(_04626_),
    .A2(_04733_),
    .B1(_04512_),
    .C1(_04739_),
    .D1(_04631_),
    .X(_04752_));
 sky130_fd_sc_hd__o2111ai_2 _10608_ (.A1(_04626_),
    .A2(_04733_),
    .B1(_04512_),
    .C1(_04739_),
    .D1(_04631_),
    .Y(_04753_));
 sky130_fd_sc_hd__o32ai_2 _10609_ (.A1(_04378_),
    .A2(_04499_),
    .A3(_04622_),
    .B1(_04750_),
    .B2(_04752_),
    .Y(_04755_));
 sky130_fd_sc_hd__o211a_1 _10610_ (.A1(_04744_),
    .A2(_04638_),
    .B1(_04748_),
    .C1(_04747_),
    .X(_04756_));
 sky130_fd_sc_hd__o211ai_2 _10611_ (.A1(_04744_),
    .A2(_04638_),
    .B1(_04748_),
    .C1(_04747_),
    .Y(_04757_));
 sky130_fd_sc_hd__nor4_1 _10612_ (.A(_04246_),
    .B(_04364_),
    .C(_04515_),
    .D(_04636_),
    .Y(_04758_));
 sky130_fd_sc_hd__o41a_1 _10613_ (.A1(_04246_),
    .A2(_04364_),
    .A3(_04515_),
    .A4(_04636_),
    .B1(_04757_),
    .X(_04759_));
 sky130_fd_sc_hd__a21oi_1 _10614_ (.A1(_04640_),
    .A2(_04755_),
    .B1(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__and4bb_1 _10615_ (.A_N(_04757_),
    .B_N(_04644_),
    .C(_04641_),
    .D(_04647_),
    .X(_04761_));
 sky130_fd_sc_hd__or4bb_2 _10616_ (.A(_04757_),
    .B(_04644_),
    .C_N(_04641_),
    .D_N(_04647_),
    .X(_04762_));
 sky130_fd_sc_hd__o211a_1 _10617_ (.A1(_04648_),
    .A2(_04760_),
    .B1(_04762_),
    .C1(_03948_),
    .X(_04763_));
 sky130_fd_sc_hd__o21ai_1 _10618_ (.A1(_04663_),
    .A2(_03948_),
    .B1(net65),
    .Y(_04764_));
 sky130_fd_sc_hd__o22ai_1 _10619_ (.A1(_02989_),
    .A2(_04661_),
    .B1(_04764_),
    .B2(_04763_),
    .Y(net86));
 sky130_fd_sc_hd__or4_1 _10620_ (.A(_04521_),
    .B(_04522_),
    .C(_04656_),
    .D(_04519_),
    .X(_04766_));
 sky130_fd_sc_hd__o31ai_2 _10621_ (.A1(_04521_),
    .A2(_04523_),
    .A3(_04654_),
    .B1(_04653_),
    .Y(_04767_));
 sky130_fd_sc_hd__xor2_1 _10622_ (.A(_01571_),
    .B(_01846_),
    .X(_04768_));
 sky130_fd_sc_hd__xnor2_1 _10623_ (.A(_04767_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__o21ai_1 _10624_ (.A1(_04086_),
    .A2(_04766_),
    .B1(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__or4_1 _10625_ (.A(_02132_),
    .B(_04766_),
    .C(_04769_),
    .D(_02976_),
    .X(_04771_));
 sky130_fd_sc_hd__a21oi_1 _10626_ (.A1(_04770_),
    .A2(_04771_),
    .B1(_02996_),
    .Y(_04772_));
 sky130_fd_sc_hd__or3_2 _10627_ (.A(_01549_),
    .B(_01945_),
    .C(_01956_),
    .X(_04773_));
 sky130_fd_sc_hd__o31a_1 _10628_ (.A1(_01549_),
    .A2(_01945_),
    .A3(_01956_),
    .B1(_01538_),
    .X(_04774_));
 sky130_fd_sc_hd__o2111ai_4 _10629_ (.A1(net54),
    .A2(net22),
    .B1(_04668_),
    .C1(_04670_),
    .D1(_04773_),
    .Y(_04776_));
 sky130_fd_sc_hd__a21o_1 _10630_ (.A1(_01538_),
    .A2(_04773_),
    .B1(_04670_),
    .X(_04777_));
 sky130_fd_sc_hd__or4_2 _10631_ (.A(_04532_),
    .B(_04663_),
    .C(_04774_),
    .D(_04399_),
    .X(_04778_));
 sky130_fd_sc_hd__o211ai_1 _10632_ (.A1(_04774_),
    .A2(_04670_),
    .B1(_04778_),
    .C1(_04776_),
    .Y(_04779_));
 sky130_fd_sc_hd__nand4b_2 _10633_ (.A_N(_04671_),
    .B(_04776_),
    .C(_04777_),
    .D(_04778_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _10634_ (.A(_04671_),
    .B(_04779_),
    .Y(_04781_));
 sky130_fd_sc_hd__a31oi_1 _10635_ (.A1(_04776_),
    .A2(_04777_),
    .A3(_04778_),
    .B1(_04671_),
    .Y(_04782_));
 sky130_fd_sc_hd__and4_1 _10636_ (.A(_04671_),
    .B(_04776_),
    .C(_04777_),
    .D(_04778_),
    .X(_04783_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(_04780_),
    .B(_04781_),
    .Y(_04784_));
 sky130_fd_sc_hd__o32ai_2 _10638_ (.A1(_04418_),
    .A2(_04539_),
    .A3(_04673_),
    .B1(_04674_),
    .B2(_04550_),
    .Y(_04785_));
 sky130_fd_sc_hd__o211ai_2 _10639_ (.A1(_04550_),
    .A2(_04674_),
    .B1(_04676_),
    .C1(_04784_),
    .Y(_04787_));
 sky130_fd_sc_hd__o21ai_2 _10640_ (.A1(_04782_),
    .A2(_04783_),
    .B1(_04785_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand2_1 _10641_ (.A(_04787_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__a21oi_1 _10642_ (.A1(_04787_),
    .A2(_04788_),
    .B1(_04685_),
    .Y(_04790_));
 sky130_fd_sc_hd__o2bb2ai_1 _10643_ (.A1_N(_04787_),
    .A2_N(_04788_),
    .B1(_04555_),
    .B2(_04679_),
    .Y(_04791_));
 sky130_fd_sc_hd__o21a_1 _10644_ (.A1(_04684_),
    .A2(_04789_),
    .B1(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__o2111ai_2 _10645_ (.A1(_04682_),
    .A2(_04554_),
    .B1(_04434_),
    .C1(_04556_),
    .D1(_04790_),
    .Y(_04793_));
 sky130_fd_sc_hd__nand3_1 _10646_ (.A(_04686_),
    .B(_04787_),
    .C(_04788_),
    .Y(_04794_));
 sky130_fd_sc_hd__o211ai_1 _10647_ (.A1(_04687_),
    .A2(_04683_),
    .B1(_04794_),
    .C1(_04791_),
    .Y(_04795_));
 sky130_fd_sc_hd__nand2_1 _10648_ (.A(_04793_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__nand3_1 _10649_ (.A(_04696_),
    .B(_04793_),
    .C(_04795_),
    .Y(_04798_));
 sky130_fd_sc_hd__nand4_2 _10650_ (.A(_04792_),
    .B(_04690_),
    .C(_04689_),
    .D(_04692_),
    .Y(_04799_));
 sky130_fd_sc_hd__o2bb2ai_2 _10651_ (.A1_N(_04798_),
    .A2_N(_04799_),
    .B1(_04572_),
    .B2(_04693_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand4_2 _10652_ (.A(_04798_),
    .B(_04565_),
    .C(_04444_),
    .D(_04694_),
    .Y(_04801_));
 sky130_fd_sc_hd__and3_1 _10653_ (.A(_04582_),
    .B(_04694_),
    .C(_04696_),
    .X(_04802_));
 sky130_fd_sc_hd__o2bb2ai_2 _10654_ (.A1_N(_04800_),
    .A2_N(_04801_),
    .B1(_04583_),
    .B2(_04698_),
    .Y(_04803_));
 sky130_fd_sc_hd__nand4_2 _10655_ (.A(_04800_),
    .B(_04801_),
    .C(_04582_),
    .D(_04697_),
    .Y(_04804_));
 sky130_fd_sc_hd__nand2_1 _10656_ (.A(_04803_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__nand2_1 _10657_ (.A(_04704_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__nand4_2 _10658_ (.A(_04803_),
    .B(_04576_),
    .C(_04700_),
    .D(_04804_),
    .Y(_04807_));
 sky130_fd_sc_hd__a2bb2oi_1 _10659_ (.A1_N(_04706_),
    .A2_N(_04587_),
    .B1(_04807_),
    .B2(_04806_),
    .Y(_04809_));
 sky130_fd_sc_hd__a22o_1 _10660_ (.A1(_04707_),
    .A2(_04588_),
    .B1(_04807_),
    .B2(_04806_),
    .X(_04810_));
 sky130_fd_sc_hd__o2111ai_1 _10661_ (.A1(_04464_),
    .A2(_04471_),
    .B1(_04807_),
    .C1(_04707_),
    .D1(_04806_),
    .Y(_04811_));
 sky130_fd_sc_hd__a41oi_2 _10662_ (.A1(_04588_),
    .A2(_04707_),
    .A3(_04806_),
    .A4(_04807_),
    .B1(_04809_),
    .Y(_04812_));
 sky130_fd_sc_hd__nand2_1 _10663_ (.A(_04810_),
    .B(_04811_),
    .Y(_04813_));
 sky130_fd_sc_hd__a2bb2oi_1 _10664_ (.A1_N(_04604_),
    .A2_N(_04713_),
    .B1(_04608_),
    .B2(_04716_),
    .Y(_04814_));
 sky130_fd_sc_hd__o211a_1 _10665_ (.A1(_04604_),
    .A2(_04713_),
    .B1(_04723_),
    .C1(_04813_),
    .X(_04815_));
 sky130_fd_sc_hd__nand2_1 _10666_ (.A(_04814_),
    .B(_04813_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _10667_ (.A(_04812_),
    .B(_04814_),
    .Y(_04817_));
 sky130_fd_sc_hd__o21ai_1 _10668_ (.A1(_04718_),
    .A2(_04722_),
    .B1(_04813_),
    .Y(_04818_));
 sky130_fd_sc_hd__o211a_1 _10669_ (.A1(_04718_),
    .A2(_04722_),
    .B1(_04810_),
    .C1(_04811_),
    .X(_04820_));
 sky130_fd_sc_hd__o21ai_1 _10670_ (.A1(_04718_),
    .A2(_04722_),
    .B1(_04812_),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _10671_ (.A(_04817_),
    .B(_04818_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand2_2 _10672_ (.A(_04816_),
    .B(_04821_),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_1 _10673_ (.A(_04618_),
    .B(_04729_),
    .Y(_04824_));
 sky130_fd_sc_hd__a21o_1 _10674_ (.A1(_04618_),
    .A2(_04729_),
    .B1(_04727_),
    .X(_04825_));
 sky130_fd_sc_hd__o211a_1 _10675_ (.A1(_04620_),
    .A2(_04727_),
    .B1(_04731_),
    .C1(_04823_),
    .X(_04826_));
 sky130_fd_sc_hd__o211ai_4 _10676_ (.A1(_04620_),
    .A2(_04727_),
    .B1(_04731_),
    .C1(_04823_),
    .Y(_04827_));
 sky130_fd_sc_hd__o211ai_4 _10677_ (.A1(_04616_),
    .A2(_04724_),
    .B1(_04822_),
    .C1(_04734_),
    .Y(_04828_));
 sky130_fd_sc_hd__o211ai_1 _10678_ (.A1(_04616_),
    .A2(_04724_),
    .B1(_04822_),
    .C1(_04824_),
    .Y(_04829_));
 sky130_fd_sc_hd__a21oi_2 _10679_ (.A1(_04731_),
    .A2(_04736_),
    .B1(_04823_),
    .Y(_04831_));
 sky130_fd_sc_hd__nor2_1 _10680_ (.A(_04826_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__a31o_1 _10681_ (.A1(_04728_),
    .A2(_04734_),
    .A3(_04816_),
    .B1(_04826_),
    .X(_04833_));
 sky130_fd_sc_hd__o22ai_4 _10682_ (.A1(_04626_),
    .A2(_04733_),
    .B1(_04826_),
    .B2(_04831_),
    .Y(_04834_));
 sky130_fd_sc_hd__nand2_1 _10683_ (.A(_04740_),
    .B(_04832_),
    .Y(_04835_));
 sky130_fd_sc_hd__and4_1 _10684_ (.A(_04735_),
    .B(_04827_),
    .C(_04828_),
    .D(_04627_),
    .X(_04836_));
 sky130_fd_sc_hd__nand4_4 _10685_ (.A(_04735_),
    .B(_04827_),
    .C(_04828_),
    .D(_04627_),
    .Y(_04837_));
 sky130_fd_sc_hd__nand2_1 _10686_ (.A(_04834_),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__nor4_1 _10687_ (.A(_04622_),
    .B(_04625_),
    .C(_04629_),
    .D(_04737_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand4b_2 _10688_ (.A_N(_04629_),
    .B(_04739_),
    .C(_04624_),
    .D(_04626_),
    .Y(_04840_));
 sky130_fd_sc_hd__a21oi_1 _10689_ (.A1(_04834_),
    .A2(_04837_),
    .B1(_04839_),
    .Y(_04842_));
 sky130_fd_sc_hd__o2bb2ai_1 _10690_ (.A1_N(_04834_),
    .A2_N(_04837_),
    .B1(_04635_),
    .B2(_04744_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand4_2 _10691_ (.A(_04624_),
    .B(_04828_),
    .C(_04628_),
    .D(_04827_),
    .Y(_04844_));
 sky130_fd_sc_hd__a21oi_1 _10692_ (.A1(_04626_),
    .A2(_04737_),
    .B1(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__a21o_1 _10693_ (.A1(_04626_),
    .A2(_04737_),
    .B1(_04844_),
    .X(_04846_));
 sky130_fd_sc_hd__a21oi_1 _10694_ (.A1(_04838_),
    .A2(_04840_),
    .B1(_04845_),
    .Y(_04847_));
 sky130_fd_sc_hd__o21ai_1 _10695_ (.A1(_04833_),
    .A2(_04840_),
    .B1(_04843_),
    .Y(_04848_));
 sky130_fd_sc_hd__o21ai_1 _10696_ (.A1(_04641_),
    .A2(_04757_),
    .B1(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__nor4_1 _10697_ (.A(_04639_),
    .B(_04838_),
    .C(_04746_),
    .D(_04749_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand4_1 _10698_ (.A(_04756_),
    .B(_04758_),
    .C(_04834_),
    .D(_04837_),
    .Y(_04851_));
 sky130_fd_sc_hd__nand4_1 _10699_ (.A(_04755_),
    .B(_04834_),
    .C(_04837_),
    .D(_04640_),
    .Y(_04853_));
 sky130_fd_sc_hd__nor3b_1 _10700_ (.A(_04744_),
    .B(_04636_),
    .C_N(_04511_),
    .Y(_04854_));
 sky130_fd_sc_hd__a21oi_1 _10701_ (.A1(_04849_),
    .A2(_04853_),
    .B1(_04751_),
    .Y(_04855_));
 sky130_fd_sc_hd__a21o_1 _10702_ (.A1(_04849_),
    .A2(_04853_),
    .B1(_04751_),
    .X(_04856_));
 sky130_fd_sc_hd__nand4_1 _10703_ (.A(_04843_),
    .B(_04637_),
    .C(_04745_),
    .D(_04846_),
    .Y(_04857_));
 sky130_fd_sc_hd__o21ai_1 _10704_ (.A1(_04753_),
    .A2(_04842_),
    .B1(_04856_),
    .Y(_04858_));
 sky130_fd_sc_hd__o21ai_1 _10705_ (.A1(_04762_),
    .A2(_04855_),
    .B1(_03948_),
    .Y(_04859_));
 sky130_fd_sc_hd__a21oi_2 _10706_ (.A1(_04762_),
    .A2(_04858_),
    .B1(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__a21oi_1 _10707_ (.A1(net65),
    .A2(_04774_),
    .B1(_03949_),
    .Y(_04861_));
 sky130_fd_sc_hd__o22ai_1 _10708_ (.A1(_04772_),
    .A2(_02989_),
    .B1(_04861_),
    .B2(_04860_),
    .Y(net87));
 sky130_fd_sc_hd__o32a_1 _10709_ (.A1(_01527_),
    .A2(_01549_),
    .A3(_01846_),
    .B1(_04768_),
    .B2(_04767_),
    .X(_04863_));
 sky130_fd_sc_hd__o21ai_1 _10710_ (.A1(_01945_),
    .A2(_01956_),
    .B1(_01549_),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_1 _10711_ (.A(_04773_),
    .B(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__xor2_1 _10712_ (.A(_04863_),
    .B(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__a21oi_1 _10713_ (.A1(_04771_),
    .A2(_04866_),
    .B1(_02996_),
    .Y(_04867_));
 sky130_fd_sc_hd__o41a_1 _10714_ (.A1(_04086_),
    .A2(_04766_),
    .A3(_04769_),
    .A4(_04866_),
    .B1(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__a21o_1 _10715_ (.A1(_01516_),
    .A2(_01934_),
    .B1(net56),
    .X(_04869_));
 sky130_fd_sc_hd__o31a_1 _10716_ (.A1(net24),
    .A2(_01505_),
    .A3(_01923_),
    .B1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__xor2_1 _10717_ (.A(_04778_),
    .B(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__a31o_1 _10718_ (.A1(_04777_),
    .A2(_04780_),
    .A3(_04788_),
    .B1(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__o2111ai_2 _10719_ (.A1(_04670_),
    .A2(_04774_),
    .B1(_04780_),
    .C1(_04788_),
    .D1(_04871_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_04872_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__o21ai_1 _10721_ (.A1(_04691_),
    .A2(_04790_),
    .B1(_04794_),
    .Y(_04876_));
 sky130_fd_sc_hd__o311a_1 _10722_ (.A1(_04683_),
    .A2(_04687_),
    .A3(_04790_),
    .B1(_04872_),
    .C1(_04874_),
    .X(_04877_));
 sky130_fd_sc_hd__a22o_1 _10723_ (.A1(_04877_),
    .A2(_04794_),
    .B1(_04875_),
    .B2(_04876_),
    .X(_04878_));
 sky130_fd_sc_hd__xor2_1 _10724_ (.A(_04799_),
    .B(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__nand4_1 _10725_ (.A(_04803_),
    .B(_04333_),
    .C(_04463_),
    .D(_04804_),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _10726_ (.A(_04706_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__nand2_1 _10727_ (.A(_04881_),
    .B(_04879_),
    .Y(_04882_));
 sky130_fd_sc_hd__o21bai_1 _10728_ (.A1(_04706_),
    .A2(_04880_),
    .B1_N(_04879_),
    .Y(_04883_));
 sky130_fd_sc_hd__nand3_1 _10729_ (.A(_04803_),
    .B(_04804_),
    .C(_04464_),
    .Y(_04885_));
 sky130_fd_sc_hd__o32a_1 _10730_ (.A1(_04586_),
    .A2(_04705_),
    .A3(_04885_),
    .B1(_04805_),
    .B2(_04703_),
    .X(_04886_));
 sky130_fd_sc_hd__a31o_1 _10731_ (.A1(_04570_),
    .A2(_04697_),
    .A3(_04796_),
    .B1(_04802_),
    .X(_04887_));
 sky130_fd_sc_hd__nand2_1 _10732_ (.A(_04800_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__nand4_1 _10733_ (.A(_04882_),
    .B(_04883_),
    .C(_04886_),
    .D(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__a22o_1 _10734_ (.A1(_04886_),
    .A2(_04888_),
    .B1(_04882_),
    .B2(_04883_),
    .X(_04890_));
 sky130_fd_sc_hd__nand2_1 _10735_ (.A(_04889_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o2bb2a_1 _10736_ (.A1_N(_04889_),
    .A2_N(_04890_),
    .B1(_04813_),
    .B2(_04814_),
    .X(_04892_));
 sky130_fd_sc_hd__and4b_1 _10737_ (.A_N(_04814_),
    .B(_04889_),
    .C(_04890_),
    .D(_04812_),
    .X(_04893_));
 sky130_fd_sc_hd__o21ai_1 _10738_ (.A1(_04892_),
    .A2(_04893_),
    .B1(_04829_),
    .Y(_04894_));
 sky130_fd_sc_hd__o31a_1 _10739_ (.A1(_04892_),
    .A2(_04893_),
    .A3(_04829_),
    .B1(_04894_),
    .X(_04896_));
 sky130_fd_sc_hd__o41ai_2 _10740_ (.A1(_04815_),
    .A2(_04891_),
    .A3(_04820_),
    .A4(_04825_),
    .B1(_04894_),
    .Y(_04897_));
 sky130_fd_sc_hd__o211ai_1 _10741_ (.A1(_04833_),
    .A2(_04840_),
    .B1(_04896_),
    .C1(_04835_),
    .Y(_04898_));
 sky130_fd_sc_hd__o211ai_1 _10742_ (.A1(_04740_),
    .A2(_04839_),
    .B1(_04897_),
    .C1(_04832_),
    .Y(_04899_));
 sky130_fd_sc_hd__o21ai_1 _10743_ (.A1(_04738_),
    .A2(_04844_),
    .B1(_04837_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_1 _10744_ (.A(_04900_),
    .B(_04896_),
    .Y(_04901_));
 sky130_fd_sc_hd__o21ai_1 _10745_ (.A1(_04738_),
    .A2(_04844_),
    .B1(_04897_),
    .Y(_04902_));
 sky130_fd_sc_hd__o211ai_1 _10746_ (.A1(_04738_),
    .A2(_04844_),
    .B1(_04897_),
    .C1(_04837_),
    .Y(_04903_));
 sky130_fd_sc_hd__o2bb2ai_1 _10747_ (.A1_N(_04896_),
    .A2_N(_04900_),
    .B1(_04836_),
    .B2(_04902_),
    .Y(_04904_));
 sky130_fd_sc_hd__nand2_1 _10748_ (.A(_04857_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__nand4_1 _10749_ (.A(_04847_),
    .B(_04854_),
    .C(_04901_),
    .D(_04903_),
    .Y(_04907_));
 sky130_fd_sc_hd__nand4_1 _10750_ (.A(_04898_),
    .B(_04751_),
    .C(_04843_),
    .D(_04899_),
    .Y(_04908_));
 sky130_fd_sc_hd__o221ai_1 _10751_ (.A1(_04836_),
    .A2(_04902_),
    .B1(_04753_),
    .B2(_04842_),
    .C1(_04901_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand3_1 _10752_ (.A(_04851_),
    .B(_04905_),
    .C(_04907_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand3_1 _10753_ (.A(_04850_),
    .B(_04908_),
    .C(_04909_),
    .Y(_04911_));
 sky130_fd_sc_hd__nand2_1 _10754_ (.A(_04910_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__o21ai_1 _10755_ (.A1(_04762_),
    .A2(_04855_),
    .B1(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__nand4_1 _10756_ (.A(_04856_),
    .B(_04910_),
    .C(_04911_),
    .D(_04761_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand3_1 _10757_ (.A(_03948_),
    .B(_04913_),
    .C(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__o31a_1 _10758_ (.A1(_03573_),
    .A2(_03947_),
    .A3(_04870_),
    .B1(net65),
    .X(_04916_));
 sky130_fd_sc_hd__o2bb2ai_1 _10759_ (.A1_N(_04915_),
    .A2_N(_04916_),
    .B1(_02989_),
    .B2(_04868_),
    .Y(net89));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(net57),
    .A1(net25),
    .S(net102),
    .X(_04918_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(_05233_),
    .A1(_04918_),
    .S(net65),
    .X(net90));
 sky130_fd_sc_hd__or4_2 _10762_ (.A(_04975_),
    .B(\adder_inst.fraction1[0] ),
    .C(_05008_),
    .D(_05029_),
    .X(_04919_));
 sky130_fd_sc_hd__a22o_1 _10763_ (.A1(_04979_),
    .A2(_05003_),
    .B1(_05009_),
    .B2(_05030_),
    .X(_04920_));
 sky130_fd_sc_hd__and2_1 _10764_ (.A(_04919_),
    .B(_04920_),
    .X(_00038_));
 sky130_fd_sc_hd__or4_1 _10765_ (.A(_04975_),
    .B(_05032_),
    .C(\adder_inst.fraction1[0] ),
    .D(_04634_),
    .X(_04921_));
 sky130_fd_sc_hd__a31o_1 _10766_ (.A1(_04979_),
    .A2(_05003_),
    .A3(_05031_),
    .B1(_04645_),
    .X(_04922_));
 sky130_fd_sc_hd__and2_1 _10767_ (.A(_04921_),
    .B(_04922_),
    .X(_00039_));
 sky130_fd_sc_hd__xor2_1 _10768_ (.A(_04317_),
    .B(_04921_),
    .X(_00040_));
 sky130_fd_sc_hd__nor4_2 _10769_ (.A(_03880_),
    .B(_04317_),
    .C(_04634_),
    .D(_04919_),
    .Y(_04924_));
 sky130_fd_sc_hd__o31a_1 _10770_ (.A1(_04317_),
    .A2(_04634_),
    .A3(_04919_),
    .B1(_03880_),
    .X(_04925_));
 sky130_fd_sc_hd__nor2_1 _10771_ (.A(_04924_),
    .B(_04925_),
    .Y(_00041_));
 sky130_fd_sc_hd__xor2_1 _10772_ (.A(_05050_),
    .B(_04924_),
    .X(_00042_));
 sky130_fd_sc_hd__or4b_1 _10773_ (.A(_05049_),
    .B(_05064_),
    .C(_05065_),
    .D_N(_04924_),
    .X(_04926_));
 sky130_fd_sc_hd__a221o_1 _10774_ (.A1(_01175_),
    .A2(_02088_),
    .B1(_05050_),
    .B2(_04924_),
    .C1(_05067_),
    .X(_04927_));
 sky130_fd_sc_hd__and2_1 _10775_ (.A(_04926_),
    .B(_04927_),
    .X(_00043_));
 sky130_fd_sc_hd__and4_1 _10776_ (.A(_05050_),
    .B(_05068_),
    .C(_05098_),
    .D(_04924_),
    .X(_04928_));
 sky130_fd_sc_hd__a31o_1 _10777_ (.A1(_05050_),
    .A2(_05068_),
    .A3(_04924_),
    .B1(_05098_),
    .X(_04929_));
 sky130_fd_sc_hd__and2b_1 _10778_ (.A_N(_04928_),
    .B(_04929_),
    .X(_00044_));
 sky130_fd_sc_hd__and3_1 _10779_ (.A(_04928_),
    .B(_05107_),
    .C(_05106_),
    .X(_04931_));
 sky130_fd_sc_hd__xor2_1 _10780_ (.A(_05110_),
    .B(_04928_),
    .X(_00045_));
 sky130_fd_sc_hd__nand3b_1 _10781_ (.A_N(_05077_),
    .B(_05110_),
    .C(_04928_),
    .Y(_04932_));
 sky130_fd_sc_hd__xnor2_1 _10782_ (.A(_05077_),
    .B(_04931_),
    .Y(_00024_));
 sky130_fd_sc_hd__or3b_2 _10783_ (.A(_05077_),
    .B(_05089_),
    .C_N(_04931_),
    .X(_04933_));
 sky130_fd_sc_hd__xor2_1 _10784_ (.A(_05089_),
    .B(_04932_),
    .X(_00025_));
 sky130_fd_sc_hd__xor2_1 _10785_ (.A(_05124_),
    .B(_04933_),
    .X(_00026_));
 sky130_fd_sc_hd__or2_1 _10786_ (.A(_05124_),
    .B(_05155_),
    .X(_04934_));
 sky130_fd_sc_hd__a2bb2o_1 _10787_ (.A1_N(_05124_),
    .A2_N(_04933_),
    .B1(_05151_),
    .B2(_05150_),
    .X(_04935_));
 sky130_fd_sc_hd__o31a_1 _10788_ (.A1(_05089_),
    .A2(_04932_),
    .A3(_04934_),
    .B1(_04935_),
    .X(_00027_));
 sky130_fd_sc_hd__or4_2 _10789_ (.A(_05124_),
    .B(_05135_),
    .C(_05155_),
    .D(_04933_),
    .X(_04937_));
 sky130_fd_sc_hd__o31ai_1 _10790_ (.A1(_05124_),
    .A2(_05155_),
    .A3(_04933_),
    .B1(_05135_),
    .Y(_04938_));
 sky130_fd_sc_hd__and2_1 _10791_ (.A(_04937_),
    .B(_04938_),
    .X(_00028_));
 sky130_fd_sc_hd__xor2_1 _10792_ (.A(_05143_),
    .B(_04937_),
    .X(_00029_));
 sky130_fd_sc_hd__nor3_1 _10793_ (.A(_05143_),
    .B(_05185_),
    .C(_04937_),
    .Y(_04939_));
 sky130_fd_sc_hd__o21a_1 _10794_ (.A1(_05143_),
    .A2(_04937_),
    .B1(_05185_),
    .X(_04940_));
 sky130_fd_sc_hd__nor2_1 _10795_ (.A(_04939_),
    .B(_04940_),
    .Y(_00030_));
 sky130_fd_sc_hd__or4_1 _10796_ (.A(_05143_),
    .B(_05179_),
    .C(_05185_),
    .D(_04937_),
    .X(_04941_));
 sky130_fd_sc_hd__or2_1 _10797_ (.A(_05178_),
    .B(_04939_),
    .X(_04942_));
 sky130_fd_sc_hd__and2_1 _10798_ (.A(_04941_),
    .B(_04942_),
    .X(_00031_));
 sky130_fd_sc_hd__and3_1 _10799_ (.A(_05165_),
    .B(_05178_),
    .C(_04939_),
    .X(_04944_));
 sky130_fd_sc_hd__o41a_1 _10800_ (.A1(_05143_),
    .A2(_05179_),
    .A3(_05185_),
    .A4(_04937_),
    .B1(_05164_),
    .X(_04945_));
 sky130_fd_sc_hd__nor2_1 _10801_ (.A(_04944_),
    .B(_04945_),
    .Y(_00032_));
 sky130_fd_sc_hd__xor2_1 _10802_ (.A(_05173_),
    .B(_04944_),
    .X(_00033_));
 sky130_fd_sc_hd__or4_2 _10803_ (.A(_05164_),
    .B(_05174_),
    .C(_05210_),
    .D(_04941_),
    .X(_04946_));
 sky130_fd_sc_hd__a41o_1 _10804_ (.A1(_05165_),
    .A2(_05173_),
    .A3(_05178_),
    .A4(_04939_),
    .B1(_05211_),
    .X(_04947_));
 sky130_fd_sc_hd__and2_1 _10805_ (.A(_04946_),
    .B(_04947_),
    .X(_00035_));
 sky130_fd_sc_hd__xnor2_1 _10806_ (.A(_05205_),
    .B(_04946_),
    .Y(_00036_));
 sky130_fd_sc_hd__a41o_1 _10807_ (.A1(_05205_),
    .A2(_04944_),
    .A3(_05211_),
    .A4(_05173_),
    .B1(_01032_),
    .X(_04948_));
 sky130_fd_sc_hd__o31a_1 _10808_ (.A1(net15),
    .A2(_05204_),
    .A3(_04946_),
    .B1(_04948_),
    .X(_00037_));
 sky130_fd_sc_hd__o311a_1 _10809_ (.A1(_01252_),
    .A2(_01989_),
    .A3(net110),
    .B1(_04936_),
    .C1(_05006_),
    .X(_04950_));
 sky130_fd_sc_hd__o311a_1 _10810_ (.A1(net33),
    .A2(_01989_),
    .A3(net110),
    .B1(_05004_),
    .C1(_04949_),
    .X(_04951_));
 sky130_fd_sc_hd__nor2_1 _10811_ (.A(_04950_),
    .B(_04951_),
    .Y(_00012_));
 sky130_fd_sc_hd__or3_2 _10812_ (.A(_04949_),
    .B(\adder_inst.fraction2[0] ),
    .C(_05034_),
    .X(_04952_));
 sky130_fd_sc_hd__a31o_1 _10813_ (.A1(_04936_),
    .A2(_04943_),
    .A3(_05006_),
    .B1(_05033_),
    .X(_04953_));
 sky130_fd_sc_hd__and2_1 _10814_ (.A(_04952_),
    .B(_04953_),
    .X(_00016_));
 sky130_fd_sc_hd__xor2_1 _10815_ (.A(_04623_),
    .B(_04952_),
    .X(_00017_));
 sky130_fd_sc_hd__and4b_1 _10816_ (.A_N(_04339_),
    .B(_04612_),
    .C(_05033_),
    .D(_04950_),
    .X(_04954_));
 sky130_fd_sc_hd__o21ai_1 _10817_ (.A1(_04623_),
    .A2(_04952_),
    .B1(_04339_),
    .Y(_04955_));
 sky130_fd_sc_hd__and2b_1 _10818_ (.A_N(_04954_),
    .B(_04955_),
    .X(_00018_));
 sky130_fd_sc_hd__or4_1 _10819_ (.A(_03814_),
    .B(_04339_),
    .C(_04623_),
    .D(_04952_),
    .X(_04957_));
 sky130_fd_sc_hd__a221o_1 _10820_ (.A1(_01197_),
    .A2(_02077_),
    .B1(_03770_),
    .B2(_03792_),
    .C1(_04954_),
    .X(_04958_));
 sky130_fd_sc_hd__and2_1 _10821_ (.A(_04957_),
    .B(_04958_),
    .X(_00019_));
 sky130_fd_sc_hd__nor2_1 _10822_ (.A(_05051_),
    .B(_04957_),
    .Y(_04959_));
 sky130_fd_sc_hd__xor2_1 _10823_ (.A(_05051_),
    .B(_04957_),
    .X(_00020_));
 sky130_fd_sc_hd__or4b_1 _10824_ (.A(_03814_),
    .B(_05051_),
    .C(_05062_),
    .D_N(_04954_),
    .X(_04960_));
 sky130_fd_sc_hd__xor2_1 _10825_ (.A(_05063_),
    .B(_04959_),
    .X(_00021_));
 sky130_fd_sc_hd__and3_1 _10826_ (.A(_05063_),
    .B(_05100_),
    .C(_04959_),
    .X(_04961_));
 sky130_fd_sc_hd__xor2_1 _10827_ (.A(_05099_),
    .B(_04960_),
    .X(_00022_));
 sky130_fd_sc_hd__xor2_1 _10828_ (.A(_05112_),
    .B(_04961_),
    .X(_00023_));
 sky130_fd_sc_hd__or4_1 _10829_ (.A(_05079_),
    .B(_05099_),
    .C(_05111_),
    .D(_04960_),
    .X(_04963_));
 sky130_fd_sc_hd__a41o_1 _10830_ (.A1(_05063_),
    .A2(_05100_),
    .A3(_05112_),
    .A4(_04959_),
    .B1(_05080_),
    .X(_04964_));
 sky130_fd_sc_hd__and2_1 _10831_ (.A(_04963_),
    .B(_04964_),
    .X(_00002_));
 sky130_fd_sc_hd__xor2_1 _10832_ (.A(_05091_),
    .B(_04963_),
    .X(_00003_));
 sky130_fd_sc_hd__or3_2 _10833_ (.A(_05091_),
    .B(_05125_),
    .C(_04963_),
    .X(_04965_));
 sky130_fd_sc_hd__a41o_1 _10834_ (.A1(_05080_),
    .A2(_05092_),
    .A3(_05112_),
    .A4(_04961_),
    .B1(_05126_),
    .X(_04966_));
 sky130_fd_sc_hd__and2_1 _10835_ (.A(_04965_),
    .B(_04966_),
    .X(_00004_));
 sky130_fd_sc_hd__xor2_1 _10836_ (.A(_05148_),
    .B(_04965_),
    .X(_00005_));
 sky130_fd_sc_hd__or3_1 _10837_ (.A(_05133_),
    .B(_05148_),
    .C(_04965_),
    .X(_04967_));
 sky130_fd_sc_hd__o21ai_1 _10838_ (.A1(_05148_),
    .A2(_04965_),
    .B1(_05133_),
    .Y(_04968_));
 sky130_fd_sc_hd__and2_1 _10839_ (.A(_04967_),
    .B(_04968_),
    .X(_00006_));
 sky130_fd_sc_hd__or4_2 _10840_ (.A(_05133_),
    .B(_05140_),
    .C(_05148_),
    .D(_04965_),
    .X(_04970_));
 sky130_fd_sc_hd__nand2_1 _10841_ (.A(_05140_),
    .B(_04967_),
    .Y(_04971_));
 sky130_fd_sc_hd__and2_1 _10842_ (.A(_04970_),
    .B(_04971_),
    .X(_00007_));
 sky130_fd_sc_hd__xor2_1 _10843_ (.A(_05187_),
    .B(_04970_),
    .X(_00008_));
 sky130_fd_sc_hd__or4_2 _10844_ (.A(_05140_),
    .B(_05182_),
    .C(_05187_),
    .D(_04967_),
    .X(_04972_));
 sky130_fd_sc_hd__o21ai_1 _10845_ (.A1(_05187_),
    .A2(_04970_),
    .B1(_05182_),
    .Y(_04973_));
 sky130_fd_sc_hd__and2_1 _10846_ (.A(_04972_),
    .B(_04973_),
    .X(_00009_));
 sky130_fd_sc_hd__xor2_1 _10847_ (.A(_05163_),
    .B(_04972_),
    .X(_00010_));
 sky130_fd_sc_hd__nor3_2 _10848_ (.A(_05163_),
    .B(_05171_),
    .C(_04972_),
    .Y(_04974_));
 sky130_fd_sc_hd__o41a_1 _10849_ (.A1(_05163_),
    .A2(_05182_),
    .A3(_05187_),
    .A4(_04970_),
    .B1(_05171_),
    .X(_04976_));
 sky130_fd_sc_hd__nor2_1 _10850_ (.A(_04974_),
    .B(_04976_),
    .Y(_00011_));
 sky130_fd_sc_hd__xor2_1 _10851_ (.A(_05219_),
    .B(_04974_),
    .X(_00013_));
 sky130_fd_sc_hd__or4b_1 _10852_ (.A(_05203_),
    .B(_05214_),
    .C(_05216_),
    .D_N(_04974_),
    .X(_04977_));
 sky130_fd_sc_hd__a22o_1 _10853_ (.A1(_05201_),
    .A2(_05202_),
    .B1(_04974_),
    .B2(_05219_),
    .X(_04978_));
 sky130_fd_sc_hd__and2_1 _10854_ (.A(_04977_),
    .B(_04978_),
    .X(_00014_));
 sky130_fd_sc_hd__xor2_1 _10855_ (.A(net47),
    .B(_04977_),
    .X(_00015_));
 sky130_fd_sc_hd__dlxtn_1 _10856_ (.D(\adder_inst.fraction1[0] ),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[0] ));
 sky130_fd_sc_hd__dlxtn_1 _10857_ (.D(_00034_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[1] ));
 sky130_fd_sc_hd__dlxtn_1 _10858_ (.D(_00038_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[2] ));
 sky130_fd_sc_hd__dlxtn_1 _10859_ (.D(_00039_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[3] ));
 sky130_fd_sc_hd__dlxtn_1 _10860_ (.D(_00040_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[4] ));
 sky130_fd_sc_hd__dlxtn_1 _10861_ (.D(_00041_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[5] ));
 sky130_fd_sc_hd__dlxtn_1 _10862_ (.D(_00042_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[6] ));
 sky130_fd_sc_hd__dlxtn_1 _10863_ (.D(_00043_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[7] ));
 sky130_fd_sc_hd__dlxtn_1 _10864_ (.D(_00044_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[8] ));
 sky130_fd_sc_hd__dlxtn_1 _10865_ (.D(_00045_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[9] ));
 sky130_fd_sc_hd__dlxtn_1 _10866_ (.D(_00024_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[10] ));
 sky130_fd_sc_hd__dlxtn_1 _10867_ (.D(_00025_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[11] ));
 sky130_fd_sc_hd__dlxtn_1 _10868_ (.D(_00026_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[12] ));
 sky130_fd_sc_hd__dlxtn_2 _10869_ (.D(_00027_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[13] ));
 sky130_fd_sc_hd__dlxtn_1 _10870_ (.D(_00028_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[14] ));
 sky130_fd_sc_hd__dlxtn_1 _10871_ (.D(_00029_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[15] ));
 sky130_fd_sc_hd__dlxtn_1 _10872_ (.D(_00030_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[16] ));
 sky130_fd_sc_hd__dlxtn_1 _10873_ (.D(_00031_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[17] ));
 sky130_fd_sc_hd__dlxtn_1 _10874_ (.D(_00032_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[18] ));
 sky130_fd_sc_hd__dlxtn_2 _10875_ (.D(_00033_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[19] ));
 sky130_fd_sc_hd__dlxtn_2 _10876_ (.D(_00035_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[20] ));
 sky130_fd_sc_hd__dlxtn_1 _10877_ (.D(_00036_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[21] ));
 sky130_fd_sc_hd__dlxtn_1 _10878_ (.D(_00037_),
    .GATE_N(_00000_),
    .Q(\adder_inst.fraction1_32neg[22] ));
 sky130_fd_sc_hd__dlxtn_1 _10879_ (.D(\adder_inst.fraction2[0] ),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[0] ));
 sky130_fd_sc_hd__dlxtn_1 _10880_ (.D(_00012_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[1] ));
 sky130_fd_sc_hd__dlxtn_1 _10881_ (.D(_00016_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[2] ));
 sky130_fd_sc_hd__dlxtn_1 _10882_ (.D(_00017_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[3] ));
 sky130_fd_sc_hd__dlxtn_1 _10883_ (.D(_00018_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[4] ));
 sky130_fd_sc_hd__dlxtn_1 _10884_ (.D(_00019_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[5] ));
 sky130_fd_sc_hd__dlxtn_1 _10885_ (.D(_00020_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[6] ));
 sky130_fd_sc_hd__dlxtn_1 _10886_ (.D(_00021_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[7] ));
 sky130_fd_sc_hd__dlxtn_1 _10887_ (.D(_00022_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[8] ));
 sky130_fd_sc_hd__dlxtn_1 _10888_ (.D(_00023_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[9] ));
 sky130_fd_sc_hd__dlxtn_1 _10889_ (.D(_00002_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[10] ));
 sky130_fd_sc_hd__dlxtn_1 _10890_ (.D(_00003_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[11] ));
 sky130_fd_sc_hd__dlxtn_1 _10891_ (.D(_00004_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[12] ));
 sky130_fd_sc_hd__dlxtn_1 _10892_ (.D(_00005_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[13] ));
 sky130_fd_sc_hd__dlxtn_1 _10893_ (.D(_00006_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[14] ));
 sky130_fd_sc_hd__dlxtn_1 _10894_ (.D(_00007_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[15] ));
 sky130_fd_sc_hd__dlxtn_1 _10895_ (.D(_00008_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[16] ));
 sky130_fd_sc_hd__dlxtn_1 _10896_ (.D(_00009_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[17] ));
 sky130_fd_sc_hd__dlxtn_1 _10897_ (.D(_00010_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[18] ));
 sky130_fd_sc_hd__dlxtn_2 _10898_ (.D(_00011_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[19] ));
 sky130_fd_sc_hd__dlxtn_1 _10899_ (.D(_00013_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[20] ));
 sky130_fd_sc_hd__dlxtn_1 _10900_ (.D(_00014_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[21] ));
 sky130_fd_sc_hd__dlxtn_1 _10901_ (.D(_00015_),
    .GATE_N(_00001_),
    .Q(\adder_inst.fraction2_32neg[22] ));
 sky130_fd_sc_hd__buf_12 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_12 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_12 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_12 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_12 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_12 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_12 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_12 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_12 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_12 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_12 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_12 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_12 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_12 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_12 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_12 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_12 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_12 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_12 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_12 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_12 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_12 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_12 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_12 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_12 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_12 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_12 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_12 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_12 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_12 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_4 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_12 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_12 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_12 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_12 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_12 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_12 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_12 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_12 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_8 input65 (.A(select),
    .X(net65));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(result[0]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(result[10]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(result[11]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(result[12]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(result[13]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(result[14]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(result[15]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(result[16]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(result[17]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(result[18]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(result[19]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(result[1]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(result[20]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(result[21]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(result[22]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(result[23]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(result[24]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(result[25]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(result[26]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(result[27]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(result[28]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(result[29]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(result[2]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(result[30]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(result[31]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(result[3]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(result[4]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(result[5]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(result[6]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(result[7]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(result[8]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(result[9]));
 sky130_fd_sc_hd__buf_12 max_cap98 (.A(_03366_),
    .X(net98));
 sky130_fd_sc_hd__buf_12 max_cap99 (.A(_03366_),
    .X(net99));
 sky130_fd_sc_hd__buf_8 max_cap100 (.A(_03365_),
    .X(net100));
 sky130_fd_sc_hd__buf_8 wire101 (.A(_03364_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 max_cap102 (.A(_05231_),
    .X(net102));
 sky130_fd_sc_hd__buf_8 max_cap103 (.A(_04092_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_8 max_cap104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_16 wire105 (.A(_02066_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 max_cap106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_8 max_cap107 (.A(_02044_),
    .X(net107));
 sky130_fd_sc_hd__buf_12 max_cap108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_6 max_cap109 (.A(_02022_),
    .X(net109));
 sky130_fd_sc_hd__buf_8 wire110 (.A(_02011_),
    .X(net110));
 sky130_fd_sc_hd__buf_12 max_cap111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_6 max_cap112 (.A(_02000_),
    .X(net112));
 sky130_fd_sc_hd__buf_6 max_cap113 (.A(_01989_),
    .X(net113));
 sky130_fd_sc_hd__buf_8 max_cap114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_8 max_cap115 (.A(_05233_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_8 max_cap116 (.A(_05232_),
    .X(net116));
endmodule
