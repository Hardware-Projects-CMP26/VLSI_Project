module sequential_multiplier (clk,
    done,
    rst,
    start,
    multiplicand,
    multiplier,
    product);
 input clk;
 output done;
 input rst;
 input start;
 input [31:0] multiplicand;
 input [31:0] multiplier;
 output [63:0] product;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire \acc[0] ;
 wire \acc[10] ;
 wire \acc[11] ;
 wire \acc[12] ;
 wire \acc[13] ;
 wire \acc[14] ;
 wire \acc[15] ;
 wire \acc[16] ;
 wire \acc[17] ;
 wire \acc[18] ;
 wire \acc[19] ;
 wire \acc[1] ;
 wire \acc[20] ;
 wire \acc[21] ;
 wire \acc[22] ;
 wire \acc[23] ;
 wire \acc[24] ;
 wire \acc[25] ;
 wire \acc[26] ;
 wire \acc[27] ;
 wire \acc[28] ;
 wire \acc[29] ;
 wire \acc[2] ;
 wire \acc[30] ;
 wire \acc[31] ;
 wire \acc[32] ;
 wire \acc[33] ;
 wire \acc[34] ;
 wire \acc[35] ;
 wire \acc[36] ;
 wire \acc[37] ;
 wire \acc[38] ;
 wire \acc[39] ;
 wire \acc[3] ;
 wire \acc[40] ;
 wire \acc[41] ;
 wire \acc[42] ;
 wire \acc[43] ;
 wire \acc[44] ;
 wire \acc[45] ;
 wire \acc[46] ;
 wire \acc[47] ;
 wire \acc[48] ;
 wire \acc[49] ;
 wire \acc[4] ;
 wire \acc[50] ;
 wire \acc[51] ;
 wire \acc[52] ;
 wire \acc[53] ;
 wire \acc[54] ;
 wire \acc[55] ;
 wire \acc[56] ;
 wire \acc[57] ;
 wire \acc[58] ;
 wire \acc[59] ;
 wire \acc[5] ;
 wire \acc[60] ;
 wire \acc[61] ;
 wire \acc[62] ;
 wire \acc[63] ;
 wire \acc[6] ;
 wire \acc[7] ;
 wire \acc[8] ;
 wire \acc[9] ;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire \m[0] ;
 wire \m[10] ;
 wire \m[11] ;
 wire \m[12] ;
 wire \m[13] ;
 wire \m[14] ;
 wire \m[15] ;
 wire \m[16] ;
 wire \m[17] ;
 wire \m[18] ;
 wire \m[19] ;
 wire \m[1] ;
 wire \m[20] ;
 wire \m[21] ;
 wire \m[22] ;
 wire \m[23] ;
 wire \m[24] ;
 wire \m[25] ;
 wire \m[26] ;
 wire \m[27] ;
 wire \m[28] ;
 wire \m[29] ;
 wire \m[2] ;
 wire \m[30] ;
 wire \m[31] ;
 wire \m[3] ;
 wire \m[4] ;
 wire \m[5] ;
 wire \m[6] ;
 wire \m[7] ;
 wire \m[8] ;
 wire \m[9] ;
 wire \q[0] ;
 wire \q[10] ;
 wire \q[11] ;
 wire \q[12] ;
 wire \q[13] ;
 wire \q[14] ;
 wire \q[15] ;
 wire \q[16] ;
 wire \q[17] ;
 wire \q[18] ;
 wire \q[19] ;
 wire \q[1] ;
 wire \q[20] ;
 wire \q[21] ;
 wire \q[22] ;
 wire \q[23] ;
 wire \q[24] ;
 wire \q[25] ;
 wire \q[26] ;
 wire \q[27] ;
 wire \q[28] ;
 wire \q[29] ;
 wire \q[2] ;
 wire \q[30] ;
 wire \q[31] ;
 wire \q[3] ;
 wire \q[4] ;
 wire \q[5] ;
 wire \q[6] ;
 wire \q[7] ;
 wire \q[8] ;
 wire \q[9] ;
 wire sign;
 wire \state[0] ;
 wire \state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_2 _2035_ (.A(\q[31] ),
    .Y(_1764_));
 sky130_fd_sc_hd__inv_2 _2036_ (.A(\q[29] ),
    .Y(_1765_));
 sky130_fd_sc_hd__inv_2 _2037_ (.A(\q[28] ),
    .Y(_1766_));
 sky130_fd_sc_hd__inv_2 _2038_ (.A(\q[27] ),
    .Y(_1767_));
 sky130_fd_sc_hd__inv_2 _2039_ (.A(\q[26] ),
    .Y(_1768_));
 sky130_fd_sc_hd__inv_2 _2040_ (.A(\q[25] ),
    .Y(_1769_));
 sky130_fd_sc_hd__inv_2 _2041_ (.A(\q[23] ),
    .Y(_1770_));
 sky130_fd_sc_hd__inv_2 _2042_ (.A(\q[22] ),
    .Y(_1771_));
 sky130_fd_sc_hd__inv_2 _2043_ (.A(\q[21] ),
    .Y(_1772_));
 sky130_fd_sc_hd__inv_2 _2044_ (.A(\q[18] ),
    .Y(_1773_));
 sky130_fd_sc_hd__inv_2 _2045_ (.A(\q[17] ),
    .Y(_1774_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(\q[16] ),
    .Y(_1775_));
 sky130_fd_sc_hd__inv_2 _2047_ (.A(\q[14] ),
    .Y(_1776_));
 sky130_fd_sc_hd__inv_2 _2048_ (.A(\q[13] ),
    .Y(_1777_));
 sky130_fd_sc_hd__inv_2 _2049_ (.A(\q[12] ),
    .Y(_1778_));
 sky130_fd_sc_hd__inv_2 _2050_ (.A(\q[11] ),
    .Y(_1779_));
 sky130_fd_sc_hd__inv_2 _2051_ (.A(\q[10] ),
    .Y(_1780_));
 sky130_fd_sc_hd__inv_2 _2052_ (.A(\q[9] ),
    .Y(_1781_));
 sky130_fd_sc_hd__inv_2 _2053_ (.A(\q[8] ),
    .Y(_1782_));
 sky130_fd_sc_hd__inv_2 _2054_ (.A(\q[7] ),
    .Y(_1783_));
 sky130_fd_sc_hd__inv_2 _2055_ (.A(\q[5] ),
    .Y(_1784_));
 sky130_fd_sc_hd__inv_2 _2056_ (.A(\q[4] ),
    .Y(_1785_));
 sky130_fd_sc_hd__inv_2 _2057_ (.A(\q[2] ),
    .Y(_1786_));
 sky130_fd_sc_hd__inv_2 _2058_ (.A(\q[1] ),
    .Y(_1787_));
 sky130_fd_sc_hd__inv_2 _2059_ (.A(\acc[43] ),
    .Y(_1788_));
 sky130_fd_sc_hd__inv_2 _2060_ (.A(\acc[40] ),
    .Y(_1789_));
 sky130_fd_sc_hd__inv_2 _2061_ (.A(\acc[38] ),
    .Y(_1790_));
 sky130_fd_sc_hd__inv_2 _2062_ (.A(\acc[37] ),
    .Y(_1791_));
 sky130_fd_sc_hd__inv_2 _2063_ (.A(\acc[36] ),
    .Y(_1792_));
 sky130_fd_sc_hd__inv_2 _2064_ (.A(\acc[35] ),
    .Y(_1793_));
 sky130_fd_sc_hd__inv_2 _2065_ (.A(\acc[34] ),
    .Y(_1794_));
 sky130_fd_sc_hd__inv_2 _2066_ (.A(\acc[33] ),
    .Y(_1795_));
 sky130_fd_sc_hd__inv_2 _2067_ (.A(\acc[27] ),
    .Y(_1796_));
 sky130_fd_sc_hd__inv_2 _2068_ (.A(\acc[21] ),
    .Y(_1797_));
 sky130_fd_sc_hd__inv_2 _2069_ (.A(\acc[8] ),
    .Y(_1798_));
 sky130_fd_sc_hd__inv_2 _2070_ (.A(\acc[5] ),
    .Y(_1799_));
 sky130_fd_sc_hd__inv_2 _2071_ (.A(\acc[4] ),
    .Y(_1800_));
 sky130_fd_sc_hd__clkinv_16 _2072_ (.A(\count[5] ),
    .Y(_1801_));
 sky130_fd_sc_hd__clkinv_16 _2073_ (.A(\count[4] ),
    .Y(_1802_));
 sky130_fd_sc_hd__clkinv_16 _2074_ (.A(\count[3] ),
    .Y(_1803_));
 sky130_fd_sc_hd__clkinv_16 _2075_ (.A(net137),
    .Y(_1804_));
 sky130_fd_sc_hd__inv_16 _2076_ (.A(\count[1] ),
    .Y(_1805_));
 sky130_fd_sc_hd__inv_4 _2077_ (.A(net140),
    .Y(_1806_));
 sky130_fd_sc_hd__inv_4 _2078_ (.A(net57),
    .Y(_1807_));
 sky130_fd_sc_hd__inv_2 _2079_ (.A(net58),
    .Y(_1808_));
 sky130_fd_sc_hd__inv_2 _2080_ (.A(net59),
    .Y(_1809_));
 sky130_fd_sc_hd__inv_2 _2081_ (.A(net61),
    .Y(_1810_));
 sky130_fd_sc_hd__inv_2 _2082_ (.A(net35),
    .Y(_1811_));
 sky130_fd_sc_hd__inv_2 _2083_ (.A(net38),
    .Y(_1812_));
 sky130_fd_sc_hd__inv_2 _2084_ (.A(net42),
    .Y(_1813_));
 sky130_fd_sc_hd__inv_2 _2085_ (.A(net10),
    .Y(_1814_));
 sky130_fd_sc_hd__inv_2 _2086_ (.A(net15),
    .Y(_1815_));
 sky130_fd_sc_hd__inv_2 _2087_ (.A(net65),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2b_4 _2088_ (.A_N(\state[0] ),
    .B(net66),
    .Y(_1816_));
 sky130_fd_sc_hd__nor2_8 _2089_ (.A(\state[1] ),
    .B(_1816_),
    .Y(_1817_));
 sky130_fd_sc_hd__or3b_4 _2090_ (.A(\state[1] ),
    .B(\state[0] ),
    .C_N(net66),
    .X(_1818_));
 sky130_fd_sc_hd__or2_1 _2091_ (.A(net1),
    .B(net12),
    .X(_1819_));
 sky130_fd_sc_hd__or3_1 _2092_ (.A(net1),
    .B(net12),
    .C(net23),
    .X(_1820_));
 sky130_fd_sc_hd__nor4_1 _2093_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(net26),
    .Y(_1821_));
 sky130_fd_sc_hd__or4_1 _2094_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(net26),
    .X(_1822_));
 sky130_fd_sc_hd__or4_2 _2095_ (.A(net23),
    .B(net26),
    .C(net27),
    .D(_1819_),
    .X(_1823_));
 sky130_fd_sc_hd__nor2_1 _2096_ (.A(net28),
    .B(net29),
    .Y(_1824_));
 sky130_fd_sc_hd__nand3b_2 _2097_ (.A_N(net27),
    .B(_1821_),
    .C(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__or2_1 _2098_ (.A(net30),
    .B(net31),
    .X(_1826_));
 sky130_fd_sc_hd__or4_1 _2099_ (.A(net28),
    .B(_1826_),
    .C(net29),
    .D(_1823_),
    .X(_1827_));
 sky130_fd_sc_hd__nor4_1 _2100_ (.A(net32),
    .B(_1826_),
    .C(net2),
    .D(_1825_),
    .Y(_1828_));
 sky130_fd_sc_hd__or4_2 _2101_ (.A(net32),
    .B(_1826_),
    .C(net2),
    .D(_1825_),
    .X(_1829_));
 sky130_fd_sc_hd__or2_1 _2102_ (.A(net3),
    .B(net4),
    .X(_1830_));
 sky130_fd_sc_hd__nor4b_1 _2103_ (.A(net5),
    .B(_1830_),
    .C(net6),
    .D_N(_1828_),
    .Y(_1831_));
 sky130_fd_sc_hd__or4_2 _2104_ (.A(net5),
    .B(_1830_),
    .C(net6),
    .D(_1829_),
    .X(_1832_));
 sky130_fd_sc_hd__nor2_1 _2105_ (.A(net7),
    .B(net8),
    .Y(_1833_));
 sky130_fd_sc_hd__or3_1 _2106_ (.A(net7),
    .B(net8),
    .C(_1832_),
    .X(_1834_));
 sky130_fd_sc_hd__nand4b_4 _2107_ (.A_N(net9),
    .B(_1831_),
    .C(_1833_),
    .D(_1814_),
    .Y(_1835_));
 sky130_fd_sc_hd__or3_1 _2108_ (.A(net11),
    .B(net13),
    .C(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__nor4_1 _2109_ (.A(net11),
    .B(net13),
    .C(net14),
    .D(_1835_),
    .Y(_1837_));
 sky130_fd_sc_hd__nand2_1 _2110_ (.A(_1837_),
    .B(_1815_),
    .Y(_1838_));
 sky130_fd_sc_hd__or3_1 _2111_ (.A(net16),
    .B(net17),
    .C(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__or3_1 _2112_ (.A(net18),
    .B(net19),
    .C(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__or3_1 _2113_ (.A(net20),
    .B(net21),
    .C(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__or4_1 _2114_ (.A(net20),
    .B(net21),
    .C(net22),
    .D(_1840_),
    .X(_1842_));
 sky130_fd_sc_hd__or4b_1 _2115_ (.A(\state[1] ),
    .B(net24),
    .C(_1816_),
    .D_N(net25),
    .X(_1843_));
 sky130_fd_sc_hd__a2bb2o_1 _2116_ (.A1_N(_1842_),
    .A2_N(_1843_),
    .B1(\q[31] ),
    .B2(_1818_),
    .X(_0403_));
 sky130_fd_sc_hd__o2111ai_1 _2117_ (.A1(net22),
    .A2(_1841_),
    .B1(net24),
    .C1(net25),
    .D1(_1817_),
    .Y(_1844_));
 sky130_fd_sc_hd__a211o_1 _2118_ (.A1(_1842_),
    .A2(net25),
    .B1(net24),
    .C1(_1818_),
    .X(_1845_));
 sky130_fd_sc_hd__o211a_1 _2119_ (.A1(\q[30] ),
    .A2(_1817_),
    .B1(_1844_),
    .C1(_1845_),
    .X(_0402_));
 sky130_fd_sc_hd__o311a_1 _2120_ (.A1(net20),
    .A2(net21),
    .A3(_1840_),
    .B1(net22),
    .C1(net25),
    .X(_1846_));
 sky130_fd_sc_hd__a21oi_1 _2121_ (.A1(_1841_),
    .A2(net25),
    .B1(net22),
    .Y(_1847_));
 sky130_fd_sc_hd__or3_1 _2122_ (.A(_1818_),
    .B(_1846_),
    .C(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__o21ai_1 _2123_ (.A1(_1765_),
    .A2(_1817_),
    .B1(_1848_),
    .Y(_0401_));
 sky130_fd_sc_hd__o41a_1 _2124_ (.A1(net18),
    .A2(net19),
    .A3(net20),
    .A4(_1839_),
    .B1(net25),
    .X(_1849_));
 sky130_fd_sc_hd__o211a_1 _2125_ (.A1(net20),
    .A2(_1840_),
    .B1(net21),
    .C1(net25),
    .X(_1850_));
 sky130_fd_sc_hd__nor2_1 _2126_ (.A(net21),
    .B(_1849_),
    .Y(_1851_));
 sky130_fd_sc_hd__or4_1 _2127_ (.A(\state[1] ),
    .B(_1816_),
    .C(_1850_),
    .D(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__o21ai_1 _2128_ (.A1(_1766_),
    .A2(_1817_),
    .B1(_1852_),
    .Y(_0400_));
 sky130_fd_sc_hd__o311a_1 _2129_ (.A1(net18),
    .A2(net19),
    .A3(_1839_),
    .B1(net20),
    .C1(net25),
    .X(_1853_));
 sky130_fd_sc_hd__a21oi_1 _2130_ (.A1(_1840_),
    .A2(net25),
    .B1(net20),
    .Y(_1854_));
 sky130_fd_sc_hd__or4_1 _2131_ (.A(\state[1] ),
    .B(_1816_),
    .C(_1853_),
    .D(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__o21ai_1 _2132_ (.A1(_1767_),
    .A2(_1817_),
    .B1(_1855_),
    .Y(_0399_));
 sky130_fd_sc_hd__o41a_1 _2133_ (.A1(net16),
    .A2(net17),
    .A3(net18),
    .A4(_1838_),
    .B1(net25),
    .X(_1856_));
 sky130_fd_sc_hd__xor2_1 _2134_ (.A(net19),
    .B(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__mux2_1 _2135_ (.A0(_1857_),
    .A1(\q[26] ),
    .S(_1818_),
    .X(_0398_));
 sky130_fd_sc_hd__o311a_1 _2136_ (.A1(net16),
    .A2(net17),
    .A3(_1838_),
    .B1(net18),
    .C1(net25),
    .X(_1858_));
 sky130_fd_sc_hd__a21oi_1 _2137_ (.A1(_1839_),
    .A2(net25),
    .B1(net18),
    .Y(_1859_));
 sky130_fd_sc_hd__or4_1 _2138_ (.A(\state[1] ),
    .B(_1816_),
    .C(_1858_),
    .D(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__o21ai_1 _2139_ (.A1(_1769_),
    .A2(_1817_),
    .B1(_1860_),
    .Y(_0397_));
 sky130_fd_sc_hd__o21ai_1 _2140_ (.A1(net16),
    .A2(_1838_),
    .B1(net25),
    .Y(_1861_));
 sky130_fd_sc_hd__xnor2_1 _2141_ (.A(net17),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__mux2_1 _2142_ (.A0(_1862_),
    .A1(\q[24] ),
    .S(_1818_),
    .X(_0396_));
 sky130_fd_sc_hd__o311a_1 _2143_ (.A1(net14),
    .A2(net15),
    .A3(_1836_),
    .B1(net16),
    .C1(net25),
    .X(_1863_));
 sky130_fd_sc_hd__a21oi_1 _2144_ (.A1(_1838_),
    .A2(net25),
    .B1(net16),
    .Y(_1864_));
 sky130_fd_sc_hd__or4_1 _2145_ (.A(\state[1] ),
    .B(_1864_),
    .C(_1816_),
    .D(_1863_),
    .X(_1865_));
 sky130_fd_sc_hd__o21ai_1 _2146_ (.A1(_1770_),
    .A2(_1817_),
    .B1(_1865_),
    .Y(_0395_));
 sky130_fd_sc_hd__o41a_1 _2147_ (.A1(net11),
    .A2(net13),
    .A3(net14),
    .A4(_1835_),
    .B1(net25),
    .X(_1866_));
 sky130_fd_sc_hd__xor2_1 _2148_ (.A(net15),
    .B(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_1 _2149_ (.A0(_1867_),
    .A1(\q[22] ),
    .S(_1818_),
    .X(_0394_));
 sky130_fd_sc_hd__o311a_1 _2150_ (.A1(net11),
    .A2(net13),
    .A3(_1835_),
    .B1(net14),
    .C1(net25),
    .X(_1868_));
 sky130_fd_sc_hd__a21oi_1 _2151_ (.A1(_1836_),
    .A2(net25),
    .B1(net14),
    .Y(_1869_));
 sky130_fd_sc_hd__o21ai_1 _2152_ (.A1(\state[1] ),
    .A2(_1816_),
    .B1(\q[21] ),
    .Y(_1870_));
 sky130_fd_sc_hd__o31ai_1 _2153_ (.A1(_1818_),
    .A2(_1868_),
    .A3(_1869_),
    .B1(_1870_),
    .Y(_0393_));
 sky130_fd_sc_hd__o21ai_1 _2154_ (.A1(net11),
    .A2(_1835_),
    .B1(net25),
    .Y(_1871_));
 sky130_fd_sc_hd__xnor2_1 _2155_ (.A(net13),
    .B(_1871_),
    .Y(_1872_));
 sky130_fd_sc_hd__mux2_1 _2156_ (.A0(_1872_),
    .A1(\q[20] ),
    .S(_1818_),
    .X(_0392_));
 sky130_fd_sc_hd__o311a_1 _2157_ (.A1(net9),
    .A2(net10),
    .A3(_1834_),
    .B1(net11),
    .C1(net25),
    .X(_1873_));
 sky130_fd_sc_hd__a21oi_1 _2158_ (.A1(_1835_),
    .A2(net25),
    .B1(net11),
    .Y(_1874_));
 sky130_fd_sc_hd__or4_1 _2159_ (.A(\state[1] ),
    .B(_1874_),
    .C(_1816_),
    .D(_1873_),
    .X(_1875_));
 sky130_fd_sc_hd__a21bo_1 _2160_ (.A1(\q[19] ),
    .A2(_1818_),
    .B1_N(_1875_),
    .X(_0391_));
 sky130_fd_sc_hd__o41a_1 _2161_ (.A1(net7),
    .A2(net8),
    .A3(net9),
    .A4(_1832_),
    .B1(net25),
    .X(_1876_));
 sky130_fd_sc_hd__xor2_1 _2162_ (.A(net10),
    .B(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__mux2_1 _2163_ (.A0(_1877_),
    .A1(\q[18] ),
    .S(_1818_),
    .X(_0390_));
 sky130_fd_sc_hd__o311a_1 _2164_ (.A1(net7),
    .A2(net8),
    .A3(_1832_),
    .B1(net9),
    .C1(net25),
    .X(_1878_));
 sky130_fd_sc_hd__a21oi_1 _2165_ (.A1(_1834_),
    .A2(net25),
    .B1(net9),
    .Y(_1879_));
 sky130_fd_sc_hd__o21ai_1 _2166_ (.A1(\state[1] ),
    .A2(_1816_),
    .B1(\q[17] ),
    .Y(_1880_));
 sky130_fd_sc_hd__o31ai_1 _2167_ (.A1(_1818_),
    .A2(_1878_),
    .A3(_1879_),
    .B1(_1880_),
    .Y(_0389_));
 sky130_fd_sc_hd__o21ai_1 _2168_ (.A1(net7),
    .A2(_1832_),
    .B1(net25),
    .Y(_1881_));
 sky130_fd_sc_hd__xnor2_1 _2169_ (.A(net8),
    .B(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__mux2_1 _2170_ (.A0(_1882_),
    .A1(\q[16] ),
    .S(_1818_),
    .X(_0388_));
 sky130_fd_sc_hd__and3_1 _2171_ (.A(_1832_),
    .B(net7),
    .C(net25),
    .X(_1883_));
 sky130_fd_sc_hd__a21oi_1 _2172_ (.A1(_1832_),
    .A2(net25),
    .B1(net7),
    .Y(_1884_));
 sky130_fd_sc_hd__or4_1 _2173_ (.A(\state[1] ),
    .B(_1884_),
    .C(_1816_),
    .D(_1883_),
    .X(_1885_));
 sky130_fd_sc_hd__a21bo_1 _2174_ (.A1(\q[15] ),
    .A2(_1818_),
    .B1_N(_1885_),
    .X(_0387_));
 sky130_fd_sc_hd__o31a_1 _2175_ (.A1(_1830_),
    .A2(net5),
    .A3(_1829_),
    .B1(net25),
    .X(_1886_));
 sky130_fd_sc_hd__xor2_1 _2176_ (.A(net6),
    .B(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__mux2_1 _2177_ (.A0(_1887_),
    .A1(\q[14] ),
    .S(_1818_),
    .X(_0386_));
 sky130_fd_sc_hd__o31a_1 _2178_ (.A1(net3),
    .A2(net4),
    .A3(_1829_),
    .B1(net25),
    .X(_1888_));
 sky130_fd_sc_hd__xor2_1 _2179_ (.A(net5),
    .B(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__mux2_1 _2180_ (.A0(_1889_),
    .A1(\q[13] ),
    .S(_1818_),
    .X(_0385_));
 sky130_fd_sc_hd__o21ai_1 _2181_ (.A1(net3),
    .A2(_1829_),
    .B1(net25),
    .Y(_1890_));
 sky130_fd_sc_hd__xnor2_1 _2182_ (.A(net4),
    .B(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__mux2_1 _2183_ (.A0(_1891_),
    .A1(\q[12] ),
    .S(_1818_),
    .X(_0384_));
 sky130_fd_sc_hd__o311a_1 _2184_ (.A1(net32),
    .A2(net2),
    .A3(_1827_),
    .B1(net3),
    .C1(net25),
    .X(_1892_));
 sky130_fd_sc_hd__a21oi_1 _2185_ (.A1(_1829_),
    .A2(net25),
    .B1(net3),
    .Y(_1893_));
 sky130_fd_sc_hd__or4_1 _2186_ (.A(\state[1] ),
    .B(_1893_),
    .C(_1816_),
    .D(_1892_),
    .X(_1894_));
 sky130_fd_sc_hd__o21ai_1 _2187_ (.A1(_1779_),
    .A2(_1817_),
    .B1(_1894_),
    .Y(_0383_));
 sky130_fd_sc_hd__o31a_1 _2188_ (.A1(_1826_),
    .A2(net32),
    .A3(_1825_),
    .B1(net25),
    .X(_1895_));
 sky130_fd_sc_hd__xor2_1 _2189_ (.A(net2),
    .B(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__mux2_1 _2190_ (.A0(_1896_),
    .A1(\q[10] ),
    .S(_1818_),
    .X(_0382_));
 sky130_fd_sc_hd__o311a_1 _2191_ (.A1(net30),
    .A2(net31),
    .A3(_1825_),
    .B1(net32),
    .C1(net25),
    .X(_1897_));
 sky130_fd_sc_hd__a21oi_1 _2192_ (.A1(_1827_),
    .A2(net25),
    .B1(net32),
    .Y(_1898_));
 sky130_fd_sc_hd__or4_1 _2193_ (.A(\state[1] ),
    .B(_1816_),
    .C(_1897_),
    .D(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__o21ai_1 _2194_ (.A1(_1781_),
    .A2(_1817_),
    .B1(_1899_),
    .Y(_0381_));
 sky130_fd_sc_hd__o41a_1 _2195_ (.A1(net28),
    .A2(net29),
    .A3(net30),
    .A4(_1823_),
    .B1(net25),
    .X(_1900_));
 sky130_fd_sc_hd__xor2_1 _2196_ (.A(net31),
    .B(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(_1901_),
    .A1(\q[8] ),
    .S(_1818_),
    .X(_0380_));
 sky130_fd_sc_hd__o311a_1 _2198_ (.A1(net28),
    .A2(net29),
    .A3(_1823_),
    .B1(net30),
    .C1(net25),
    .X(_1902_));
 sky130_fd_sc_hd__a21oi_1 _2199_ (.A1(_1825_),
    .A2(net25),
    .B1(net30),
    .Y(_1903_));
 sky130_fd_sc_hd__or4_1 _2200_ (.A(\state[1] ),
    .B(_1903_),
    .C(_1816_),
    .D(_1902_),
    .X(_1904_));
 sky130_fd_sc_hd__o21ai_1 _2201_ (.A1(_1783_),
    .A2(_1817_),
    .B1(_1904_),
    .Y(_0379_));
 sky130_fd_sc_hd__o21ai_1 _2202_ (.A1(net28),
    .A2(_1823_),
    .B1(net25),
    .Y(_1905_));
 sky130_fd_sc_hd__xnor2_1 _2203_ (.A(net29),
    .B(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__mux2_1 _2204_ (.A0(_1906_),
    .A1(\q[6] ),
    .S(_1818_),
    .X(_0378_));
 sky130_fd_sc_hd__o311a_1 _2205_ (.A1(net26),
    .A2(net27),
    .A3(_1820_),
    .B1(net28),
    .C1(net25),
    .X(_1907_));
 sky130_fd_sc_hd__a21oi_1 _2206_ (.A1(_1823_),
    .A2(net25),
    .B1(net28),
    .Y(_1908_));
 sky130_fd_sc_hd__o21ai_1 _2207_ (.A1(\state[1] ),
    .A2(_1816_),
    .B1(\q[5] ),
    .Y(_1909_));
 sky130_fd_sc_hd__o31ai_1 _2208_ (.A1(_1818_),
    .A2(_1907_),
    .A3(_1908_),
    .B1(_1909_),
    .Y(_0377_));
 sky130_fd_sc_hd__o311a_1 _2209_ (.A1(net23),
    .A2(net26),
    .A3(_1819_),
    .B1(net27),
    .C1(net25),
    .X(_1910_));
 sky130_fd_sc_hd__a21oi_1 _2210_ (.A1(_1822_),
    .A2(net25),
    .B1(net27),
    .Y(_1911_));
 sky130_fd_sc_hd__or4_1 _2211_ (.A(\state[1] ),
    .B(_1816_),
    .C(_1910_),
    .D(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__o21ai_1 _2212_ (.A1(_1785_),
    .A2(_1817_),
    .B1(_1912_),
    .Y(_0376_));
 sky130_fd_sc_hd__o311a_1 _2213_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .B1(net26),
    .C1(net25),
    .X(_1913_));
 sky130_fd_sc_hd__a21oi_1 _2214_ (.A1(_1820_),
    .A2(net25),
    .B1(net26),
    .Y(_1914_));
 sky130_fd_sc_hd__or4_1 _2215_ (.A(\state[1] ),
    .B(_1816_),
    .C(_1913_),
    .D(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__a21bo_1 _2216_ (.A1(\q[3] ),
    .A2(_1818_),
    .B1_N(_1915_),
    .X(_0375_));
 sky130_fd_sc_hd__and3_1 _2217_ (.A(_1819_),
    .B(net23),
    .C(net25),
    .X(_1916_));
 sky130_fd_sc_hd__a21oi_1 _2218_ (.A1(_1819_),
    .A2(net25),
    .B1(net23),
    .Y(_1917_));
 sky130_fd_sc_hd__or4_1 _2219_ (.A(\state[1] ),
    .B(_1917_),
    .C(_1816_),
    .D(_1916_),
    .X(_1918_));
 sky130_fd_sc_hd__o21ai_1 _2220_ (.A1(_1786_),
    .A2(_1817_),
    .B1(_1918_),
    .Y(_0374_));
 sky130_fd_sc_hd__and3_1 _2221_ (.A(net1),
    .B(net12),
    .C(net25),
    .X(_1919_));
 sky130_fd_sc_hd__a21oi_1 _2222_ (.A1(net1),
    .A2(net25),
    .B1(net12),
    .Y(_1920_));
 sky130_fd_sc_hd__or4_1 _2223_ (.A(\state[1] ),
    .B(_1920_),
    .C(_1816_),
    .D(_1919_),
    .X(_1921_));
 sky130_fd_sc_hd__o21ai_1 _2224_ (.A1(_1787_),
    .A2(_1817_),
    .B1(_1921_),
    .Y(_0373_));
 sky130_fd_sc_hd__mux2_1 _2225_ (.A0(\q[0] ),
    .A1(net1),
    .S(_1817_),
    .X(_0372_));
 sky130_fd_sc_hd__and2b_4 _2226_ (.A_N(\state[1] ),
    .B(\state[0] ),
    .X(_1922_));
 sky130_fd_sc_hd__nand2b_4 _2227_ (.A_N(\state[1] ),
    .B(\state[0] ),
    .Y(_1923_));
 sky130_fd_sc_hd__nor2_8 _2228_ (.A(net135),
    .B(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__o22a_4 _2229_ (.A1(\state[1] ),
    .A2(_1816_),
    .B1(_1923_),
    .B2(\count[5] ),
    .X(_1925_));
 sky130_fd_sc_hd__inv_2 _2230_ (.A(_1925_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor3_1 _2231_ (.A(net33),
    .B(net44),
    .C(net55),
    .Y(_1926_));
 sky130_fd_sc_hd__or3_1 _2232_ (.A(net33),
    .B(net44),
    .C(net55),
    .X(_1927_));
 sky130_fd_sc_hd__or3_1 _2233_ (.A(net58),
    .B(net59),
    .C(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__or4_1 _2234_ (.A(net58),
    .B(net59),
    .C(net60),
    .D(_1927_),
    .X(_1929_));
 sky130_fd_sc_hd__nor2_1 _2235_ (.A(net60),
    .B(net61),
    .Y(_1930_));
 sky130_fd_sc_hd__and4_1 _2236_ (.A(_1926_),
    .B(_1930_),
    .C(_1808_),
    .D(_1809_),
    .X(_1931_));
 sky130_fd_sc_hd__or4_1 _2237_ (.A(net60),
    .B(net61),
    .C(net62),
    .D(_1928_),
    .X(_1932_));
 sky130_fd_sc_hd__nor2_1 _2238_ (.A(net62),
    .B(net63),
    .Y(_1933_));
 sky130_fd_sc_hd__and4bb_1 _2239_ (.A_N(net64),
    .B_N(_1928_),
    .C(_1930_),
    .D(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__nor2_1 _2240_ (.A(net64),
    .B(net34),
    .Y(_1935_));
 sky130_fd_sc_hd__or4_1 _2241_ (.A(net63),
    .B(net64),
    .C(net34),
    .D(_1932_),
    .X(_1936_));
 sky130_fd_sc_hd__nand4_2 _2242_ (.A(_1931_),
    .B(_1933_),
    .C(_1935_),
    .D(_1811_),
    .Y(_1937_));
 sky130_fd_sc_hd__nor2_1 _2243_ (.A(net36),
    .B(net37),
    .Y(_1938_));
 sky130_fd_sc_hd__or3_1 _2244_ (.A(net36),
    .B(net37),
    .C(_1937_),
    .X(_1939_));
 sky130_fd_sc_hd__and4b_1 _2245_ (.A_N(_1936_),
    .B(_1938_),
    .C(_1811_),
    .D(_1812_),
    .X(_1940_));
 sky130_fd_sc_hd__nor4b_2 _2246_ (.A(net38),
    .B(net39),
    .C(_1937_),
    .D_N(_1938_),
    .Y(_1941_));
 sky130_fd_sc_hd__nor2_1 _2247_ (.A(net40),
    .B(net41),
    .Y(_1942_));
 sky130_fd_sc_hd__or4b_1 _2248_ (.A(net38),
    .B(net39),
    .C(_1939_),
    .D_N(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__nor2_1 _2249_ (.A(net43),
    .B(net45),
    .Y(_1944_));
 sky130_fd_sc_hd__nand4_2 _2250_ (.A(_1941_),
    .B(_1942_),
    .C(_1944_),
    .D(_1813_),
    .Y(_1945_));
 sky130_fd_sc_hd__nor3_1 _2251_ (.A(net46),
    .B(net47),
    .C(_1945_),
    .Y(_1946_));
 sky130_fd_sc_hd__nor4_1 _2252_ (.A(net46),
    .B(net47),
    .C(net48),
    .D(_1945_),
    .Y(_1947_));
 sky130_fd_sc_hd__or3b_1 _2253_ (.A(net48),
    .B(net49),
    .C_N(_1946_),
    .X(_1948_));
 sky130_fd_sc_hd__or3_2 _2254_ (.A(net50),
    .B(net51),
    .C(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__nor2_1 _2255_ (.A(net52),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nor4_1 _2256_ (.A(net52),
    .B(net53),
    .C(net54),
    .D(_1949_),
    .Y(_1951_));
 sky130_fd_sc_hd__and4b_1 _2257_ (.A_N(net56),
    .B(_1817_),
    .C(_1951_),
    .D(net57),
    .X(_1952_));
 sky130_fd_sc_hd__a21o_1 _2258_ (.A1(\m[31] ),
    .A2(_1925_),
    .B1(_1952_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _2259_ (.A(_1807_),
    .B(_1951_),
    .X(_1953_));
 sky130_fd_sc_hd__a21oi_1 _2260_ (.A1(_1953_),
    .A2(net56),
    .B1(_1922_),
    .Y(_1954_));
 sky130_fd_sc_hd__o21ai_1 _2261_ (.A1(net56),
    .A2(_1953_),
    .B1(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__o22a_1 _2262_ (.A1(\m[31] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .X(_1956_));
 sky130_fd_sc_hd__a22o_1 _2263_ (.A1(\m[30] ),
    .A2(_1925_),
    .B1(_1955_),
    .B2(_1956_),
    .X(_0370_));
 sky130_fd_sc_hd__o31ai_1 _2264_ (.A1(net52),
    .A2(net53),
    .A3(_1949_),
    .B1(net57),
    .Y(_1957_));
 sky130_fd_sc_hd__a21oi_1 _2265_ (.A1(_1957_),
    .A2(net54),
    .B1(_1922_),
    .Y(_1958_));
 sky130_fd_sc_hd__o21ai_1 _2266_ (.A1(net54),
    .A2(_1957_),
    .B1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__o221a_1 _2267_ (.A1(\m[30] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_1959_),
    .X(_1960_));
 sky130_fd_sc_hd__a21o_1 _2268_ (.A1(\m[29] ),
    .A2(_1925_),
    .B1(_1960_),
    .X(_0369_));
 sky130_fd_sc_hd__nor2_1 _2269_ (.A(net53),
    .B(_1950_),
    .Y(_1961_));
 sky130_fd_sc_hd__o21a_1 _2270_ (.A1(_1807_),
    .A2(_1950_),
    .B1(net53),
    .X(_1962_));
 sky130_fd_sc_hd__a211o_1 _2271_ (.A1(net57),
    .A2(_1961_),
    .B1(_1962_),
    .C1(_1922_),
    .X(_1963_));
 sky130_fd_sc_hd__o221a_1 _2272_ (.A1(\m[29] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__a21o_1 _2273_ (.A1(\m[28] ),
    .A2(_1925_),
    .B1(_1964_),
    .X(_0368_));
 sky130_fd_sc_hd__or3b_1 _2274_ (.A(_1807_),
    .B(net52),
    .C_N(_1949_),
    .X(_1965_));
 sky130_fd_sc_hd__a21bo_1 _2275_ (.A1(_1949_),
    .A2(net57),
    .B1_N(net52),
    .X(_1966_));
 sky130_fd_sc_hd__and3_1 _2276_ (.A(_1923_),
    .B(_1965_),
    .C(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__o21ai_1 _2277_ (.A1(\m[28] ),
    .A2(_1923_),
    .B1(_0274_),
    .Y(_1968_));
 sky130_fd_sc_hd__a2bb2o_1 _2278_ (.A1_N(_1968_),
    .A2_N(_1967_),
    .B1(_1925_),
    .B2(\m[27] ),
    .X(_0367_));
 sky130_fd_sc_hd__o21ai_1 _2279_ (.A1(net50),
    .A2(_1948_),
    .B1(net57),
    .Y(_1969_));
 sky130_fd_sc_hd__a21oi_1 _2280_ (.A1(_1969_),
    .A2(net51),
    .B1(_1922_),
    .Y(_1970_));
 sky130_fd_sc_hd__o21ai_1 _2281_ (.A1(net51),
    .A2(_1969_),
    .B1(_1970_),
    .Y(_1971_));
 sky130_fd_sc_hd__o221a_1 _2282_ (.A1(\m[27] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__a21o_1 _2283_ (.A1(\m[26] ),
    .A2(_1925_),
    .B1(_1972_),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _2284_ (.A(_1948_),
    .B(net57),
    .Y(_1973_));
 sky130_fd_sc_hd__a21oi_1 _2285_ (.A1(_1973_),
    .A2(net50),
    .B1(_1922_),
    .Y(_1974_));
 sky130_fd_sc_hd__o21ai_1 _2286_ (.A1(net50),
    .A2(_1973_),
    .B1(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__o221a_1 _2287_ (.A1(\m[26] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__a21o_1 _2288_ (.A1(\m[25] ),
    .A2(_1925_),
    .B1(_1976_),
    .X(_0365_));
 sky130_fd_sc_hd__or3_1 _2289_ (.A(_1807_),
    .B(net49),
    .C(_1947_),
    .X(_1977_));
 sky130_fd_sc_hd__o21ai_1 _2290_ (.A1(_1807_),
    .A2(_1947_),
    .B1(net49),
    .Y(_1978_));
 sky130_fd_sc_hd__and3_1 _2291_ (.A(_1923_),
    .B(_1977_),
    .C(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__o21ai_1 _2292_ (.A1(\m[25] ),
    .A2(_1923_),
    .B1(_0274_),
    .Y(_1980_));
 sky130_fd_sc_hd__a2bb2o_1 _2293_ (.A1_N(_1980_),
    .A2_N(_1979_),
    .B1(_1925_),
    .B2(\m[24] ),
    .X(_0364_));
 sky130_fd_sc_hd__o21ai_1 _2294_ (.A1(_1807_),
    .A2(_1946_),
    .B1(net48),
    .Y(_1981_));
 sky130_fd_sc_hd__o31a_1 _2295_ (.A1(_1807_),
    .A2(net48),
    .A3(_1946_),
    .B1(_1923_),
    .X(_1982_));
 sky130_fd_sc_hd__o2bb2a_1 _2296_ (.A1_N(_1982_),
    .A2_N(_1981_),
    .B1(_1923_),
    .B2(\m[24] ),
    .X(_1983_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(_1983_),
    .A1(\m[23] ),
    .S(_1925_),
    .X(_0363_));
 sky130_fd_sc_hd__o21ai_1 _2298_ (.A1(net46),
    .A2(_1945_),
    .B1(net57),
    .Y(_1984_));
 sky130_fd_sc_hd__a21oi_1 _2299_ (.A1(_1984_),
    .A2(net47),
    .B1(_1922_),
    .Y(_1985_));
 sky130_fd_sc_hd__o21ai_1 _2300_ (.A1(net47),
    .A2(_1984_),
    .B1(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__o221a_1 _2301_ (.A1(\m[23] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__a21o_1 _2302_ (.A1(\m[22] ),
    .A2(_1925_),
    .B1(_1987_),
    .X(_0362_));
 sky130_fd_sc_hd__a41o_1 _2303_ (.A1(_1941_),
    .A2(_1942_),
    .A3(_1944_),
    .A4(_1813_),
    .B1(_1807_),
    .X(_1988_));
 sky130_fd_sc_hd__a21oi_1 _2304_ (.A1(_1988_),
    .A2(net46),
    .B1(_1922_),
    .Y(_1989_));
 sky130_fd_sc_hd__o21ai_1 _2305_ (.A1(net46),
    .A2(_1988_),
    .B1(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__o22a_1 _2306_ (.A1(\m[22] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .X(_1991_));
 sky130_fd_sc_hd__a22o_1 _2307_ (.A1(\m[21] ),
    .A2(_1925_),
    .B1(_1990_),
    .B2(_1991_),
    .X(_0361_));
 sky130_fd_sc_hd__o31ai_1 _2308_ (.A1(net42),
    .A2(net43),
    .A3(_1943_),
    .B1(net57),
    .Y(_1992_));
 sky130_fd_sc_hd__a21oi_1 _2309_ (.A1(_1992_),
    .A2(net45),
    .B1(_1922_),
    .Y(_1993_));
 sky130_fd_sc_hd__o21ai_1 _2310_ (.A1(net45),
    .A2(_1992_),
    .B1(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__o221a_1 _2311_ (.A1(\m[21] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__a21o_1 _2312_ (.A1(\m[20] ),
    .A2(_1925_),
    .B1(_1995_),
    .X(_0360_));
 sky130_fd_sc_hd__a31o_1 _2313_ (.A1(_1941_),
    .A2(_1942_),
    .A3(_1813_),
    .B1(_1807_),
    .X(_1996_));
 sky130_fd_sc_hd__a21oi_1 _2314_ (.A1(_1996_),
    .A2(net43),
    .B1(_1922_),
    .Y(_1997_));
 sky130_fd_sc_hd__o21ai_1 _2315_ (.A1(net43),
    .A2(_1996_),
    .B1(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__o22a_1 _2316_ (.A1(\m[20] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .X(_1999_));
 sky130_fd_sc_hd__a22o_1 _2317_ (.A1(\m[19] ),
    .A2(_1925_),
    .B1(_1998_),
    .B2(_1999_),
    .X(_0359_));
 sky130_fd_sc_hd__a21oi_1 _2318_ (.A1(_1943_),
    .A2(net57),
    .B1(_1813_),
    .Y(_2000_));
 sky130_fd_sc_hd__a31o_1 _2319_ (.A1(_1943_),
    .A2(net57),
    .A3(_1813_),
    .B1(_1922_),
    .X(_2001_));
 sky130_fd_sc_hd__o22a_1 _2320_ (.A1(\m[19] ),
    .A2(_1923_),
    .B1(_2000_),
    .B2(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _2321_ (.A0(_2002_),
    .A1(\m[18] ),
    .S(_1925_),
    .X(_0358_));
 sky130_fd_sc_hd__o41a_1 _2322_ (.A1(net38),
    .A2(net39),
    .A3(net40),
    .A4(_1939_),
    .B1(net57),
    .X(_2003_));
 sky130_fd_sc_hd__xor2_1 _2323_ (.A(net41),
    .B(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(_2004_),
    .A1(\m[18] ),
    .S(_1922_),
    .X(_2005_));
 sky130_fd_sc_hd__mux2_1 _2325_ (.A0(_2005_),
    .A1(\m[17] ),
    .S(_1925_),
    .X(_0357_));
 sky130_fd_sc_hd__or3_1 _2326_ (.A(_1807_),
    .B(net40),
    .C(_1941_),
    .X(_2006_));
 sky130_fd_sc_hd__o21ai_1 _2327_ (.A1(_1807_),
    .A2(_1941_),
    .B1(net40),
    .Y(_2007_));
 sky130_fd_sc_hd__and3_1 _2328_ (.A(_1923_),
    .B(_2006_),
    .C(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__o21ai_1 _2329_ (.A1(\m[17] ),
    .A2(_1923_),
    .B1(_0274_),
    .Y(_2009_));
 sky130_fd_sc_hd__a2bb2o_1 _2330_ (.A1_N(_2009_),
    .A2_N(_2008_),
    .B1(_1925_),
    .B2(\m[16] ),
    .X(_0356_));
 sky130_fd_sc_hd__o21ai_1 _2331_ (.A1(_1807_),
    .A2(_1940_),
    .B1(net39),
    .Y(_2010_));
 sky130_fd_sc_hd__o31a_1 _2332_ (.A1(_1807_),
    .A2(net39),
    .A3(_1940_),
    .B1(_1923_),
    .X(_2011_));
 sky130_fd_sc_hd__o2bb2a_1 _2333_ (.A1_N(_2011_),
    .A2_N(_2010_),
    .B1(_1923_),
    .B2(\m[16] ),
    .X(_2012_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(_2012_),
    .A1(\m[15] ),
    .S(_1925_),
    .X(_0355_));
 sky130_fd_sc_hd__a21oi_1 _2335_ (.A1(_1939_),
    .A2(net57),
    .B1(_1812_),
    .Y(_2013_));
 sky130_fd_sc_hd__a31o_1 _2336_ (.A1(_1939_),
    .A2(net57),
    .A3(_1812_),
    .B1(_1922_),
    .X(_2014_));
 sky130_fd_sc_hd__o221a_1 _2337_ (.A1(\m[15] ),
    .A2(_1923_),
    .B1(_2013_),
    .B2(_2014_),
    .C1(_0274_),
    .X(_2015_));
 sky130_fd_sc_hd__a21o_1 _2338_ (.A1(\m[14] ),
    .A2(_1925_),
    .B1(_2015_),
    .X(_0354_));
 sky130_fd_sc_hd__o21ai_1 _2339_ (.A1(net36),
    .A2(_1937_),
    .B1(net57),
    .Y(_2016_));
 sky130_fd_sc_hd__a21oi_1 _2340_ (.A1(_2016_),
    .A2(net37),
    .B1(_1922_),
    .Y(_2017_));
 sky130_fd_sc_hd__o21ai_1 _2341_ (.A1(net37),
    .A2(_2016_),
    .B1(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__o221a_1 _2342_ (.A1(\m[14] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__a21o_1 _2343_ (.A1(\m[13] ),
    .A2(_1925_),
    .B1(_2019_),
    .X(_0353_));
 sky130_fd_sc_hd__and3b_1 _2344_ (.A_N(net36),
    .B(_1937_),
    .C(net57),
    .X(_2020_));
 sky130_fd_sc_hd__a21boi_1 _2345_ (.A1(_1937_),
    .A2(net57),
    .B1_N(net36),
    .Y(_2021_));
 sky130_fd_sc_hd__or3_1 _2346_ (.A(_1922_),
    .B(_2020_),
    .C(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__o221a_1 _2347_ (.A1(\m[13] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__a21o_1 _2348_ (.A1(\m[12] ),
    .A2(_1925_),
    .B1(_2023_),
    .X(_0352_));
 sky130_fd_sc_hd__a21oi_1 _2349_ (.A1(_1936_),
    .A2(net57),
    .B1(_1811_),
    .Y(_2024_));
 sky130_fd_sc_hd__a31o_1 _2350_ (.A1(_1936_),
    .A2(net57),
    .A3(_1811_),
    .B1(_1922_),
    .X(_2025_));
 sky130_fd_sc_hd__o22a_1 _2351_ (.A1(\m[12] ),
    .A2(_1923_),
    .B1(_2024_),
    .B2(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__mux2_1 _2352_ (.A0(_2026_),
    .A1(\m[11] ),
    .S(_1925_),
    .X(_0351_));
 sky130_fd_sc_hd__o21ai_1 _2353_ (.A1(_1807_),
    .A2(_1934_),
    .B1(net34),
    .Y(_2027_));
 sky130_fd_sc_hd__or3_1 _2354_ (.A(_1807_),
    .B(net34),
    .C(_1934_),
    .X(_2028_));
 sky130_fd_sc_hd__and3_1 _2355_ (.A(_1923_),
    .B(_2027_),
    .C(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__o21ai_1 _2356_ (.A1(\m[11] ),
    .A2(_1923_),
    .B1(_0274_),
    .Y(_2030_));
 sky130_fd_sc_hd__a2bb2o_1 _2357_ (.A1_N(_2030_),
    .A2_N(_2029_),
    .B1(_1925_),
    .B2(\m[10] ),
    .X(_0350_));
 sky130_fd_sc_hd__a21o_1 _2358_ (.A1(_1931_),
    .A2(_1933_),
    .B1(_1807_),
    .X(_2031_));
 sky130_fd_sc_hd__a21oi_1 _2359_ (.A1(_2031_),
    .A2(net64),
    .B1(_1922_),
    .Y(_2032_));
 sky130_fd_sc_hd__o21ai_1 _2360_ (.A1(net64),
    .A2(_2031_),
    .B1(_2032_),
    .Y(_2033_));
 sky130_fd_sc_hd__o221a_1 _2361_ (.A1(\m[10] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__a21o_1 _2362_ (.A1(\m[9] ),
    .A2(_1925_),
    .B1(_2034_),
    .X(_0349_));
 sky130_fd_sc_hd__and3b_1 _2363_ (.A_N(net63),
    .B(_1932_),
    .C(net57),
    .X(_0404_));
 sky130_fd_sc_hd__a21boi_1 _2364_ (.A1(_1932_),
    .A2(net57),
    .B1_N(net63),
    .Y(_0405_));
 sky130_fd_sc_hd__or3_1 _2365_ (.A(_1922_),
    .B(_0404_),
    .C(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__o221a_1 _2366_ (.A1(\m[9] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__a21o_1 _2367_ (.A1(\m[8] ),
    .A2(_1925_),
    .B1(_0407_),
    .X(_0348_));
 sky130_fd_sc_hd__o21a_1 _2368_ (.A1(_1807_),
    .A2(_1931_),
    .B1(net62),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_1 _2369_ (.A(_1922_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__o31ai_1 _2370_ (.A1(_1807_),
    .A2(net62),
    .A3(_1931_),
    .B1(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__o221a_1 _2371_ (.A1(\m[8] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__a21o_1 _2372_ (.A1(\m[7] ),
    .A2(_1925_),
    .B1(_0411_),
    .X(_0347_));
 sky130_fd_sc_hd__o21ai_1 _2373_ (.A1(net60),
    .A2(_1928_),
    .B1(net57),
    .Y(_0412_));
 sky130_fd_sc_hd__a31o_1 _2374_ (.A1(_1929_),
    .A2(net57),
    .A3(_1810_),
    .B1(_1922_),
    .X(_0413_));
 sky130_fd_sc_hd__a21oi_1 _2375_ (.A1(net61),
    .A2(_0412_),
    .B1(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__o21ai_1 _2376_ (.A1(\m[7] ),
    .A2(_1923_),
    .B1(_0274_),
    .Y(_0415_));
 sky130_fd_sc_hd__a2bb2o_1 _2377_ (.A1_N(_0415_),
    .A2_N(_0414_),
    .B1(_1925_),
    .B2(\m[6] ),
    .X(_0346_));
 sky130_fd_sc_hd__a31o_1 _2378_ (.A1(_1926_),
    .A2(_1809_),
    .A3(_1808_),
    .B1(_1807_),
    .X(_0416_));
 sky130_fd_sc_hd__a21oi_1 _2379_ (.A1(_0416_),
    .A2(net60),
    .B1(_1922_),
    .Y(_0417_));
 sky130_fd_sc_hd__o21ai_1 _2380_ (.A1(net60),
    .A2(_0416_),
    .B1(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__o22a_1 _2381_ (.A1(\m[6] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _2382_ (.A1(\m[5] ),
    .A2(_1925_),
    .B1(_0418_),
    .B2(_0419_),
    .X(_0345_));
 sky130_fd_sc_hd__a21o_1 _2383_ (.A1(_1926_),
    .A2(_1808_),
    .B1(_1807_),
    .X(_0420_));
 sky130_fd_sc_hd__o21ai_1 _2384_ (.A1(net59),
    .A2(_0420_),
    .B1(_1923_),
    .Y(_0421_));
 sky130_fd_sc_hd__a21o_1 _2385_ (.A1(net59),
    .A2(_0420_),
    .B1(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__o221a_1 _2386_ (.A1(\m[5] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__a21o_1 _2387_ (.A1(\m[4] ),
    .A2(_1925_),
    .B1(_0423_),
    .X(_0344_));
 sky130_fd_sc_hd__o311a_1 _2388_ (.A1(net33),
    .A2(net44),
    .A3(net55),
    .B1(_1808_),
    .C1(net57),
    .X(_0424_));
 sky130_fd_sc_hd__o21a_1 _2389_ (.A1(_1807_),
    .A2(_1926_),
    .B1(net58),
    .X(_0425_));
 sky130_fd_sc_hd__or3_1 _2390_ (.A(_1922_),
    .B(_0424_),
    .C(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o221a_1 _2391_ (.A1(\m[4] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__a21o_1 _2392_ (.A1(\m[3] ),
    .A2(_1925_),
    .B1(_0427_),
    .X(_0343_));
 sky130_fd_sc_hd__o21ai_1 _2393_ (.A1(net33),
    .A2(net44),
    .B1(net57),
    .Y(_0428_));
 sky130_fd_sc_hd__a21oi_1 _2394_ (.A1(_0428_),
    .A2(net55),
    .B1(_1922_),
    .Y(_0429_));
 sky130_fd_sc_hd__o21ai_1 _2395_ (.A1(net55),
    .A2(_0428_),
    .B1(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__o22a_1 _2396_ (.A1(\m[3] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _2397_ (.A1(\m[2] ),
    .A2(_1925_),
    .B1(_0431_),
    .B2(_0430_),
    .X(_0342_));
 sky130_fd_sc_hd__and3_1 _2398_ (.A(net33),
    .B(net57),
    .C(net44),
    .X(_0432_));
 sky130_fd_sc_hd__a21oi_1 _2399_ (.A1(net33),
    .A2(net57),
    .B1(net44),
    .Y(_0433_));
 sky130_fd_sc_hd__o21ai_1 _2400_ (.A1(_0432_),
    .A2(_0433_),
    .B1(_1923_),
    .Y(_0434_));
 sky130_fd_sc_hd__o221a_1 _2401_ (.A1(\m[2] ),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_1817_),
    .C1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__a21o_1 _2402_ (.A1(\m[1] ),
    .A2(_1925_),
    .B1(_0435_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(net33),
    .A1(\m[1] ),
    .S(_1922_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(_0436_),
    .A1(\m[0] ),
    .S(_1925_),
    .X(_0340_));
 sky130_fd_sc_hd__o21ai_2 _2405_ (.A1(\m[0] ),
    .A2(_1923_),
    .B1(_0274_),
    .Y(_0437_));
 sky130_fd_sc_hd__and2_1 _2406_ (.A(net133),
    .B(\acc[63] ),
    .X(_0438_));
 sky130_fd_sc_hd__nand2b_1 _2407_ (.A_N(\q[8] ),
    .B(\count[0] ),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _2408_ (.A(\q[8] ),
    .B(net139),
    .Y(_0440_));
 sky130_fd_sc_hd__o211ai_1 _2409_ (.A1(net139),
    .A2(_1781_),
    .B1(net138),
    .C1(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2b_1 _2410_ (.A_N(\q[10] ),
    .B(\count[0] ),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _2411_ (.A(\q[10] ),
    .B(net139),
    .Y(_0443_));
 sky130_fd_sc_hd__o211ai_1 _2412_ (.A1(net139),
    .A2(_1779_),
    .B1(_1805_),
    .C1(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__o211ai_1 _2413_ (.A1(\q[11] ),
    .A2(\count[0] ),
    .B1(_0442_),
    .C1(_1805_),
    .Y(_0445_));
 sky130_fd_sc_hd__o211ai_1 _2414_ (.A1(\q[9] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0439_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand3_1 _2415_ (.A(_0445_),
    .B(_0446_),
    .C(net137),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2b_1 _2416_ (.A_N(\q[12] ),
    .B(\count[0] ),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _2417_ (.A(\q[12] ),
    .B(net139),
    .Y(_0449_));
 sky130_fd_sc_hd__o211ai_1 _2418_ (.A1(net139),
    .A2(_1777_),
    .B1(net138),
    .C1(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2b_1 _2419_ (.A_N(\q[14] ),
    .B(\count[0] ),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _2420_ (.A(\q[14] ),
    .B(net139),
    .Y(_0452_));
 sky130_fd_sc_hd__nand2b_1 _2421_ (.A_N(net139),
    .B(\q[15] ),
    .Y(_0453_));
 sky130_fd_sc_hd__o211ai_1 _2422_ (.A1(_1776_),
    .A2(_1806_),
    .B1(_0453_),
    .C1(_1805_),
    .Y(_0454_));
 sky130_fd_sc_hd__o211ai_1 _2423_ (.A1(\q[15] ),
    .A2(\count[0] ),
    .B1(_0451_),
    .C1(_1805_),
    .Y(_0455_));
 sky130_fd_sc_hd__o211ai_1 _2424_ (.A1(\q[13] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0448_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand3_1 _2425_ (.A(_1804_),
    .B(_0455_),
    .C(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__nand3_1 _2426_ (.A(_1804_),
    .B(_0450_),
    .C(_0454_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand3_1 _2427_ (.A(_0441_),
    .B(_0444_),
    .C(net137),
    .Y(_0459_));
 sky130_fd_sc_hd__nand3_2 _2428_ (.A(_1803_),
    .B(_0458_),
    .C(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nor2_1 _2429_ (.A(\q[7] ),
    .B(\count[0] ),
    .Y(_0461_));
 sky130_fd_sc_hd__and2b_1 _2430_ (.A_N(\q[6] ),
    .B(\count[0] ),
    .X(_0462_));
 sky130_fd_sc_hd__nand2b_1 _2431_ (.A_N(\q[6] ),
    .B(\count[0] ),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _2432_ (.A(\q[6] ),
    .B(net139),
    .Y(_0464_));
 sky130_fd_sc_hd__o211ai_2 _2433_ (.A1(net139),
    .A2(_1783_),
    .B1(_1805_),
    .C1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2b_1 _2434_ (.A_N(\q[4] ),
    .B(\count[0] ),
    .Y(_0466_));
 sky130_fd_sc_hd__nand2_1 _2435_ (.A(\q[4] ),
    .B(net139),
    .Y(_0467_));
 sky130_fd_sc_hd__o211ai_2 _2436_ (.A1(net139),
    .A2(_1784_),
    .B1(net138),
    .C1(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__o211ai_2 _2437_ (.A1(\q[5] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0466_),
    .Y(_0469_));
 sky130_fd_sc_hd__o311ai_4 _2438_ (.A1(\count[1] ),
    .A2(_0461_),
    .A3(_0462_),
    .B1(_0469_),
    .C1(_1804_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2b_1 _2439_ (.A_N(\q[2] ),
    .B(\count[0] ),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_1 _2440_ (.A(\q[2] ),
    .B(net139),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2b_1 _2441_ (.A_N(net139),
    .B(\q[3] ),
    .Y(_0473_));
 sky130_fd_sc_hd__o211ai_2 _2442_ (.A1(_1786_),
    .A2(_1806_),
    .B1(_0473_),
    .C1(_1805_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2b_4 _2443_ (.A_N(\q[0] ),
    .B(net139),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _2444_ (.A(\q[0] ),
    .B(net139),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_1 _2445_ (.A1(net139),
    .A2(_1787_),
    .B1(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__o21ai_1 _2446_ (.A1(\q[1] ),
    .A2(net139),
    .B1(_0475_),
    .Y(_0478_));
 sky130_fd_sc_hd__o211ai_1 _2447_ (.A1(net139),
    .A2(_1787_),
    .B1(net138),
    .C1(_0476_),
    .Y(_0479_));
 sky130_fd_sc_hd__o211ai_2 _2448_ (.A1(\q[1] ),
    .A2(net139),
    .B1(net138),
    .C1(_0475_),
    .Y(_0480_));
 sky130_fd_sc_hd__o211ai_2 _2449_ (.A1(\q[3] ),
    .A2(\count[0] ),
    .B1(_0471_),
    .C1(_1805_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand3_2 _2450_ (.A(_0481_),
    .B(net137),
    .C(_0480_),
    .Y(_0482_));
 sky130_fd_sc_hd__o211ai_1 _2451_ (.A1(_1805_),
    .A2(_0477_),
    .B1(_0474_),
    .C1(net137),
    .Y(_0483_));
 sky130_fd_sc_hd__nand3_1 _2452_ (.A(_1804_),
    .B(_0465_),
    .C(_0468_),
    .Y(_0484_));
 sky130_fd_sc_hd__nand2_1 _2453_ (.A(_0470_),
    .B(_0482_),
    .Y(_0485_));
 sky130_fd_sc_hd__nand3_2 _2454_ (.A(_0483_),
    .B(_0484_),
    .C(net136),
    .Y(_0486_));
 sky130_fd_sc_hd__nand3_2 _2455_ (.A(_1803_),
    .B(_0447_),
    .C(_0457_),
    .Y(_0487_));
 sky130_fd_sc_hd__o211ai_4 _2456_ (.A1(_1803_),
    .A2(_0485_),
    .B1(_0487_),
    .C1(\count[4] ),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _2457_ (.A(\q[17] ),
    .B(\count[0] ),
    .Y(_0489_));
 sky130_fd_sc_hd__and2b_1 _2458_ (.A_N(\q[16] ),
    .B(\count[0] ),
    .X(_0490_));
 sky130_fd_sc_hd__nand2b_1 _2459_ (.A_N(\q[16] ),
    .B(\count[0] ),
    .Y(_0491_));
 sky130_fd_sc_hd__nand2_1 _2460_ (.A(\q[16] ),
    .B(net139),
    .Y(_0492_));
 sky130_fd_sc_hd__o211ai_1 _2461_ (.A1(net139),
    .A2(_1774_),
    .B1(net138),
    .C1(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2b_1 _2462_ (.A_N(\q[18] ),
    .B(\count[0] ),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _2463_ (.A(\q[18] ),
    .B(net139),
    .Y(_0495_));
 sky130_fd_sc_hd__nand2b_1 _2464_ (.A_N(net139),
    .B(\q[19] ),
    .Y(_0496_));
 sky130_fd_sc_hd__o211ai_1 _2465_ (.A1(_1773_),
    .A2(_1806_),
    .B1(_0496_),
    .C1(_1805_),
    .Y(_0497_));
 sky130_fd_sc_hd__o211ai_1 _2466_ (.A1(\q[19] ),
    .A2(\count[0] ),
    .B1(_0494_),
    .C1(_1805_),
    .Y(_0498_));
 sky130_fd_sc_hd__o211ai_1 _2467_ (.A1(\q[17] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0491_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand3_1 _2468_ (.A(_0498_),
    .B(_0499_),
    .C(net137),
    .Y(_0500_));
 sky130_fd_sc_hd__nor2_1 _2469_ (.A(\q[21] ),
    .B(\count[0] ),
    .Y(_0501_));
 sky130_fd_sc_hd__and2b_1 _2470_ (.A_N(\q[20] ),
    .B(\count[0] ),
    .X(_0502_));
 sky130_fd_sc_hd__nand2b_1 _2471_ (.A_N(\q[20] ),
    .B(\count[0] ),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _2472_ (.A(\q[20] ),
    .B(net139),
    .Y(_0504_));
 sky130_fd_sc_hd__o211ai_1 _2473_ (.A1(net139),
    .A2(_1772_),
    .B1(net138),
    .C1(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__nand2b_1 _2474_ (.A_N(\q[22] ),
    .B(\count[0] ),
    .Y(_0506_));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(\q[22] ),
    .B(net139),
    .Y(_0507_));
 sky130_fd_sc_hd__o211ai_1 _2476_ (.A1(net139),
    .A2(_1770_),
    .B1(_1805_),
    .C1(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__o211ai_1 _2477_ (.A1(\q[23] ),
    .A2(\count[0] ),
    .B1(_0506_),
    .C1(_1805_),
    .Y(_0509_));
 sky130_fd_sc_hd__o211ai_1 _2478_ (.A1(\q[21] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0503_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand3_1 _2479_ (.A(_1804_),
    .B(_0509_),
    .C(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand3_1 _2480_ (.A(_1804_),
    .B(_0505_),
    .C(_0508_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand3_1 _2481_ (.A(_0497_),
    .B(net137),
    .C(_0493_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_2 _2482_ (.A(_0500_),
    .B(_0511_),
    .Y(_0514_));
 sky130_fd_sc_hd__nand3_1 _2483_ (.A(_0512_),
    .B(_0513_),
    .C(net136),
    .Y(_0515_));
 sky130_fd_sc_hd__nor2_2 _2484_ (.A(\q[25] ),
    .B(\count[0] ),
    .Y(_0516_));
 sky130_fd_sc_hd__and2b_1 _2485_ (.A_N(\q[24] ),
    .B(\count[0] ),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_1 _2486_ (.A(\q[24] ),
    .B(\count[0] ),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2b_1 _2487_ (.A_N(\count[0] ),
    .B(\q[25] ),
    .Y(_0519_));
 sky130_fd_sc_hd__nand3_1 _2488_ (.A(_0519_),
    .B(\count[1] ),
    .C(_0518_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2b_1 _2489_ (.A_N(\q[26] ),
    .B(\count[0] ),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _2490_ (.A(\q[26] ),
    .B(net139),
    .Y(_0522_));
 sky130_fd_sc_hd__o211ai_1 _2491_ (.A1(net139),
    .A2(_1767_),
    .B1(_1805_),
    .C1(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__o211ai_2 _2492_ (.A1(\q[27] ),
    .A2(\count[0] ),
    .B1(_0521_),
    .C1(_1805_),
    .Y(_0524_));
 sky130_fd_sc_hd__o311ai_4 _2493_ (.A1(_1805_),
    .A2(_0516_),
    .A3(_0517_),
    .B1(net137),
    .C1(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__nor2_2 _2494_ (.A(\q[29] ),
    .B(net140),
    .Y(_0526_));
 sky130_fd_sc_hd__and2b_2 _2495_ (.A_N(\q[28] ),
    .B(net140),
    .X(_0527_));
 sky130_fd_sc_hd__nand2_1 _2496_ (.A(\q[28] ),
    .B(net140),
    .Y(_0528_));
 sky130_fd_sc_hd__o211ai_1 _2497_ (.A1(net140),
    .A2(_1765_),
    .B1(\count[1] ),
    .C1(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2b_2 _2498_ (.A_N(\q[30] ),
    .B(net140),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _2499_ (.A(\q[30] ),
    .B(net140),
    .Y(_0531_));
 sky130_fd_sc_hd__o211ai_1 _2500_ (.A1(net140),
    .A2(_1764_),
    .B1(_1805_),
    .C1(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__o211ai_2 _2501_ (.A1(\q[31] ),
    .A2(net140),
    .B1(_0530_),
    .C1(_1805_),
    .Y(_0533_));
 sky130_fd_sc_hd__o311ai_4 _2502_ (.A1(_1805_),
    .A2(_0526_),
    .A3(_0527_),
    .B1(_0533_),
    .C1(_1804_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand3_1 _2503_ (.A(_1804_),
    .B(_0529_),
    .C(_0532_),
    .Y(_0535_));
 sky130_fd_sc_hd__nand3_1 _2504_ (.A(_0523_),
    .B(net137),
    .C(_0520_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand3_1 _2505_ (.A(_1803_),
    .B(_0535_),
    .C(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand3_1 _2506_ (.A(_1803_),
    .B(_0525_),
    .C(_0534_),
    .Y(_0538_));
 sky130_fd_sc_hd__o211ai_4 _2507_ (.A1(_1803_),
    .A2(_0514_),
    .B1(_0538_),
    .C1(_1802_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _2508_ (.A(_0488_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__and4b_1 _2509_ (.A_N(\acc[63] ),
    .B(_0488_),
    .C(_0539_),
    .D(net135),
    .X(_0541_));
 sky130_fd_sc_hd__o21a_1 _2510_ (.A1(_1801_),
    .A2(_0540_),
    .B1(\acc[63] ),
    .X(_0542_));
 sky130_fd_sc_hd__nor2_1 _2511_ (.A(_0541_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__nor2_8 _2512_ (.A(net135),
    .B(_1802_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_8 _2513_ (.A(_1801_),
    .B(\count[4] ),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _2514_ (.A(\count[1] ),
    .B(\count[0] ),
    .Y(_0546_));
 sky130_fd_sc_hd__nand3_4 _2515_ (.A(\q[31] ),
    .B(\count[1] ),
    .C(net140),
    .Y(_0547_));
 sky130_fd_sc_hd__and2_1 _2516_ (.A(net136),
    .B(\count[2] ),
    .X(_0548_));
 sky130_fd_sc_hd__and3_1 _2517_ (.A(\count[1] ),
    .B(\count[0] ),
    .C(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__and4_2 _2518_ (.A(\q[31] ),
    .B(\count[1] ),
    .C(net140),
    .D(_0548_),
    .X(_0550_));
 sky130_fd_sc_hd__nor2_1 _2519_ (.A(\q[18] ),
    .B(net139),
    .Y(_0551_));
 sky130_fd_sc_hd__and2b_1 _2520_ (.A_N(\q[17] ),
    .B(net139),
    .X(_0552_));
 sky130_fd_sc_hd__nand2b_1 _2521_ (.A_N(\q[17] ),
    .B(net139),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_1 _2522_ (.A(\q[17] ),
    .B(net139),
    .Y(_0554_));
 sky130_fd_sc_hd__o21ai_1 _2523_ (.A1(net139),
    .A2(_1773_),
    .B1(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand2b_1 _2524_ (.A_N(\q[15] ),
    .B(net139),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _2525_ (.A(\q[15] ),
    .B(net140),
    .Y(_0557_));
 sky130_fd_sc_hd__o211ai_1 _2526_ (.A1(net140),
    .A2(_1775_),
    .B1(net138),
    .C1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__o211ai_4 _2527_ (.A1(\q[16] ),
    .A2(net139),
    .B1(net138),
    .C1(_0556_),
    .Y(_0559_));
 sky130_fd_sc_hd__o311ai_4 _2528_ (.A1(net138),
    .A2(_0551_),
    .A3(_0552_),
    .B1(net137),
    .C1(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2b_1 _2529_ (.A_N(\q[19] ),
    .B(net139),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _2530_ (.A(\q[19] ),
    .B(net140),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2b_1 _2531_ (.A_N(net140),
    .B(\q[20] ),
    .Y(_0563_));
 sky130_fd_sc_hd__nand3_1 _2532_ (.A(_0563_),
    .B(net138),
    .C(_0562_),
    .Y(_0564_));
 sky130_fd_sc_hd__nor2_1 _2533_ (.A(\q[22] ),
    .B(net139),
    .Y(_0565_));
 sky130_fd_sc_hd__and2b_1 _2534_ (.A_N(\q[21] ),
    .B(net139),
    .X(_0566_));
 sky130_fd_sc_hd__nand2b_1 _2535_ (.A_N(\q[21] ),
    .B(net140),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _2536_ (.A(\q[21] ),
    .B(net140),
    .Y(_0568_));
 sky130_fd_sc_hd__o211ai_1 _2537_ (.A1(net140),
    .A2(_1771_),
    .B1(_1805_),
    .C1(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__o211ai_2 _2538_ (.A1(\q[20] ),
    .A2(net139),
    .B1(net138),
    .C1(_0561_),
    .Y(_0570_));
 sky130_fd_sc_hd__o31ai_1 _2539_ (.A1(net138),
    .A2(_0565_),
    .A3(_0566_),
    .B1(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__o311ai_4 _2540_ (.A1(net138),
    .A2(_0565_),
    .A3(_0566_),
    .B1(_0570_),
    .C1(_1804_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2b_1 _2541_ (.A_N(\q[23] ),
    .B(\count[0] ),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2b_1 _2542_ (.A_N(net140),
    .B(\q[24] ),
    .Y(_0574_));
 sky130_fd_sc_hd__o211ai_1 _2543_ (.A1(_1770_),
    .A2(_1806_),
    .B1(_0574_),
    .C1(net138),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2b_1 _2544_ (.A_N(\q[25] ),
    .B(net140),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _2545_ (.A(\q[25] ),
    .B(net140),
    .Y(_0577_));
 sky130_fd_sc_hd__o211ai_1 _2546_ (.A1(net140),
    .A2(_1768_),
    .B1(_1805_),
    .C1(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__o211ai_1 _2547_ (.A1(\q[26] ),
    .A2(net139),
    .B1(_0576_),
    .C1(_1805_),
    .Y(_0579_));
 sky130_fd_sc_hd__o211ai_1 _2548_ (.A1(\q[24] ),
    .A2(net140),
    .B1(net138),
    .C1(_0573_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand3_1 _2549_ (.A(_0579_),
    .B(_0580_),
    .C(net137),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _2550_ (.A(\q[29] ),
    .B(net140),
    .Y(_0582_));
 sky130_fd_sc_hd__nand2b_1 _2551_ (.A_N(net140),
    .B(\q[30] ),
    .Y(_0583_));
 sky130_fd_sc_hd__a21boi_1 _2552_ (.A1(_1806_),
    .A2(\q[30] ),
    .B1_N(_0582_),
    .Y(_0584_));
 sky130_fd_sc_hd__o211ai_1 _2553_ (.A1(_1765_),
    .A2(_1806_),
    .B1(_0583_),
    .C1(_1805_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2b_1 _2554_ (.A_N(\q[27] ),
    .B(net140),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _2555_ (.A(\q[27] ),
    .B(net140),
    .Y(_0587_));
 sky130_fd_sc_hd__o211ai_1 _2556_ (.A1(net140),
    .A2(_1766_),
    .B1(\count[1] ),
    .C1(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__o211ai_1 _2557_ (.A1(\q[28] ),
    .A2(net140),
    .B1(\count[1] ),
    .C1(_0586_),
    .Y(_0589_));
 sky130_fd_sc_hd__o211ai_2 _2558_ (.A1(\count[1] ),
    .A2(_0584_),
    .B1(_0589_),
    .C1(_1804_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand3_2 _2559_ (.A(_1803_),
    .B(_0581_),
    .C(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand3_2 _2560_ (.A(_0572_),
    .B(net136),
    .C(_0560_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand3_2 _2561_ (.A(_1802_),
    .B(_0591_),
    .C(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__and2b_2 _2562_ (.A_N(net139),
    .B(\q[0] ),
    .X(_0594_));
 sky130_fd_sc_hd__nand2b_2 _2563_ (.A_N(net139),
    .B(\q[0] ),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2b_1 _2564_ (.A_N(\q[1] ),
    .B(net139),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _2565_ (.A(\q[1] ),
    .B(net140),
    .Y(_0597_));
 sky130_fd_sc_hd__o211ai_4 _2566_ (.A1(net140),
    .A2(_1786_),
    .B1(_1805_),
    .C1(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__o211ai_2 _2567_ (.A1(\q[2] ),
    .A2(net139),
    .B1(_0596_),
    .C1(_1805_),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_1 _2568_ (.A1(_1805_),
    .A2(_0594_),
    .B1(_0598_),
    .Y(_0600_));
 sky130_fd_sc_hd__o211ai_4 _2569_ (.A1(_1805_),
    .A2(_0595_),
    .B1(net137),
    .C1(_0599_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2b_1 _2570_ (.A_N(\q[3] ),
    .B(net139),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _2571_ (.A(\q[3] ),
    .B(\count[0] ),
    .Y(_0603_));
 sky130_fd_sc_hd__o211ai_2 _2572_ (.A1(net140),
    .A2(_1785_),
    .B1(net138),
    .C1(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__nand2b_1 _2573_ (.A_N(\q[5] ),
    .B(net139),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_1 _2574_ (.A(\q[5] ),
    .B(net140),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2b_1 _2575_ (.A_N(net140),
    .B(\q[6] ),
    .Y(_0607_));
 sky130_fd_sc_hd__o211ai_2 _2576_ (.A1(_1784_),
    .A2(_1806_),
    .B1(_0607_),
    .C1(_1805_),
    .Y(_0608_));
 sky130_fd_sc_hd__o211ai_2 _2577_ (.A1(\q[6] ),
    .A2(net139),
    .B1(_0605_),
    .C1(_1805_),
    .Y(_0609_));
 sky130_fd_sc_hd__o211ai_2 _2578_ (.A1(\q[4] ),
    .A2(net139),
    .B1(net138),
    .C1(_0602_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand3_2 _2579_ (.A(_1804_),
    .B(_0609_),
    .C(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__nand3_2 _2580_ (.A(_1804_),
    .B(_0604_),
    .C(_0608_),
    .Y(_0612_));
 sky130_fd_sc_hd__o211ai_4 _2581_ (.A1(_1804_),
    .A2(_0600_),
    .B1(_0612_),
    .C1(net136),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2_1 _2582_ (.A(\q[8] ),
    .B(net139),
    .Y(_0614_));
 sky130_fd_sc_hd__and2b_1 _2583_ (.A_N(\q[7] ),
    .B(net139),
    .X(_0615_));
 sky130_fd_sc_hd__nand2b_1 _2584_ (.A_N(\q[7] ),
    .B(net139),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _2585_ (.A(\q[7] ),
    .B(net140),
    .Y(_0617_));
 sky130_fd_sc_hd__o211ai_1 _2586_ (.A1(net140),
    .A2(_1782_),
    .B1(net138),
    .C1(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2b_1 _2587_ (.A_N(\q[9] ),
    .B(net140),
    .Y(_0619_));
 sky130_fd_sc_hd__nand2_1 _2588_ (.A(\q[9] ),
    .B(net140),
    .Y(_0620_));
 sky130_fd_sc_hd__o211ai_1 _2589_ (.A1(net140),
    .A2(_1780_),
    .B1(_1805_),
    .C1(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__o211ai_1 _2590_ (.A1(\q[10] ),
    .A2(net139),
    .B1(_0619_),
    .C1(_1805_),
    .Y(_0622_));
 sky130_fd_sc_hd__o211ai_1 _2591_ (.A1(\q[8] ),
    .A2(net139),
    .B1(net138),
    .C1(_0616_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand3_1 _2592_ (.A(_0622_),
    .B(_0623_),
    .C(net137),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2b_1 _2593_ (.A_N(\q[11] ),
    .B(net139),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _2594_ (.A(\q[11] ),
    .B(net140),
    .Y(_0626_));
 sky130_fd_sc_hd__o211ai_1 _2595_ (.A1(net140),
    .A2(_1778_),
    .B1(net138),
    .C1(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2b_1 _2596_ (.A_N(\q[13] ),
    .B(net139),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _2597_ (.A(\q[13] ),
    .B(net140),
    .Y(_0629_));
 sky130_fd_sc_hd__o211ai_1 _2598_ (.A1(net140),
    .A2(_1776_),
    .B1(_1805_),
    .C1(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__o211ai_1 _2599_ (.A1(\q[14] ),
    .A2(net139),
    .B1(_0628_),
    .C1(_1805_),
    .Y(_0631_));
 sky130_fd_sc_hd__o211ai_2 _2600_ (.A1(\q[12] ),
    .A2(net139),
    .B1(net138),
    .C1(_0625_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand3_1 _2601_ (.A(_1804_),
    .B(_0631_),
    .C(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand3_1 _2602_ (.A(_1804_),
    .B(_0627_),
    .C(_0630_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand3_1 _2603_ (.A(_0618_),
    .B(_0621_),
    .C(net137),
    .Y(_0635_));
 sky130_fd_sc_hd__nand3_2 _2604_ (.A(_1803_),
    .B(_0634_),
    .C(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand3_1 _2605_ (.A(_1803_),
    .B(_0624_),
    .C(_0633_),
    .Y(_0637_));
 sky130_fd_sc_hd__nand3_1 _2606_ (.A(_0611_),
    .B(net136),
    .C(_0601_),
    .Y(_0638_));
 sky130_fd_sc_hd__nand3_4 _2607_ (.A(_0637_),
    .B(_0638_),
    .C(\count[4] ),
    .Y(_0639_));
 sky130_fd_sc_hd__a32oi_4 _2608_ (.A1(_0593_),
    .A2(_0639_),
    .A3(net135),
    .B1(_0544_),
    .B2(_0550_),
    .Y(_0640_));
 sky130_fd_sc_hd__a32o_1 _2609_ (.A1(_0593_),
    .A2(_0639_),
    .A3(net135),
    .B1(_0544_),
    .B2(_0550_),
    .X(_0641_));
 sky130_fd_sc_hd__and2_1 _2610_ (.A(_0641_),
    .B(\acc[62] ),
    .X(_0642_));
 sky130_fd_sc_hd__nand2_1 _2611_ (.A(_0641_),
    .B(\acc[62] ),
    .Y(_0643_));
 sky130_fd_sc_hd__nor2_1 _2612_ (.A(\count[4] ),
    .B(_1801_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_8 _2613_ (.A(_1802_),
    .B(net135),
    .Y(_0645_));
 sky130_fd_sc_hd__nand3_1 _2614_ (.A(_0460_),
    .B(_0486_),
    .C(_0644_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand3_1 _2615_ (.A(_0515_),
    .B(_0537_),
    .C(_0544_),
    .Y(_0647_));
 sky130_fd_sc_hd__nor2_8 _2616_ (.A(\count[5] ),
    .B(\count[4] ),
    .Y(_0648_));
 sky130_fd_sc_hd__or2_4 _2617_ (.A(net135),
    .B(\count[4] ),
    .X(_0649_));
 sky130_fd_sc_hd__a21bo_1 _2618_ (.A1(_0646_),
    .A2(_0647_),
    .B1_N(\acc[47] ),
    .X(_0650_));
 sky130_fd_sc_hd__o31a_1 _2619_ (.A1(_1803_),
    .A2(_1804_),
    .A3(_0547_),
    .B1(_0648_),
    .X(_0651_));
 sky130_fd_sc_hd__nand3_1 _2620_ (.A(_0591_),
    .B(_0592_),
    .C(_0544_),
    .Y(_0652_));
 sky130_fd_sc_hd__a31oi_2 _2621_ (.A1(_1802_),
    .A2(_0613_),
    .A3(_0636_),
    .B1(_1801_),
    .Y(_0653_));
 sky130_fd_sc_hd__a31o_1 _2622_ (.A1(_1802_),
    .A2(_0613_),
    .A3(_0636_),
    .B1(_1801_),
    .X(_0654_));
 sky130_fd_sc_hd__a31oi_2 _2623_ (.A1(_0591_),
    .A2(_0592_),
    .A3(_0544_),
    .B1(_0651_),
    .Y(_0655_));
 sky130_fd_sc_hd__o211ai_2 _2624_ (.A1(_0550_),
    .A2(_0649_),
    .B1(\acc[46] ),
    .C1(_0652_),
    .Y(_0656_));
 sky130_fd_sc_hd__and3_1 _2625_ (.A(_0654_),
    .B(_0655_),
    .C(\acc[46] ),
    .X(_0657_));
 sky130_fd_sc_hd__nand3b_2 _2626_ (.A_N(\acc[47] ),
    .B(_0646_),
    .C(_0647_),
    .Y(_0658_));
 sky130_fd_sc_hd__a21boi_1 _2627_ (.A1(_0657_),
    .A2(_0658_),
    .B1_N(_0650_),
    .Y(_0659_));
 sky130_fd_sc_hd__a21oi_1 _2628_ (.A1(_0654_),
    .A2(_0655_),
    .B1(\acc[46] ),
    .Y(_0660_));
 sky130_fd_sc_hd__a21o_1 _2629_ (.A1(_0654_),
    .A2(_0655_),
    .B1(\acc[46] ),
    .X(_0661_));
 sky130_fd_sc_hd__o21ai_1 _2630_ (.A1(_0653_),
    .A2(_0656_),
    .B1(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__o211ai_1 _2631_ (.A1(_0653_),
    .A2(_0656_),
    .B1(_0658_),
    .C1(_0650_),
    .Y(_0663_));
 sky130_fd_sc_hd__nor2_1 _2632_ (.A(_0660_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__o2111ai_1 _2633_ (.A1(_0653_),
    .A2(_0656_),
    .B1(_0658_),
    .C1(_0661_),
    .D1(_0650_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand3_1 _2634_ (.A(_0453_),
    .B(net138),
    .C(_0452_),
    .Y(_0666_));
 sky130_fd_sc_hd__o211ai_1 _2635_ (.A1(net139),
    .A2(_1774_),
    .B1(_1805_),
    .C1(_0492_),
    .Y(_0667_));
 sky130_fd_sc_hd__o211ai_2 _2636_ (.A1(\q[15] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0451_),
    .Y(_0668_));
 sky130_fd_sc_hd__o311ai_2 _2637_ (.A1(\count[1] ),
    .A2(_0489_),
    .A3(_0490_),
    .B1(net137),
    .C1(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__o211ai_1 _2638_ (.A1(net139),
    .A2(_1772_),
    .B1(_1805_),
    .C1(_0504_),
    .Y(_0670_));
 sky130_fd_sc_hd__nand3_1 _2639_ (.A(_0496_),
    .B(net138),
    .C(_0495_),
    .Y(_0671_));
 sky130_fd_sc_hd__o211ai_2 _2640_ (.A1(\q[19] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0494_),
    .Y(_0672_));
 sky130_fd_sc_hd__o31ai_1 _2641_ (.A1(\count[1] ),
    .A2(_0501_),
    .A3(_0502_),
    .B1(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__o311ai_2 _2642_ (.A1(\count[1] ),
    .A2(_0501_),
    .A3(_0502_),
    .B1(_0672_),
    .C1(_1804_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand3_1 _2643_ (.A(_1804_),
    .B(_0670_),
    .C(_0671_),
    .Y(_0675_));
 sky130_fd_sc_hd__nand3_1 _2644_ (.A(_0667_),
    .B(net137),
    .C(_0666_),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_1 _2645_ (.A(_0675_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand3_1 _2646_ (.A(_0675_),
    .B(_0676_),
    .C(net136),
    .Y(_0678_));
 sky130_fd_sc_hd__o211ai_1 _2647_ (.A1(net139),
    .A2(_1770_),
    .B1(\count[1] ),
    .C1(_0507_),
    .Y(_0679_));
 sky130_fd_sc_hd__o211ai_2 _2648_ (.A1(\count[0] ),
    .A2(_1769_),
    .B1(_1805_),
    .C1(_0518_),
    .Y(_0680_));
 sky130_fd_sc_hd__o211ai_2 _2649_ (.A1(\q[23] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0506_),
    .Y(_0681_));
 sky130_fd_sc_hd__o311ai_1 _2650_ (.A1(\count[1] ),
    .A2(_0516_),
    .A3(_0517_),
    .B1(net137),
    .C1(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__o211ai_1 _2651_ (.A1(net139),
    .A2(_1767_),
    .B1(\count[1] ),
    .C1(_0522_),
    .Y(_0683_));
 sky130_fd_sc_hd__o211ai_1 _2652_ (.A1(net140),
    .A2(_1765_),
    .B1(_1805_),
    .C1(_0528_),
    .Y(_0684_));
 sky130_fd_sc_hd__o211ai_2 _2653_ (.A1(\q[27] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0521_),
    .Y(_0685_));
 sky130_fd_sc_hd__o311ai_2 _2654_ (.A1(\count[1] ),
    .A2(_0526_),
    .A3(_0527_),
    .B1(_0685_),
    .C1(_1804_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand3_1 _2655_ (.A(_1804_),
    .B(_0683_),
    .C(_0684_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand3_1 _2656_ (.A(_0679_),
    .B(_0680_),
    .C(net137),
    .Y(_0688_));
 sky130_fd_sc_hd__nand3_1 _2657_ (.A(_1803_),
    .B(_0687_),
    .C(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand3_1 _2658_ (.A(_1803_),
    .B(_0682_),
    .C(_0686_),
    .Y(_0690_));
 sky130_fd_sc_hd__nand3_1 _2659_ (.A(_0674_),
    .B(\count[3] ),
    .C(_0669_),
    .Y(_0691_));
 sky130_fd_sc_hd__a21oi_1 _2660_ (.A1(_0678_),
    .A2(_0689_),
    .B1(_0545_),
    .Y(_0692_));
 sky130_fd_sc_hd__o211ai_1 _2661_ (.A1(net139),
    .A2(_1779_),
    .B1(net138),
    .C1(_0443_),
    .Y(_0693_));
 sky130_fd_sc_hd__o211ai_1 _2662_ (.A1(net139),
    .A2(_1777_),
    .B1(_1805_),
    .C1(_0449_),
    .Y(_0694_));
 sky130_fd_sc_hd__o211ai_1 _2663_ (.A1(\q[13] ),
    .A2(\count[0] ),
    .B1(_0448_),
    .C1(_1805_),
    .Y(_0695_));
 sky130_fd_sc_hd__o211ai_1 _2664_ (.A1(\q[11] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0442_),
    .Y(_0696_));
 sky130_fd_sc_hd__nand3_1 _2665_ (.A(_1804_),
    .B(_0695_),
    .C(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__o211ai_1 _2666_ (.A1(net139),
    .A2(_1783_),
    .B1(net138),
    .C1(_0464_),
    .Y(_0698_));
 sky130_fd_sc_hd__o211ai_1 _2667_ (.A1(net139),
    .A2(_1781_),
    .B1(_1805_),
    .C1(_0440_),
    .Y(_0699_));
 sky130_fd_sc_hd__o211ai_1 _2668_ (.A1(\q[9] ),
    .A2(\count[0] ),
    .B1(_0439_),
    .C1(_1805_),
    .Y(_0700_));
 sky130_fd_sc_hd__o211ai_1 _2669_ (.A1(\q[7] ),
    .A2(\count[0] ),
    .B1(\count[1] ),
    .C1(_0463_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand3_1 _2670_ (.A(_0700_),
    .B(_0701_),
    .C(net137),
    .Y(_0702_));
 sky130_fd_sc_hd__nand3_1 _2671_ (.A(_0698_),
    .B(_0699_),
    .C(net137),
    .Y(_0703_));
 sky130_fd_sc_hd__nand3_1 _2672_ (.A(_1804_),
    .B(_0693_),
    .C(_0694_),
    .Y(_0704_));
 sky130_fd_sc_hd__nand3_2 _2673_ (.A(_1803_),
    .B(_0703_),
    .C(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__nand3_1 _2674_ (.A(_0473_),
    .B(net138),
    .C(_0472_),
    .Y(_0706_));
 sky130_fd_sc_hd__o211ai_1 _2675_ (.A1(net139),
    .A2(_1784_),
    .B1(_1805_),
    .C1(_0467_),
    .Y(_0707_));
 sky130_fd_sc_hd__o211ai_2 _2676_ (.A1(\q[5] ),
    .A2(\count[0] ),
    .B1(_0466_),
    .C1(_1805_),
    .Y(_0708_));
 sky130_fd_sc_hd__o211ai_2 _2677_ (.A1(\q[3] ),
    .A2(\count[0] ),
    .B1(net138),
    .C1(_0471_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand3_4 _2678_ (.A(_1804_),
    .B(_0708_),
    .C(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o211a_1 _2679_ (.A1(\q[1] ),
    .A2(net139),
    .B1(_0475_),
    .C1(_1805_),
    .X(_0711_));
 sky130_fd_sc_hd__o21ai_1 _2680_ (.A1(net138),
    .A2(_0478_),
    .B1(net137),
    .Y(_0712_));
 sky130_fd_sc_hd__o2111ai_4 _2681_ (.A1(\q[1] ),
    .A2(net139),
    .B1(net137),
    .C1(_1805_),
    .D1(_0475_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand3_1 _2682_ (.A(_1804_),
    .B(_0706_),
    .C(_0707_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand3_2 _2683_ (.A(_0714_),
    .B(net136),
    .C(_0713_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand3_1 _2684_ (.A(_1803_),
    .B(_0697_),
    .C(_0702_),
    .Y(_0716_));
 sky130_fd_sc_hd__o211ai_1 _2685_ (.A1(_1804_),
    .A2(_0711_),
    .B1(\count[3] ),
    .C1(_0710_),
    .Y(_0717_));
 sky130_fd_sc_hd__o211a_1 _2686_ (.A1(\q[31] ),
    .A2(net140),
    .B1(\count[1] ),
    .C1(_0530_),
    .X(_0718_));
 sky130_fd_sc_hd__o211ai_2 _2687_ (.A1(\q[31] ),
    .A2(net140),
    .B1(\count[1] ),
    .C1(_0530_),
    .Y(_0719_));
 sky130_fd_sc_hd__o2111a_1 _2688_ (.A1(\q[31] ),
    .A2(net140),
    .B1(_0548_),
    .C1(\count[1] ),
    .D1(_0530_),
    .X(_0720_));
 sky130_fd_sc_hd__o21a_1 _2689_ (.A1(\count[4] ),
    .A2(_0720_),
    .B1(_1801_),
    .X(_0721_));
 sky130_fd_sc_hd__a31oi_1 _2690_ (.A1(_0705_),
    .A2(_0715_),
    .A3(_0644_),
    .B1(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__a31o_1 _2691_ (.A1(_0705_),
    .A2(_0715_),
    .A3(_0644_),
    .B1(_0721_),
    .X(_0723_));
 sky130_fd_sc_hd__nand3b_1 _2692_ (.A_N(_0692_),
    .B(_0723_),
    .C(\acc[45] ),
    .Y(_0724_));
 sky130_fd_sc_hd__o21bai_2 _2693_ (.A1(_0692_),
    .A2(_0722_),
    .B1_N(\acc[45] ),
    .Y(_0725_));
 sky130_fd_sc_hd__a21oi_1 _2694_ (.A1(\q[31] ),
    .A2(net140),
    .B1(\count[1] ),
    .Y(_0726_));
 sky130_fd_sc_hd__a31o_2 _2695_ (.A1(_0583_),
    .A2(\count[1] ),
    .A3(_0582_),
    .B1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__a21oi_1 _2696_ (.A1(_0584_),
    .A2(\count[1] ),
    .B1(_0726_),
    .Y(_0728_));
 sky130_fd_sc_hd__nor2_1 _2697_ (.A(_1804_),
    .B(_0727_),
    .Y(_0729_));
 sky130_fd_sc_hd__o311a_1 _2698_ (.A1(_1803_),
    .A2(_1804_),
    .A3(_0727_),
    .B1(_1802_),
    .C1(_1801_),
    .X(_0730_));
 sky130_fd_sc_hd__a31o_1 _2699_ (.A1(_0728_),
    .A2(\count[2] ),
    .A3(net136),
    .B1(_0649_),
    .X(_0731_));
 sky130_fd_sc_hd__o211ai_1 _2700_ (.A1(net140),
    .A2(_1776_),
    .B1(net138),
    .C1(_0629_),
    .Y(_0732_));
 sky130_fd_sc_hd__o211ai_1 _2701_ (.A1(net140),
    .A2(_1775_),
    .B1(_1805_),
    .C1(_0557_),
    .Y(_0733_));
 sky130_fd_sc_hd__o211ai_1 _2702_ (.A1(\q[16] ),
    .A2(net139),
    .B1(_0556_),
    .C1(_1805_),
    .Y(_0734_));
 sky130_fd_sc_hd__o211ai_1 _2703_ (.A1(\q[14] ),
    .A2(net139),
    .B1(net138),
    .C1(_0628_),
    .Y(_0735_));
 sky130_fd_sc_hd__nand3_1 _2704_ (.A(_0734_),
    .B(_0735_),
    .C(net137),
    .Y(_0736_));
 sky130_fd_sc_hd__nand3_1 _2705_ (.A(_1805_),
    .B(_0562_),
    .C(_0563_),
    .Y(_0737_));
 sky130_fd_sc_hd__o211ai_1 _2706_ (.A1(\q[20] ),
    .A2(net139),
    .B1(_0561_),
    .C1(_1805_),
    .Y(_0738_));
 sky130_fd_sc_hd__o211ai_1 _2707_ (.A1(\q[18] ),
    .A2(net139),
    .B1(net138),
    .C1(_0553_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand3_1 _2708_ (.A(_1804_),
    .B(_0738_),
    .C(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__o211ai_1 _2709_ (.A1(_1805_),
    .A2(_0555_),
    .B1(_0737_),
    .C1(_1804_),
    .Y(_0741_));
 sky130_fd_sc_hd__nand3_1 _2710_ (.A(_0732_),
    .B(_0733_),
    .C(net137),
    .Y(_0742_));
 sky130_fd_sc_hd__o21ai_1 _2711_ (.A1(_0565_),
    .A2(_0566_),
    .B1(net138),
    .Y(_0743_));
 sky130_fd_sc_hd__o211ai_1 _2712_ (.A1(_1770_),
    .A2(_1806_),
    .B1(_0574_),
    .C1(_1805_),
    .Y(_0744_));
 sky130_fd_sc_hd__o211ai_1 _2713_ (.A1(\q[24] ),
    .A2(net140),
    .B1(_0573_),
    .C1(_1805_),
    .Y(_0745_));
 sky130_fd_sc_hd__o211ai_1 _2714_ (.A1(\q[22] ),
    .A2(net140),
    .B1(net138),
    .C1(_0567_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand3_1 _2715_ (.A(_0745_),
    .B(_0746_),
    .C(net137),
    .Y(_0747_));
 sky130_fd_sc_hd__o211ai_2 _2716_ (.A1(net140),
    .A2(_1768_),
    .B1(net138),
    .C1(_0577_),
    .Y(_0748_));
 sky130_fd_sc_hd__o211ai_2 _2717_ (.A1(net140),
    .A2(_1766_),
    .B1(_1805_),
    .C1(_0587_),
    .Y(_0749_));
 sky130_fd_sc_hd__o211ai_1 _2718_ (.A1(\q[28] ),
    .A2(net140),
    .B1(_0586_),
    .C1(_1805_),
    .Y(_0750_));
 sky130_fd_sc_hd__o211ai_1 _2719_ (.A1(\q[26] ),
    .A2(net139),
    .B1(net138),
    .C1(_0576_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand3_1 _2720_ (.A(_1804_),
    .B(_0750_),
    .C(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand3_1 _2721_ (.A(_1804_),
    .B(_0748_),
    .C(_0749_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand3_1 _2722_ (.A(_0743_),
    .B(_0744_),
    .C(net137),
    .Y(_0754_));
 sky130_fd_sc_hd__nand3_2 _2723_ (.A(_1803_),
    .B(_0747_),
    .C(_0752_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand3_2 _2724_ (.A(_0740_),
    .B(\count[3] ),
    .C(_0736_),
    .Y(_0756_));
 sky130_fd_sc_hd__nand2_2 _2725_ (.A(_0755_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__a31o_1 _2726_ (.A1(_1805_),
    .A2(_1806_),
    .A3(\q[0] ),
    .B1(_1804_),
    .X(_0758_));
 sky130_fd_sc_hd__o211ai_2 _2727_ (.A1(net140),
    .A2(_1786_),
    .B1(net138),
    .C1(_0597_),
    .Y(_0759_));
 sky130_fd_sc_hd__o211ai_2 _2728_ (.A1(net140),
    .A2(_1785_),
    .B1(_1805_),
    .C1(_0603_),
    .Y(_0760_));
 sky130_fd_sc_hd__o211ai_2 _2729_ (.A1(\q[4] ),
    .A2(net139),
    .B1(_0602_),
    .C1(_1805_),
    .Y(_0761_));
 sky130_fd_sc_hd__o211ai_2 _2730_ (.A1(\q[2] ),
    .A2(net139),
    .B1(net138),
    .C1(_0596_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand3_2 _2731_ (.A(_1804_),
    .B(_0761_),
    .C(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand3_2 _2732_ (.A(_1804_),
    .B(_0759_),
    .C(_0760_),
    .Y(_0764_));
 sky130_fd_sc_hd__nand4_4 _2733_ (.A(_1805_),
    .B(_1806_),
    .C(\q[0] ),
    .D(net137),
    .Y(_0765_));
 sky130_fd_sc_hd__nand3_2 _2734_ (.A(_0764_),
    .B(_0765_),
    .C(net136),
    .Y(_0766_));
 sky130_fd_sc_hd__o211ai_1 _2735_ (.A1(net140),
    .A2(_1780_),
    .B1(net138),
    .C1(_0620_),
    .Y(_0767_));
 sky130_fd_sc_hd__o211ai_1 _2736_ (.A1(net140),
    .A2(_1778_),
    .B1(_1805_),
    .C1(_0626_),
    .Y(_0768_));
 sky130_fd_sc_hd__o211ai_1 _2737_ (.A1(\q[12] ),
    .A2(net139),
    .B1(_0625_),
    .C1(_1805_),
    .Y(_0769_));
 sky130_fd_sc_hd__o211ai_1 _2738_ (.A1(\q[10] ),
    .A2(net139),
    .B1(net138),
    .C1(_0619_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand3_1 _2739_ (.A(_1804_),
    .B(_0769_),
    .C(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__o211ai_1 _2740_ (.A1(net140),
    .A2(_1782_),
    .B1(_1805_),
    .C1(_0617_),
    .Y(_0772_));
 sky130_fd_sc_hd__nand3_1 _2741_ (.A(_0607_),
    .B(net138),
    .C(_0606_),
    .Y(_0773_));
 sky130_fd_sc_hd__o211ai_2 _2742_ (.A1(\q[6] ),
    .A2(net139),
    .B1(net138),
    .C1(_0605_),
    .Y(_0774_));
 sky130_fd_sc_hd__o311ai_2 _2743_ (.A1(net138),
    .A2(_0614_),
    .A3(_0615_),
    .B1(net137),
    .C1(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand3_1 _2744_ (.A(_0772_),
    .B(_0773_),
    .C(net137),
    .Y(_0776_));
 sky130_fd_sc_hd__nand3_1 _2745_ (.A(_1804_),
    .B(_0767_),
    .C(_0768_),
    .Y(_0777_));
 sky130_fd_sc_hd__nand3_2 _2746_ (.A(_1803_),
    .B(_0776_),
    .C(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand3_1 _2747_ (.A(_0763_),
    .B(\count[3] ),
    .C(_0758_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand3_1 _2748_ (.A(_1803_),
    .B(_0771_),
    .C(_0775_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand3_1 _2749_ (.A(_1802_),
    .B(_0766_),
    .C(_0778_),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_1 _2750_ (.A(_0781_),
    .B(net135),
    .Y(_0782_));
 sky130_fd_sc_hd__a31oi_1 _2751_ (.A1(_0544_),
    .A2(_0755_),
    .A3(_0756_),
    .B1(_0730_),
    .Y(_0783_));
 sky130_fd_sc_hd__o2111a_1 _2752_ (.A1(_0757_),
    .A2(_0545_),
    .B1(\acc[44] ),
    .C1(_0731_),
    .D1(_0782_),
    .X(_0784_));
 sky130_fd_sc_hd__o2111ai_2 _2753_ (.A1(_0757_),
    .A2(_0545_),
    .B1(\acc[44] ),
    .C1(_0731_),
    .D1(_0782_),
    .Y(_0785_));
 sky130_fd_sc_hd__a21bo_1 _2754_ (.A1(_0724_),
    .A2(_0785_),
    .B1_N(_0725_),
    .X(_0786_));
 sky130_fd_sc_hd__and3_2 _2755_ (.A(_0529_),
    .B(_0532_),
    .C(\count[2] ),
    .X(_0787_));
 sky130_fd_sc_hd__a21oi_2 _2756_ (.A1(net136),
    .A2(_0787_),
    .B1(_0649_),
    .Y(_0788_));
 sky130_fd_sc_hd__nand3_1 _2757_ (.A(_0455_),
    .B(_0456_),
    .C(net137),
    .Y(_0789_));
 sky130_fd_sc_hd__nand3_1 _2758_ (.A(_1804_),
    .B(_0498_),
    .C(_0499_),
    .Y(_0790_));
 sky130_fd_sc_hd__nand3_1 _2759_ (.A(_1804_),
    .B(_0493_),
    .C(_0497_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand3_1 _2760_ (.A(_0454_),
    .B(net137),
    .C(_0450_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_1 _2761_ (.A(_0791_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__nand3_1 _2762_ (.A(_0791_),
    .B(_0792_),
    .C(net136),
    .Y(_0794_));
 sky130_fd_sc_hd__nand3_1 _2763_ (.A(_1804_),
    .B(_0520_),
    .C(_0523_),
    .Y(_0795_));
 sky130_fd_sc_hd__nand3_1 _2764_ (.A(_0505_),
    .B(_0508_),
    .C(net137),
    .Y(_0796_));
 sky130_fd_sc_hd__nand3_2 _2765_ (.A(_1803_),
    .B(_0795_),
    .C(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__o21a_1 _2766_ (.A1(_1803_),
    .A2(_0793_),
    .B1(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__o311ai_1 _2767_ (.A1(\count[1] ),
    .A2(_0461_),
    .A3(_0462_),
    .B1(net137),
    .C1(_0469_),
    .Y(_0799_));
 sky130_fd_sc_hd__nand3_1 _2768_ (.A(_1804_),
    .B(_0445_),
    .C(_0446_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand3_1 _2769_ (.A(_1804_),
    .B(_0441_),
    .C(_0444_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand3_2 _2770_ (.A(_0465_),
    .B(_0468_),
    .C(net137),
    .Y(_0802_));
 sky130_fd_sc_hd__nand3_4 _2771_ (.A(_1803_),
    .B(_0801_),
    .C(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__a31o_2 _2772_ (.A1(_1804_),
    .A2(_0474_),
    .A3(_0479_),
    .B1(_1803_),
    .X(_0804_));
 sky130_fd_sc_hd__a21oi_2 _2773_ (.A1(_0794_),
    .A2(_0797_),
    .B1(_0545_),
    .Y(_0805_));
 sky130_fd_sc_hd__nand3_1 _2774_ (.A(_1802_),
    .B(_0803_),
    .C(_0804_),
    .Y(_0806_));
 sky130_fd_sc_hd__a31oi_1 _2775_ (.A1(_1802_),
    .A2(_0803_),
    .A3(_0804_),
    .B1(_1801_),
    .Y(_0807_));
 sky130_fd_sc_hd__a2111oi_1 _2776_ (.A1(_0806_),
    .A2(net135),
    .B1(_1788_),
    .C1(_0788_),
    .D1(_0805_),
    .Y(_0808_));
 sky130_fd_sc_hd__a2111o_2 _2777_ (.A1(_0806_),
    .A2(net135),
    .B1(_1788_),
    .C1(_0788_),
    .D1(_0805_),
    .X(_0809_));
 sky130_fd_sc_hd__o31a_1 _2778_ (.A1(_0788_),
    .A2(_0805_),
    .A3(_0807_),
    .B1(_1788_),
    .X(_0810_));
 sky130_fd_sc_hd__o31ai_1 _2779_ (.A1(_0788_),
    .A2(_0805_),
    .A3(_0807_),
    .B1(_1788_),
    .Y(_0811_));
 sky130_fd_sc_hd__nor2_1 _2780_ (.A(_0808_),
    .B(_0810_),
    .Y(_0812_));
 sky130_fd_sc_hd__nand2_1 _2781_ (.A(_0809_),
    .B(_0811_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand3_1 _2782_ (.A(_0631_),
    .B(_0632_),
    .C(net137),
    .Y(_0814_));
 sky130_fd_sc_hd__o311ai_2 _2783_ (.A1(net138),
    .A2(_0551_),
    .A3(_0552_),
    .B1(_0559_),
    .C1(_1804_),
    .Y(_0815_));
 sky130_fd_sc_hd__o211ai_1 _2784_ (.A1(net138),
    .A2(_0555_),
    .B1(_0558_),
    .C1(_1804_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand3_1 _2785_ (.A(_0627_),
    .B(_0630_),
    .C(net137),
    .Y(_0817_));
 sky130_fd_sc_hd__nand3_1 _2786_ (.A(_1804_),
    .B(_0579_),
    .C(_0580_),
    .Y(_0818_));
 sky130_fd_sc_hd__nand3_1 _2787_ (.A(_0569_),
    .B(net137),
    .C(_0564_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand3_1 _2788_ (.A(_1804_),
    .B(_0575_),
    .C(_0578_),
    .Y(_0820_));
 sky130_fd_sc_hd__o211ai_2 _2789_ (.A1(_1804_),
    .A2(_0571_),
    .B1(_0818_),
    .C1(_1803_),
    .Y(_0821_));
 sky130_fd_sc_hd__nand3_2 _2790_ (.A(_0815_),
    .B(net136),
    .C(_0814_),
    .Y(_0822_));
 sky130_fd_sc_hd__nand2_2 _2791_ (.A(_0821_),
    .B(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__nand4_1 _2792_ (.A(_1801_),
    .B(_0821_),
    .C(_0822_),
    .D(\count[4] ),
    .Y(_0824_));
 sky130_fd_sc_hd__nand3_1 _2793_ (.A(_0609_),
    .B(_0610_),
    .C(net137),
    .Y(_0825_));
 sky130_fd_sc_hd__nand3_1 _2794_ (.A(_1804_),
    .B(_0622_),
    .C(_0623_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand3_1 _2795_ (.A(_1804_),
    .B(_0618_),
    .C(_0621_),
    .Y(_0827_));
 sky130_fd_sc_hd__nand3_1 _2796_ (.A(_0608_),
    .B(net137),
    .C(_0604_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand3_2 _2797_ (.A(_1803_),
    .B(_0827_),
    .C(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__a21oi_2 _2798_ (.A1(_0595_),
    .A2(net138),
    .B1(net137),
    .Y(_0830_));
 sky130_fd_sc_hd__o211ai_4 _2799_ (.A1(_0594_),
    .A2(_1805_),
    .B1(_1804_),
    .C1(_0598_),
    .Y(_0831_));
 sky130_fd_sc_hd__a21o_1 _2800_ (.A1(_0830_),
    .A2(_0598_),
    .B1(_1803_),
    .X(_0832_));
 sky130_fd_sc_hd__nand3_1 _2801_ (.A(_1803_),
    .B(_0825_),
    .C(_0826_),
    .Y(_0833_));
 sky130_fd_sc_hd__nand3_1 _2802_ (.A(_0585_),
    .B(_0588_),
    .C(\count[2] ),
    .Y(_0834_));
 sky130_fd_sc_hd__and3_1 _2803_ (.A(_1804_),
    .B(\count[1] ),
    .C(net140),
    .X(_0835_));
 sky130_fd_sc_hd__a32o_1 _2804_ (.A1(_0585_),
    .A2(_0588_),
    .A3(\count[2] ),
    .B1(_0835_),
    .B2(\q[31] ),
    .X(_0836_));
 sky130_fd_sc_hd__a21oi_1 _2805_ (.A1(_0831_),
    .A2(net136),
    .B1(\count[4] ),
    .Y(_0837_));
 sky130_fd_sc_hd__a21o_1 _2806_ (.A1(_0837_),
    .A2(_0829_),
    .B1(_1801_),
    .X(_0838_));
 sky130_fd_sc_hd__a21o_1 _2807_ (.A1(_0836_),
    .A2(net136),
    .B1(_0649_),
    .X(_0839_));
 sky130_fd_sc_hd__a31oi_1 _2808_ (.A1(_0824_),
    .A2(_0838_),
    .A3(_0839_),
    .B1(\acc[42] ),
    .Y(_0840_));
 sky130_fd_sc_hd__a31o_1 _2809_ (.A1(_0824_),
    .A2(_0838_),
    .A3(_0839_),
    .B1(\acc[42] ),
    .X(_0841_));
 sky130_fd_sc_hd__and4_1 _2810_ (.A(_0824_),
    .B(_0838_),
    .C(_0839_),
    .D(\acc[42] ),
    .X(_0842_));
 sky130_fd_sc_hd__o2111ai_4 _2811_ (.A1(_0545_),
    .A2(_0823_),
    .B1(_0839_),
    .C1(\acc[42] ),
    .D1(_0838_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _2812_ (.A(_0840_),
    .B(_0842_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _2813_ (.A(_0841_),
    .B(_0843_),
    .Y(_0845_));
 sky130_fd_sc_hd__and4_1 _2814_ (.A(_0809_),
    .B(_0811_),
    .C(_0841_),
    .D(_0843_),
    .X(_0846_));
 sky130_fd_sc_hd__nand4_1 _2815_ (.A(_0809_),
    .B(_0811_),
    .C(_0841_),
    .D(_0843_),
    .Y(_0847_));
 sky130_fd_sc_hd__nand3_1 _2816_ (.A(_0695_),
    .B(_0696_),
    .C(net137),
    .Y(_0848_));
 sky130_fd_sc_hd__o311ai_2 _2817_ (.A1(\count[1] ),
    .A2(_0489_),
    .A3(_0490_),
    .B1(_0668_),
    .C1(_1804_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand3_1 _2818_ (.A(_1804_),
    .B(_0666_),
    .C(_0667_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand3_1 _2819_ (.A(_0693_),
    .B(_0694_),
    .C(net137),
    .Y(_0851_));
 sky130_fd_sc_hd__o311ai_2 _2820_ (.A1(\count[1] ),
    .A2(_0516_),
    .A3(_0517_),
    .B1(_0681_),
    .C1(_1804_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand3_1 _2821_ (.A(_1804_),
    .B(_0679_),
    .C(_0680_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand3_1 _2822_ (.A(_0670_),
    .B(_0671_),
    .C(net137),
    .Y(_0854_));
 sky130_fd_sc_hd__o211ai_2 _2823_ (.A1(_1804_),
    .A2(_0673_),
    .B1(_0852_),
    .C1(_1803_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand3_2 _2824_ (.A(_0849_),
    .B(\count[3] ),
    .C(_0848_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand3_1 _2825_ (.A(_0855_),
    .B(_0856_),
    .C(_0544_),
    .Y(_0857_));
 sky130_fd_sc_hd__nand3_1 _2826_ (.A(_0708_),
    .B(_0709_),
    .C(net137),
    .Y(_0858_));
 sky130_fd_sc_hd__nand3_1 _2827_ (.A(_1804_),
    .B(_0700_),
    .C(_0701_),
    .Y(_0859_));
 sky130_fd_sc_hd__nand3_1 _2828_ (.A(_1804_),
    .B(_0698_),
    .C(_0699_),
    .Y(_0860_));
 sky130_fd_sc_hd__nand3_1 _2829_ (.A(_0707_),
    .B(net137),
    .C(_0706_),
    .Y(_0861_));
 sky130_fd_sc_hd__nand3_2 _2830_ (.A(_1803_),
    .B(_0860_),
    .C(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__o21ba_1 _2831_ (.A1(\q[1] ),
    .A2(net139),
    .B1_N(net137),
    .X(_0863_));
 sky130_fd_sc_hd__o2111ai_1 _2832_ (.A1(\q[1] ),
    .A2(net139),
    .B1(_0475_),
    .C1(_1804_),
    .D1(_1805_),
    .Y(_0864_));
 sky130_fd_sc_hd__a31o_1 _2833_ (.A1(_0863_),
    .A2(_0475_),
    .A3(_1805_),
    .B1(_1803_),
    .X(_0865_));
 sky130_fd_sc_hd__o311ai_2 _2834_ (.A1(\count[1] ),
    .A2(_0526_),
    .A3(_0527_),
    .B1(\count[2] ),
    .C1(_0685_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand3_1 _2835_ (.A(_0683_),
    .B(_0684_),
    .C(\count[2] ),
    .Y(_0867_));
 sky130_fd_sc_hd__o21ai_1 _2836_ (.A1(\count[2] ),
    .A2(_0718_),
    .B1(_0866_),
    .Y(_0868_));
 sky130_fd_sc_hd__o211a_1 _2837_ (.A1(\count[2] ),
    .A2(_0718_),
    .B1(net136),
    .C1(_0866_),
    .X(_0869_));
 sky130_fd_sc_hd__a21oi_1 _2838_ (.A1(_0864_),
    .A2(net136),
    .B1(\count[4] ),
    .Y(_0870_));
 sky130_fd_sc_hd__a21o_1 _2839_ (.A1(_0862_),
    .A2(_0870_),
    .B1(_1801_),
    .X(_0871_));
 sky130_fd_sc_hd__o21ai_1 _2840_ (.A1(_1803_),
    .A2(_0868_),
    .B1(_0648_),
    .Y(_0872_));
 sky130_fd_sc_hd__and4_1 _2841_ (.A(_0871_),
    .B(\acc[41] ),
    .C(_0857_),
    .D(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__o2111ai_1 _2842_ (.A1(_0869_),
    .A2(_0649_),
    .B1(\acc[41] ),
    .C1(_0857_),
    .D1(_0871_),
    .Y(_0874_));
 sky130_fd_sc_hd__a31oi_2 _2843_ (.A1(_0857_),
    .A2(_0871_),
    .A3(_0872_),
    .B1(\acc[41] ),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _2844_ (.A(_0727_),
    .B(_1804_),
    .Y(_0876_));
 sky130_fd_sc_hd__a21o_1 _2845_ (.A1(_0748_),
    .A2(_0749_),
    .B1(_1804_),
    .X(_0877_));
 sky130_fd_sc_hd__nand3_1 _2846_ (.A(_0748_),
    .B(_0749_),
    .C(\count[2] ),
    .Y(_0878_));
 sky130_fd_sc_hd__a31o_1 _2847_ (.A1(_0876_),
    .A2(_0877_),
    .A3(net136),
    .B1(_0649_),
    .X(_0879_));
 sky130_fd_sc_hd__nand3_1 _2848_ (.A(_0769_),
    .B(_0770_),
    .C(net137),
    .Y(_0880_));
 sky130_fd_sc_hd__nand3_1 _2849_ (.A(_1804_),
    .B(_0734_),
    .C(_0735_),
    .Y(_0881_));
 sky130_fd_sc_hd__nand3_1 _2850_ (.A(_1804_),
    .B(_0732_),
    .C(_0733_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand3_1 _2851_ (.A(_0767_),
    .B(_0768_),
    .C(net137),
    .Y(_0883_));
 sky130_fd_sc_hd__nand3_1 _2852_ (.A(_0738_),
    .B(_0739_),
    .C(net137),
    .Y(_0884_));
 sky130_fd_sc_hd__nand3_1 _2853_ (.A(_1804_),
    .B(_0745_),
    .C(_0746_),
    .Y(_0885_));
 sky130_fd_sc_hd__nand3_1 _2854_ (.A(_1804_),
    .B(_0743_),
    .C(_0744_),
    .Y(_0886_));
 sky130_fd_sc_hd__o211ai_1 _2855_ (.A1(_1805_),
    .A2(_0555_),
    .B1(_0737_),
    .C1(net137),
    .Y(_0887_));
 sky130_fd_sc_hd__nand3_2 _2856_ (.A(_1803_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0888_));
 sky130_fd_sc_hd__nand3_2 _2857_ (.A(_0881_),
    .B(\count[3] ),
    .C(_0880_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand2_2 _2858_ (.A(_0888_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__o311ai_1 _2859_ (.A1(net138),
    .A2(_0614_),
    .A3(_0615_),
    .B1(_0774_),
    .C1(_1804_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand3_1 _2860_ (.A(_0761_),
    .B(_0762_),
    .C(net137),
    .Y(_0892_));
 sky130_fd_sc_hd__nand3_2 _2861_ (.A(_0759_),
    .B(_0760_),
    .C(net137),
    .Y(_0893_));
 sky130_fd_sc_hd__nand3_1 _2862_ (.A(_1804_),
    .B(_0772_),
    .C(_0773_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand3_4 _2863_ (.A(_1803_),
    .B(_0893_),
    .C(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__nor2_1 _2864_ (.A(net137),
    .B(net138),
    .Y(_0896_));
 sky130_fd_sc_hd__and3_1 _2865_ (.A(\q[0] ),
    .B(_0896_),
    .C(_1806_),
    .X(_0897_));
 sky130_fd_sc_hd__a31o_2 _2866_ (.A1(\q[0] ),
    .A2(_0896_),
    .A3(_1806_),
    .B1(_1803_),
    .X(_0898_));
 sky130_fd_sc_hd__a31oi_4 _2867_ (.A1(_1802_),
    .A2(_0895_),
    .A3(_0898_),
    .B1(_1801_),
    .Y(_0899_));
 sky130_fd_sc_hd__a31o_1 _2868_ (.A1(_1802_),
    .A2(_0895_),
    .A3(_0898_),
    .B1(_1801_),
    .X(_0900_));
 sky130_fd_sc_hd__o21ai_1 _2869_ (.A1(_0545_),
    .A2(_0890_),
    .B1(_0879_),
    .Y(_0901_));
 sky130_fd_sc_hd__o311a_1 _2870_ (.A1(net135),
    .A2(_1802_),
    .A3(_0890_),
    .B1(_0900_),
    .C1(_0879_),
    .X(_0902_));
 sky130_fd_sc_hd__o211ai_1 _2871_ (.A1(_0545_),
    .A2(_0890_),
    .B1(\acc[40] ),
    .C1(_0879_),
    .Y(_0903_));
 sky130_fd_sc_hd__o2111a_1 _2872_ (.A1(_0890_),
    .A2(_0545_),
    .B1(\acc[40] ),
    .C1(_0879_),
    .D1(_0900_),
    .X(_0904_));
 sky130_fd_sc_hd__o21bai_2 _2873_ (.A1(_0873_),
    .A2(_0904_),
    .B1_N(_0875_),
    .Y(_0905_));
 sky130_fd_sc_hd__o221ai_4 _2874_ (.A1(_0810_),
    .A2(_0843_),
    .B1(_0905_),
    .B2(_0847_),
    .C1(_0809_),
    .Y(_0906_));
 sky130_fd_sc_hd__and2_1 _2875_ (.A(_0724_),
    .B(_0725_),
    .X(_0907_));
 sky130_fd_sc_hd__nand2_1 _2876_ (.A(_0724_),
    .B(_0725_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21oi_1 _2877_ (.A1(_0783_),
    .A2(_0782_),
    .B1(\acc[44] ),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_1 _2878_ (.A(_0784_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nor3_1 _2879_ (.A(_0784_),
    .B(_0909_),
    .C(_0908_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand3_1 _2880_ (.A(_0664_),
    .B(_0907_),
    .C(_0910_),
    .Y(_0912_));
 sky130_fd_sc_hd__o21ai_1 _2881_ (.A1(_0786_),
    .A2(_0665_),
    .B1(_0659_),
    .Y(_0913_));
 sky130_fd_sc_hd__a31oi_1 _2882_ (.A1(_0906_),
    .A2(_0911_),
    .A3(_0664_),
    .B1(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__nor2_1 _2883_ (.A(_0873_),
    .B(_0875_),
    .Y(_0915_));
 sky130_fd_sc_hd__o21ai_1 _2884_ (.A1(_0899_),
    .A2(_0901_),
    .B1(_1789_),
    .Y(_0916_));
 sky130_fd_sc_hd__o21ai_1 _2885_ (.A1(_0899_),
    .A2(_0901_),
    .B1(\acc[40] ),
    .Y(_0917_));
 sky130_fd_sc_hd__o2111ai_1 _2886_ (.A1(_0890_),
    .A2(_0545_),
    .B1(_1789_),
    .C1(_0879_),
    .D1(_0900_),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _2887_ (.A(_0917_),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__o21ai_1 _2888_ (.A1(_0899_),
    .A2(_0903_),
    .B1(_0916_),
    .Y(_0920_));
 sky130_fd_sc_hd__o211a_1 _2889_ (.A1(_0899_),
    .A2(_0903_),
    .B1(_0916_),
    .C1(_0915_),
    .X(_0921_));
 sky130_fd_sc_hd__nand4_1 _2890_ (.A(_0812_),
    .B(_0844_),
    .C(_0915_),
    .D(_0919_),
    .Y(_0922_));
 sky130_fd_sc_hd__nor2_1 _2891_ (.A(_0912_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__nand4_1 _2892_ (.A(_0664_),
    .B(_0846_),
    .C(_0911_),
    .D(_0921_),
    .Y(_0924_));
 sky130_fd_sc_hd__a31o_1 _2893_ (.A1(_1801_),
    .A2(_0488_),
    .A3(_0539_),
    .B1(\acc[31] ),
    .X(_0925_));
 sky130_fd_sc_hd__nand3_2 _2894_ (.A(_0780_),
    .B(\count[4] ),
    .C(_0779_),
    .Y(_0926_));
 sky130_fd_sc_hd__nand3_1 _2895_ (.A(_1802_),
    .B(_0755_),
    .C(_0756_),
    .Y(_0927_));
 sky130_fd_sc_hd__o2111ai_2 _2896_ (.A1(\count[4] ),
    .A2(_0757_),
    .B1(_0926_),
    .C1(_1801_),
    .D1(\acc[28] ),
    .Y(_0928_));
 sky130_fd_sc_hd__nand3_2 _2897_ (.A(_0716_),
    .B(_0717_),
    .C(\count[4] ),
    .Y(_0929_));
 sky130_fd_sc_hd__nand3_2 _2898_ (.A(_1802_),
    .B(_0690_),
    .C(_0691_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand4_2 _2899_ (.A(_1801_),
    .B(_0929_),
    .C(_0930_),
    .D(\acc[29] ),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _2900_ (.A(_0928_),
    .B(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__a31o_1 _2901_ (.A1(_1801_),
    .A2(_0593_),
    .A3(_0639_),
    .B1(\acc[30] ),
    .X(_0933_));
 sky130_fd_sc_hd__a31o_1 _2902_ (.A1(_1801_),
    .A2(_0929_),
    .A3(_0930_),
    .B1(\acc[29] ),
    .X(_0934_));
 sky130_fd_sc_hd__nand4_1 _2903_ (.A(_1801_),
    .B(_0488_),
    .C(_0539_),
    .D(\acc[31] ),
    .Y(_0935_));
 sky130_fd_sc_hd__nand4_2 _2904_ (.A(_0593_),
    .B(\acc[30] ),
    .C(_1801_),
    .D(_0639_),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2_1 _2905_ (.A(_0935_),
    .B(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__a31o_1 _2906_ (.A1(_0932_),
    .A2(_0933_),
    .A3(_0934_),
    .B1(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__nand2_1 _2907_ (.A(_0925_),
    .B(_0935_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_1 _2908_ (.A(_0933_),
    .B(_0936_),
    .Y(_0940_));
 sky130_fd_sc_hd__a31o_1 _2909_ (.A1(_1801_),
    .A2(_0926_),
    .A3(_0927_),
    .B1(\acc[28] ),
    .X(_0941_));
 sky130_fd_sc_hd__nand2_1 _2910_ (.A(_0928_),
    .B(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand4_1 _2911_ (.A(_0928_),
    .B(_0931_),
    .C(_0934_),
    .D(_0941_),
    .Y(_0943_));
 sky130_fd_sc_hd__nand4_1 _2912_ (.A(_0925_),
    .B(_0933_),
    .C(_0935_),
    .D(_0936_),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_1 _2913_ (.A(_0943_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__a21oi_1 _2914_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_1802_),
    .Y(_0946_));
 sky130_fd_sc_hd__a21o_1 _2915_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_1802_),
    .X(_0947_));
 sky130_fd_sc_hd__a21oi_2 _2916_ (.A1(_0794_),
    .A2(_0797_),
    .B1(\count[4] ),
    .Y(_0948_));
 sky130_fd_sc_hd__o21a_1 _2917_ (.A1(\count[4] ),
    .A2(_0798_),
    .B1(_0947_),
    .X(_0949_));
 sky130_fd_sc_hd__o2111ai_4 _2918_ (.A1(\count[4] ),
    .A2(_0798_),
    .B1(_0947_),
    .C1(_1801_),
    .D1(\acc[27] ),
    .Y(_0950_));
 sky130_fd_sc_hd__o31a_1 _2919_ (.A1(net135),
    .A2(_0946_),
    .A3(_0948_),
    .B1(_1796_),
    .X(_0951_));
 sky130_fd_sc_hd__o31ai_2 _2920_ (.A1(net135),
    .A2(_0946_),
    .A3(_0948_),
    .B1(_1796_),
    .Y(_0952_));
 sky130_fd_sc_hd__o211ai_4 _2921_ (.A1(_1803_),
    .A2(_0831_),
    .B1(\count[4] ),
    .C1(_0833_),
    .Y(_0953_));
 sky130_fd_sc_hd__nand3_1 _2922_ (.A(_1802_),
    .B(_0821_),
    .C(_0822_),
    .Y(_0954_));
 sky130_fd_sc_hd__o2111ai_4 _2923_ (.A1(\count[4] ),
    .A2(_0823_),
    .B1(_0953_),
    .C1(_1801_),
    .D1(\acc[26] ),
    .Y(_0955_));
 sky130_fd_sc_hd__o41a_1 _2924_ (.A1(_1796_),
    .A2(net135),
    .A3(_0946_),
    .A4(_0948_),
    .B1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__a21o_1 _2925_ (.A1(_0950_),
    .A2(_0955_),
    .B1(_0951_),
    .X(_0957_));
 sky130_fd_sc_hd__nand2_1 _2926_ (.A(_0950_),
    .B(_0952_),
    .Y(_0958_));
 sky130_fd_sc_hd__a31o_1 _2927_ (.A1(_1801_),
    .A2(_0953_),
    .A3(_0954_),
    .B1(\acc[26] ),
    .X(_0959_));
 sky130_fd_sc_hd__and4_1 _2928_ (.A(_0950_),
    .B(_0952_),
    .C(_0955_),
    .D(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__nand4_2 _2929_ (.A(_0950_),
    .B(_0952_),
    .C(_0955_),
    .D(_0959_),
    .Y(_0961_));
 sky130_fd_sc_hd__a21o_1 _2930_ (.A1(_0862_),
    .A2(_0865_),
    .B1(_1802_),
    .X(_0962_));
 sky130_fd_sc_hd__nand3_1 _2931_ (.A(_1802_),
    .B(_0855_),
    .C(_0856_),
    .Y(_0963_));
 sky130_fd_sc_hd__a31o_1 _2932_ (.A1(_1801_),
    .A2(_0962_),
    .A3(_0963_),
    .B1(\acc[25] ),
    .X(_0964_));
 sky130_fd_sc_hd__a21o_1 _2933_ (.A1(_0895_),
    .A2(_0898_),
    .B1(_1802_),
    .X(_0965_));
 sky130_fd_sc_hd__nand3_2 _2934_ (.A(_1802_),
    .B(_0888_),
    .C(_0889_),
    .Y(_0966_));
 sky130_fd_sc_hd__o2111ai_2 _2935_ (.A1(\count[4] ),
    .A2(_0890_),
    .B1(\acc[24] ),
    .C1(_0965_),
    .D1(_1801_),
    .Y(_0967_));
 sky130_fd_sc_hd__nand4_1 _2936_ (.A(_0962_),
    .B(\acc[25] ),
    .C(_1801_),
    .D(_0963_),
    .Y(_0968_));
 sky130_fd_sc_hd__nand2_1 _2937_ (.A(_0967_),
    .B(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__nand2_1 _2938_ (.A(_0964_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__o22ai_2 _2939_ (.A1(_0951_),
    .A2(_0956_),
    .B1(_0961_),
    .B2(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__a22oi_4 _2940_ (.A1(_0925_),
    .A2(_0938_),
    .B1(_0971_),
    .B2(_0945_),
    .Y(_0972_));
 sky130_fd_sc_hd__a31o_1 _2941_ (.A1(_1801_),
    .A2(_0965_),
    .A3(_0966_),
    .B1(\acc[24] ),
    .X(_0973_));
 sky130_fd_sc_hd__nand2_1 _2942_ (.A(_0967_),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_1 _2943_ (.A(_0964_),
    .B(_0968_),
    .Y(_0975_));
 sky130_fd_sc_hd__nand4_1 _2944_ (.A(_0964_),
    .B(_0967_),
    .C(_0968_),
    .D(_0973_),
    .Y(_0976_));
 sky130_fd_sc_hd__nor4_2 _2945_ (.A(_0943_),
    .B(_0944_),
    .C(_0961_),
    .D(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__nand3_2 _2946_ (.A(_1803_),
    .B(_0601_),
    .C(_0611_),
    .Y(_0978_));
 sky130_fd_sc_hd__a31o_2 _2947_ (.A1(_1803_),
    .A2(_0601_),
    .A3(_0611_),
    .B1(_1802_),
    .X(_0979_));
 sky130_fd_sc_hd__nand3_2 _2948_ (.A(_1803_),
    .B(_0560_),
    .C(_0572_),
    .Y(_0980_));
 sky130_fd_sc_hd__nand3_2 _2949_ (.A(_0633_),
    .B(net136),
    .C(_0624_),
    .Y(_0981_));
 sky130_fd_sc_hd__nand3_4 _2950_ (.A(_1802_),
    .B(_0980_),
    .C(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__a31oi_1 _2951_ (.A1(_1801_),
    .A2(_0979_),
    .A3(_0982_),
    .B1(\acc[22] ),
    .Y(_0983_));
 sky130_fd_sc_hd__a31o_1 _2952_ (.A1(_1801_),
    .A2(_0979_),
    .A3(_0982_),
    .B1(\acc[22] ),
    .X(_0984_));
 sky130_fd_sc_hd__and4_1 _2953_ (.A(_1801_),
    .B(_0979_),
    .C(_0982_),
    .D(\acc[22] ),
    .X(_0985_));
 sky130_fd_sc_hd__nand4_1 _2954_ (.A(_1801_),
    .B(_0979_),
    .C(_0982_),
    .D(\acc[22] ),
    .Y(_0986_));
 sky130_fd_sc_hd__nor2_1 _2955_ (.A(_0983_),
    .B(_0985_),
    .Y(_0987_));
 sky130_fd_sc_hd__and3_1 _2956_ (.A(_1803_),
    .B(_0470_),
    .C(_0482_),
    .X(_0988_));
 sky130_fd_sc_hd__a31o_1 _2957_ (.A1(_1803_),
    .A2(_0470_),
    .A3(_0482_),
    .B1(_1802_),
    .X(_0989_));
 sky130_fd_sc_hd__nand3_1 _2958_ (.A(_1803_),
    .B(_0500_),
    .C(_0511_),
    .Y(_0990_));
 sky130_fd_sc_hd__nand3_2 _2959_ (.A(_0457_),
    .B(\count[3] ),
    .C(_0447_),
    .Y(_0991_));
 sky130_fd_sc_hd__nand3_4 _2960_ (.A(_1802_),
    .B(_0990_),
    .C(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__o2111a_1 _2961_ (.A1(_1802_),
    .A2(_0988_),
    .B1(_0992_),
    .C1(_1801_),
    .D1(\acc[23] ),
    .X(_0993_));
 sky130_fd_sc_hd__o2111ai_1 _2962_ (.A1(_1802_),
    .A2(_0988_),
    .B1(_0992_),
    .C1(_1801_),
    .D1(\acc[23] ),
    .Y(_0994_));
 sky130_fd_sc_hd__a31oi_1 _2963_ (.A1(_1801_),
    .A2(_0989_),
    .A3(_0992_),
    .B1(\acc[23] ),
    .Y(_0995_));
 sky130_fd_sc_hd__a31o_1 _2964_ (.A1(_1801_),
    .A2(_0989_),
    .A3(_0992_),
    .B1(\acc[23] ),
    .X(_0996_));
 sky130_fd_sc_hd__nor2_1 _2965_ (.A(_0993_),
    .B(_0995_),
    .Y(_0997_));
 sky130_fd_sc_hd__nand4_1 _2966_ (.A(_0984_),
    .B(_0986_),
    .C(_0994_),
    .D(_0996_),
    .Y(_0998_));
 sky130_fd_sc_hd__a21oi_4 _2967_ (.A1(_0764_),
    .A2(_0765_),
    .B1(net136),
    .Y(_0999_));
 sky130_fd_sc_hd__a21o_1 _2968_ (.A1(_0764_),
    .A2(_0765_),
    .B1(net136),
    .X(_1000_));
 sky130_fd_sc_hd__a31o_1 _2969_ (.A1(_1803_),
    .A2(_0758_),
    .A3(_0763_),
    .B1(_1802_),
    .X(_1001_));
 sky130_fd_sc_hd__nand3_1 _2970_ (.A(_0777_),
    .B(\count[3] ),
    .C(_0776_),
    .Y(_1002_));
 sky130_fd_sc_hd__nand3_1 _2971_ (.A(_1803_),
    .B(_0741_),
    .C(_0742_),
    .Y(_1003_));
 sky130_fd_sc_hd__nand3_1 _2972_ (.A(_1803_),
    .B(_0736_),
    .C(_0740_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand3_1 _2973_ (.A(_0771_),
    .B(_0775_),
    .C(\count[3] ),
    .Y(_1005_));
 sky130_fd_sc_hd__nand3_4 _2974_ (.A(_1802_),
    .B(_1004_),
    .C(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__o21ai_2 _2975_ (.A1(_1802_),
    .A2(_0999_),
    .B1(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__o2111a_1 _2976_ (.A1(_0999_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[20] ),
    .D1(_1006_),
    .X(_1008_));
 sky130_fd_sc_hd__o2111ai_2 _2977_ (.A1(_0999_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[20] ),
    .D1(_1006_),
    .Y(_1009_));
 sky130_fd_sc_hd__a31oi_1 _2978_ (.A1(_1801_),
    .A2(_1001_),
    .A3(_1006_),
    .B1(\acc[20] ),
    .Y(_1010_));
 sky130_fd_sc_hd__a31o_1 _2979_ (.A1(_1801_),
    .A2(_1001_),
    .A3(_1006_),
    .B1(\acc[20] ),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_1 _2980_ (.A(_1008_),
    .B(_1010_),
    .Y(_1012_));
 sky130_fd_sc_hd__nand2_1 _2981_ (.A(_1009_),
    .B(_1011_),
    .Y(_1013_));
 sky130_fd_sc_hd__o211a_1 _2982_ (.A1(_0711_),
    .A2(_1804_),
    .B1(_1803_),
    .C1(_0710_),
    .X(_1014_));
 sky130_fd_sc_hd__a21o_1 _2983_ (.A1(_0713_),
    .A2(_0714_),
    .B1(net136),
    .X(_1015_));
 sky130_fd_sc_hd__a31o_1 _2984_ (.A1(_1803_),
    .A2(_0710_),
    .A3(_0712_),
    .B1(_1802_),
    .X(_1016_));
 sky130_fd_sc_hd__nand3_1 _2985_ (.A(_0703_),
    .B(_0704_),
    .C(net136),
    .Y(_1017_));
 sky130_fd_sc_hd__nand3_1 _2986_ (.A(_0697_),
    .B(_0702_),
    .C(\count[3] ),
    .Y(_1018_));
 sky130_fd_sc_hd__nand3_1 _2987_ (.A(_1803_),
    .B(_0669_),
    .C(_0674_),
    .Y(_1019_));
 sky130_fd_sc_hd__nand3_4 _2988_ (.A(_1802_),
    .B(_1018_),
    .C(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__o2111a_1 _2989_ (.A1(_1802_),
    .A2(_1014_),
    .B1(\acc[21] ),
    .C1(_1020_),
    .D1(_1801_),
    .X(_1021_));
 sky130_fd_sc_hd__o2111ai_1 _2990_ (.A1(_1802_),
    .A2(_1014_),
    .B1(\acc[21] ),
    .C1(_1020_),
    .D1(_1801_),
    .Y(_1022_));
 sky130_fd_sc_hd__a31oi_1 _2991_ (.A1(_1801_),
    .A2(_1016_),
    .A3(_1020_),
    .B1(\acc[21] ),
    .Y(_1023_));
 sky130_fd_sc_hd__a31o_1 _2992_ (.A1(_1801_),
    .A2(_1016_),
    .A3(_1020_),
    .B1(\acc[21] ),
    .X(_1024_));
 sky130_fd_sc_hd__nor2_1 _2993_ (.A(_1021_),
    .B(_1023_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand4_1 _2994_ (.A(_1009_),
    .B(_1011_),
    .C(_1022_),
    .D(_1024_),
    .Y(_1026_));
 sky130_fd_sc_hd__nand4_1 _2995_ (.A(_0987_),
    .B(_0997_),
    .C(_1012_),
    .D(_1025_),
    .Y(_1027_));
 sky130_fd_sc_hd__and3_2 _2996_ (.A(_0711_),
    .B(_1804_),
    .C(_1803_),
    .X(_1028_));
 sky130_fd_sc_hd__o2111ai_2 _2997_ (.A1(\q[0] ),
    .A2(_1806_),
    .B1(_1805_),
    .C1(_1803_),
    .D1(_0863_),
    .Y(_1029_));
 sky130_fd_sc_hd__nand3_1 _2998_ (.A(_0860_),
    .B(_0861_),
    .C(net136),
    .Y(_1030_));
 sky130_fd_sc_hd__nand3_1 _2999_ (.A(_1803_),
    .B(_0850_),
    .C(_0851_),
    .Y(_1031_));
 sky130_fd_sc_hd__nand3_1 _3000_ (.A(_0859_),
    .B(\count[3] ),
    .C(_0858_),
    .Y(_1032_));
 sky130_fd_sc_hd__nand3_1 _3001_ (.A(_1803_),
    .B(_0848_),
    .C(_0849_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand3_4 _3002_ (.A(_1802_),
    .B(_1032_),
    .C(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__a21oi_1 _3003_ (.A1(_1029_),
    .A2(\count[4] ),
    .B1(net135),
    .Y(_1035_));
 sky130_fd_sc_hd__a21oi_2 _3004_ (.A1(_1034_),
    .A2(_1035_),
    .B1(\acc[17] ),
    .Y(_1036_));
 sky130_fd_sc_hd__a21o_1 _3005_ (.A1(_1034_),
    .A2(_1035_),
    .B1(\acc[17] ),
    .X(_1037_));
 sky130_fd_sc_hd__o2111a_1 _3006_ (.A1(_1028_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[17] ),
    .D1(_1034_),
    .X(_1038_));
 sky130_fd_sc_hd__o2111ai_1 _3007_ (.A1(_1028_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[17] ),
    .D1(_1034_),
    .Y(_1039_));
 sky130_fd_sc_hd__nand3_1 _3008_ (.A(_1803_),
    .B(_0882_),
    .C(_0883_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand3_1 _3009_ (.A(_0893_),
    .B(_0894_),
    .C(\count[3] ),
    .Y(_1041_));
 sky130_fd_sc_hd__nand3_1 _3010_ (.A(_0891_),
    .B(_0892_),
    .C(\count[3] ),
    .Y(_1042_));
 sky130_fd_sc_hd__nand3_1 _3011_ (.A(_1803_),
    .B(_0880_),
    .C(_0881_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand3_4 _3012_ (.A(_1802_),
    .B(_1042_),
    .C(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__and3_2 _3013_ (.A(_0594_),
    .B(_0896_),
    .C(_1803_),
    .X(_1045_));
 sky130_fd_sc_hd__or4_1 _3014_ (.A(net136),
    .B(net137),
    .C(net138),
    .D(_0595_),
    .X(_1046_));
 sky130_fd_sc_hd__o21a_1 _3015_ (.A1(_1802_),
    .A2(_1045_),
    .B1(_1801_),
    .X(_1047_));
 sky130_fd_sc_hd__o2111a_1 _3016_ (.A1(_1045_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[16] ),
    .D1(_1044_),
    .X(_1048_));
 sky130_fd_sc_hd__o2111ai_4 _3017_ (.A1(_1045_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[16] ),
    .D1(_1044_),
    .Y(_1049_));
 sky130_fd_sc_hd__o21ai_2 _3018_ (.A1(_1049_),
    .A2(_1036_),
    .B1(_1039_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand3_1 _3019_ (.A(_1803_),
    .B(_0816_),
    .C(_0817_),
    .Y(_1051_));
 sky130_fd_sc_hd__nand3_1 _3020_ (.A(_0827_),
    .B(_0828_),
    .C(\count[3] ),
    .Y(_1052_));
 sky130_fd_sc_hd__nand3_1 _3021_ (.A(_0826_),
    .B(net136),
    .C(_0825_),
    .Y(_1053_));
 sky130_fd_sc_hd__nand3_1 _3022_ (.A(_1803_),
    .B(_0814_),
    .C(_0815_),
    .Y(_1054_));
 sky130_fd_sc_hd__nand3_4 _3023_ (.A(_1802_),
    .B(_1053_),
    .C(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__and3_1 _3024_ (.A(_0830_),
    .B(_0598_),
    .C(_1803_),
    .X(_1056_));
 sky130_fd_sc_hd__o2111ai_4 _3025_ (.A1(_0594_),
    .A2(_1805_),
    .B1(_1804_),
    .C1(_1803_),
    .D1(_0598_),
    .Y(_1057_));
 sky130_fd_sc_hd__a31o_1 _3026_ (.A1(_0830_),
    .A2(_0598_),
    .A3(_1803_),
    .B1(_1802_),
    .X(_1058_));
 sky130_fd_sc_hd__a21oi_1 _3027_ (.A1(_1057_),
    .A2(\count[4] ),
    .B1(net135),
    .Y(_1059_));
 sky130_fd_sc_hd__a21oi_1 _3028_ (.A1(_1055_),
    .A2(_1059_),
    .B1(\acc[18] ),
    .Y(_1060_));
 sky130_fd_sc_hd__a31o_1 _3029_ (.A1(_1801_),
    .A2(_1055_),
    .A3(_1058_),
    .B1(\acc[18] ),
    .X(_1061_));
 sky130_fd_sc_hd__o2111a_1 _3030_ (.A1(_1056_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[18] ),
    .D1(_1055_),
    .X(_1062_));
 sky130_fd_sc_hd__o2111ai_1 _3031_ (.A1(_1056_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[18] ),
    .D1(_1055_),
    .Y(_1063_));
 sky130_fd_sc_hd__nor2_1 _3032_ (.A(_1060_),
    .B(_1062_),
    .Y(_1064_));
 sky130_fd_sc_hd__o2111a_2 _3033_ (.A1(_1805_),
    .A2(_0477_),
    .B1(_0474_),
    .C1(_1803_),
    .D1(_1804_),
    .X(_1065_));
 sky130_fd_sc_hd__a41o_1 _3034_ (.A1(_1803_),
    .A2(_1804_),
    .A3(_0474_),
    .A4(_0479_),
    .B1(_1802_),
    .X(_1066_));
 sky130_fd_sc_hd__nand3_1 _3035_ (.A(_0801_),
    .B(_0802_),
    .C(net136),
    .Y(_1067_));
 sky130_fd_sc_hd__nand3_1 _3036_ (.A(_0800_),
    .B(\count[3] ),
    .C(_0799_),
    .Y(_1068_));
 sky130_fd_sc_hd__nand3_1 _3037_ (.A(_1803_),
    .B(_0789_),
    .C(_0790_),
    .Y(_1069_));
 sky130_fd_sc_hd__nand3_4 _3038_ (.A(_1802_),
    .B(_1068_),
    .C(_1069_),
    .Y(_1070_));
 sky130_fd_sc_hd__o21a_1 _3039_ (.A1(_1802_),
    .A2(_1065_),
    .B1(_1801_),
    .X(_1071_));
 sky130_fd_sc_hd__o2111a_1 _3040_ (.A1(_1065_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[19] ),
    .D1(_1070_),
    .X(_1072_));
 sky130_fd_sc_hd__o2111ai_4 _3041_ (.A1(_1065_),
    .A2(_1802_),
    .B1(_1801_),
    .C1(\acc[19] ),
    .D1(_1070_),
    .Y(_1073_));
 sky130_fd_sc_hd__a21oi_1 _3042_ (.A1(_1071_),
    .A2(_1070_),
    .B1(\acc[19] ),
    .Y(_1074_));
 sky130_fd_sc_hd__a31o_1 _3043_ (.A1(_1801_),
    .A2(_1066_),
    .A3(_1070_),
    .B1(\acc[19] ),
    .X(_1075_));
 sky130_fd_sc_hd__nor2_1 _3044_ (.A(_1072_),
    .B(_1074_),
    .Y(_1076_));
 sky130_fd_sc_hd__o21ai_1 _3045_ (.A1(_1063_),
    .A2(_1074_),
    .B1(_1073_),
    .Y(_1077_));
 sky130_fd_sc_hd__a41oi_4 _3046_ (.A1(_1050_),
    .A2(_1064_),
    .A3(_1073_),
    .A4(_1075_),
    .B1(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__a21oi_1 _3047_ (.A1(_1009_),
    .A2(_1022_),
    .B1(_1023_),
    .Y(_1079_));
 sky130_fd_sc_hd__o21ai_1 _3048_ (.A1(_0986_),
    .A2(_0995_),
    .B1(_0994_),
    .Y(_1080_));
 sky130_fd_sc_hd__a31oi_1 _3049_ (.A1(_0987_),
    .A2(_0997_),
    .A3(_1079_),
    .B1(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__o21ai_2 _3050_ (.A1(_1027_),
    .A2(_1078_),
    .B1(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__a21oi_1 _3051_ (.A1(_1044_),
    .A2(_1047_),
    .B1(\acc[16] ),
    .Y(_1083_));
 sky130_fd_sc_hd__a21o_1 _3052_ (.A1(_1044_),
    .A2(_1047_),
    .B1(\acc[16] ),
    .X(_1084_));
 sky130_fd_sc_hd__nor2_1 _3053_ (.A(_1048_),
    .B(_1083_),
    .Y(_1085_));
 sky130_fd_sc_hd__nor2_1 _3054_ (.A(_1036_),
    .B(_1038_),
    .Y(_1086_));
 sky130_fd_sc_hd__nand4_1 _3055_ (.A(_1064_),
    .B(_1076_),
    .C(_1085_),
    .D(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__nor3_1 _3056_ (.A(_0998_),
    .B(_1026_),
    .C(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__nand4_2 _3057_ (.A(_0460_),
    .B(_0486_),
    .C(_0648_),
    .D(\acc[15] ),
    .Y(_1089_));
 sky130_fd_sc_hd__a31o_1 _3058_ (.A1(_0460_),
    .A2(_0486_),
    .A3(_0648_),
    .B1(\acc[15] ),
    .X(_1090_));
 sky130_fd_sc_hd__nand4_1 _3059_ (.A(_0613_),
    .B(_0636_),
    .C(_0648_),
    .D(\acc[14] ),
    .Y(_1091_));
 sky130_fd_sc_hd__a31o_1 _3060_ (.A1(_0613_),
    .A2(_0636_),
    .A3(_0648_),
    .B1(\acc[14] ),
    .X(_1092_));
 sky130_fd_sc_hd__nand2_1 _3061_ (.A(_1091_),
    .B(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__nand4_1 _3062_ (.A(_1089_),
    .B(_1090_),
    .C(_1091_),
    .D(_1092_),
    .Y(_1094_));
 sky130_fd_sc_hd__a31o_1 _3063_ (.A1(_0778_),
    .A2(_0648_),
    .A3(_0766_),
    .B1(\acc[12] ),
    .X(_1095_));
 sky130_fd_sc_hd__nand4_4 _3064_ (.A(_0778_),
    .B(\acc[12] ),
    .C(_0766_),
    .D(_0648_),
    .Y(_1096_));
 sky130_fd_sc_hd__nand2_1 _3065_ (.A(_1095_),
    .B(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__a31oi_1 _3066_ (.A1(_0705_),
    .A2(_0715_),
    .A3(_0648_),
    .B1(\acc[13] ),
    .Y(_1098_));
 sky130_fd_sc_hd__a31o_1 _3067_ (.A1(_0705_),
    .A2(_0715_),
    .A3(_0648_),
    .B1(\acc[13] ),
    .X(_1099_));
 sky130_fd_sc_hd__nand4_2 _3068_ (.A(_0705_),
    .B(_0715_),
    .C(\acc[13] ),
    .D(_0648_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _3069_ (.A(_1099_),
    .B(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__nand4_1 _3070_ (.A(_1095_),
    .B(_1096_),
    .C(_1099_),
    .D(_1100_),
    .Y(_1102_));
 sky130_fd_sc_hd__nor2_1 _3071_ (.A(_1094_),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__a21o_1 _3072_ (.A1(_1096_),
    .A2(_1100_),
    .B1(_1098_),
    .X(_1104_));
 sky130_fd_sc_hd__nand2b_1 _3073_ (.A_N(_1091_),
    .B(_1090_),
    .Y(_1105_));
 sky130_fd_sc_hd__o211a_1 _3074_ (.A1(_1094_),
    .A2(_1104_),
    .B1(_1105_),
    .C1(_1089_),
    .X(_1106_));
 sky130_fd_sc_hd__nor3_4 _3075_ (.A(net135),
    .B(\count[4] ),
    .C(\count[3] ),
    .Y(_1107_));
 sky130_fd_sc_hd__or4_1 _3076_ (.A(_1800_),
    .B(net135),
    .C(\count[4] ),
    .D(_1000_),
    .X(_1108_));
 sky130_fd_sc_hd__and4_2 _3077_ (.A(_1107_),
    .B(_0763_),
    .C(_0758_),
    .D(_1800_),
    .X(_1109_));
 sky130_fd_sc_hd__a31oi_4 _3078_ (.A1(_0758_),
    .A2(_0763_),
    .A3(_1107_),
    .B1(_1800_),
    .Y(_1110_));
 sky130_fd_sc_hd__a31o_2 _3079_ (.A1(_1065_),
    .A2(_1802_),
    .A3(_1801_),
    .B1(\acc[3] ),
    .X(_1111_));
 sky130_fd_sc_hd__nand2_1 _3080_ (.A(\acc[3] ),
    .B(_1065_),
    .Y(_1112_));
 sky130_fd_sc_hd__a31o_1 _3081_ (.A1(_0830_),
    .A2(_1107_),
    .A3(_0598_),
    .B1(\acc[2] ),
    .X(_1113_));
 sky130_fd_sc_hd__nand4_1 _3082_ (.A(\acc[2] ),
    .B(_0830_),
    .C(_1107_),
    .D(_0598_),
    .Y(_1114_));
 sky130_fd_sc_hd__a41oi_4 _3083_ (.A1(_1805_),
    .A2(_0863_),
    .A3(_1107_),
    .A4(_0475_),
    .B1(\acc[1] ),
    .Y(_1115_));
 sky130_fd_sc_hd__nand4_2 _3084_ (.A(\acc[0] ),
    .B(_0594_),
    .C(_0896_),
    .D(_1107_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand4_1 _3085_ (.A(\acc[1] ),
    .B(_0711_),
    .C(_1107_),
    .D(_1804_),
    .Y(_1117_));
 sky130_fd_sc_hd__a21oi_1 _3086_ (.A1(_1116_),
    .A2(_1117_),
    .B1(_1115_),
    .Y(_1118_));
 sky130_fd_sc_hd__o211ai_1 _3087_ (.A1(_1116_),
    .A2(_1115_),
    .B1(_1114_),
    .C1(_1117_),
    .Y(_1119_));
 sky130_fd_sc_hd__and2_1 _3088_ (.A(_1113_),
    .B(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__o2bb2ai_2 _3089_ (.A1_N(_1113_),
    .A2_N(_1119_),
    .B1(_0649_),
    .B2(_1112_),
    .Y(_1121_));
 sky130_fd_sc_hd__o211ai_2 _3090_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1111_),
    .C1(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__and4_1 _3091_ (.A(_0710_),
    .B(_0712_),
    .C(_1107_),
    .D(\acc[5] ),
    .X(_1123_));
 sky130_fd_sc_hd__a31o_1 _3092_ (.A1(_0710_),
    .A2(_0712_),
    .A3(_1107_),
    .B1(\acc[5] ),
    .X(_1124_));
 sky130_fd_sc_hd__a31o_1 _3093_ (.A1(_0710_),
    .A2(_0712_),
    .A3(_1107_),
    .B1(_1799_),
    .X(_1125_));
 sky130_fd_sc_hd__o2111ai_2 _3094_ (.A1(_1804_),
    .A2(_0711_),
    .B1(_1107_),
    .C1(_0710_),
    .D1(_1799_),
    .Y(_1126_));
 sky130_fd_sc_hd__nand2_1 _3095_ (.A(_1125_),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__o2111ai_4 _3096_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1111_),
    .C1(_1127_),
    .D1(_1121_),
    .Y(_1128_));
 sky130_fd_sc_hd__a41oi_4 _3097_ (.A1(_1124_),
    .A2(_0999_),
    .A3(_0648_),
    .A4(\acc[4] ),
    .B1(_1123_),
    .Y(_1129_));
 sky130_fd_sc_hd__a31o_1 _3098_ (.A1(_0470_),
    .A2(_0482_),
    .A3(_1107_),
    .B1(\acc[7] ),
    .X(_1130_));
 sky130_fd_sc_hd__or3b_1 _3099_ (.A(net135),
    .B(\count[4] ),
    .C_N(\acc[6] ),
    .X(_1131_));
 sky130_fd_sc_hd__and4_1 _3100_ (.A(_0601_),
    .B(_0611_),
    .C(_1107_),
    .D(\acc[6] ),
    .X(_1132_));
 sky130_fd_sc_hd__nand2_1 _3101_ (.A(_1132_),
    .B(_1130_),
    .Y(_1133_));
 sky130_fd_sc_hd__nand4_2 _3102_ (.A(_0470_),
    .B(_0482_),
    .C(_1107_),
    .D(\acc[7] ),
    .Y(_1134_));
 sky130_fd_sc_hd__a31o_1 _3103_ (.A1(_0601_),
    .A2(_0611_),
    .A3(_1107_),
    .B1(\acc[6] ),
    .X(_1135_));
 sky130_fd_sc_hd__a21boi_1 _3104_ (.A1(_1130_),
    .A2(_1135_),
    .B1_N(_1134_),
    .Y(_1136_));
 sky130_fd_sc_hd__a41oi_4 _3105_ (.A1(_1128_),
    .A2(_1129_),
    .A3(_1133_),
    .A4(_1134_),
    .B1(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__a31oi_1 _3106_ (.A1(_0803_),
    .A2(_0804_),
    .A3(_0648_),
    .B1(\acc[11] ),
    .Y(_1138_));
 sky130_fd_sc_hd__a31o_1 _3107_ (.A1(_0803_),
    .A2(_0804_),
    .A3(_0648_),
    .B1(\acc[11] ),
    .X(_1139_));
 sky130_fd_sc_hd__nand4_2 _3108_ (.A(_0803_),
    .B(_0804_),
    .C(\acc[11] ),
    .D(_0648_),
    .Y(_1140_));
 sky130_fd_sc_hd__a31o_1 _3109_ (.A1(_0829_),
    .A2(_0832_),
    .A3(_0648_),
    .B1(\acc[10] ),
    .X(_1141_));
 sky130_fd_sc_hd__and4_1 _3110_ (.A(_0829_),
    .B(_0832_),
    .C(\acc[10] ),
    .D(_0648_),
    .X(_1142_));
 sky130_fd_sc_hd__nand4_1 _3111_ (.A(_0829_),
    .B(_0832_),
    .C(\acc[10] ),
    .D(_0648_),
    .Y(_1143_));
 sky130_fd_sc_hd__and2_1 _3112_ (.A(_1141_),
    .B(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__nand4_1 _3113_ (.A(_1139_),
    .B(_1140_),
    .C(_1141_),
    .D(_1143_),
    .Y(_1145_));
 sky130_fd_sc_hd__a31o_1 _3114_ (.A1(_0895_),
    .A2(_0898_),
    .A3(_0648_),
    .B1(\acc[8] ),
    .X(_1146_));
 sky130_fd_sc_hd__o2111ai_4 _3115_ (.A1(_1803_),
    .A2(_0897_),
    .B1(_0648_),
    .C1(\acc[8] ),
    .D1(_0895_),
    .Y(_1147_));
 sky130_fd_sc_hd__a31o_1 _3116_ (.A1(_0862_),
    .A2(_0865_),
    .A3(_0648_),
    .B1(\acc[9] ),
    .X(_1148_));
 sky130_fd_sc_hd__nand4_1 _3117_ (.A(_0862_),
    .B(_0865_),
    .C(\acc[9] ),
    .D(_0648_),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _3118_ (.A(_1148_),
    .B(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand4_1 _3119_ (.A(_1146_),
    .B(_1147_),
    .C(_1148_),
    .D(_1149_),
    .Y(_1151_));
 sky130_fd_sc_hd__nor2_1 _3120_ (.A(_1145_),
    .B(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _3121_ (.A(_1137_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_1 _3122_ (.A(_1147_),
    .B(_1149_),
    .Y(_1154_));
 sky130_fd_sc_hd__nand2_1 _3123_ (.A(_1148_),
    .B(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__and2_1 _3124_ (.A(_1140_),
    .B(_1143_),
    .X(_1156_));
 sky130_fd_sc_hd__o221a_1 _3125_ (.A1(_1143_),
    .A2(_1138_),
    .B1(_1155_),
    .B2(_1145_),
    .C1(_1140_),
    .X(_1157_));
 sky130_fd_sc_hd__o22ai_1 _3126_ (.A1(_1138_),
    .A2(_1156_),
    .B1(_1155_),
    .B2(_1145_),
    .Y(_1158_));
 sky130_fd_sc_hd__nand3_2 _3127_ (.A(_1103_),
    .B(_1137_),
    .C(_1152_),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_1 _3128_ (.A(_1103_),
    .B(_1158_),
    .Y(_1160_));
 sky130_fd_sc_hd__nand3_4 _3129_ (.A(_1159_),
    .B(_1160_),
    .C(_1106_),
    .Y(_1161_));
 sky130_fd_sc_hd__a21oi_2 _3130_ (.A1(_1088_),
    .A2(_1161_),
    .B1(_1082_),
    .Y(_1162_));
 sky130_fd_sc_hd__nand2_2 _3131_ (.A(_1082_),
    .B(_0977_),
    .Y(_1163_));
 sky130_fd_sc_hd__nand3_2 _3132_ (.A(_0977_),
    .B(_1088_),
    .C(_1161_),
    .Y(_1164_));
 sky130_fd_sc_hd__nand3_4 _3133_ (.A(_1163_),
    .B(_1164_),
    .C(_0972_),
    .Y(_1165_));
 sky130_fd_sc_hd__o21ai_2 _3134_ (.A1(_1804_),
    .A2(_0719_),
    .B1(_1803_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand3_2 _3135_ (.A(_0687_),
    .B(_0688_),
    .C(net136),
    .Y(_1167_));
 sky130_fd_sc_hd__nand4_4 _3136_ (.A(_1801_),
    .B(_1802_),
    .C(_1166_),
    .D(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__a211o_1 _3137_ (.A1(_0713_),
    .A2(_0714_),
    .B1(net136),
    .C1(_0645_),
    .X(_1169_));
 sky130_fd_sc_hd__o211ai_4 _3138_ (.A1(net136),
    .A2(_0677_),
    .B1(_1017_),
    .C1(_0544_),
    .Y(_1170_));
 sky130_fd_sc_hd__o211ai_2 _3139_ (.A1(_0645_),
    .A2(_1015_),
    .B1(_1168_),
    .C1(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__and4_1 _3140_ (.A(_1791_),
    .B(_1168_),
    .C(_1169_),
    .D(_1170_),
    .X(_1172_));
 sky130_fd_sc_hd__o2111ai_4 _3141_ (.A1(_0645_),
    .A2(_1015_),
    .B1(_1168_),
    .C1(_1170_),
    .D1(_1791_),
    .Y(_1173_));
 sky130_fd_sc_hd__a31o_1 _3142_ (.A1(_1168_),
    .A2(_1169_),
    .A3(_1170_),
    .B1(_1791_),
    .X(_1174_));
 sky130_fd_sc_hd__o21a_1 _3143_ (.A1(_1804_),
    .A2(_0727_),
    .B1(_1803_),
    .X(_1175_));
 sky130_fd_sc_hd__and3_1 _3144_ (.A(_0754_),
    .B(net136),
    .C(_0753_),
    .X(_1176_));
 sky130_fd_sc_hd__nand3_1 _3145_ (.A(_0754_),
    .B(net136),
    .C(_0753_),
    .Y(_1177_));
 sky130_fd_sc_hd__o211ai_4 _3146_ (.A1(net136),
    .A2(_0729_),
    .B1(_0648_),
    .C1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__nand4_4 _3147_ (.A(_1801_),
    .B(_1003_),
    .C(\count[4] ),
    .D(_1002_),
    .Y(_1179_));
 sky130_fd_sc_hd__o211ai_2 _3148_ (.A1(_0645_),
    .A2(_1000_),
    .B1(_1178_),
    .C1(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__and2_1 _3149_ (.A(_1180_),
    .B(\acc[36] ),
    .X(_1181_));
 sky130_fd_sc_hd__nand2_1 _3150_ (.A(_1180_),
    .B(\acc[36] ),
    .Y(_1182_));
 sky130_fd_sc_hd__o2111ai_4 _3151_ (.A1(_0645_),
    .A2(_1000_),
    .B1(_1178_),
    .C1(_1179_),
    .D1(_1792_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _3152_ (.A(_1182_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__nand4_1 _3153_ (.A(_1173_),
    .B(_1174_),
    .C(_1182_),
    .D(_1183_),
    .Y(_1185_));
 sky130_fd_sc_hd__a21o_1 _3154_ (.A1(_0980_),
    .A2(_0981_),
    .B1(_0545_),
    .X(_1186_));
 sky130_fd_sc_hd__nand3_1 _3155_ (.A(_0590_),
    .B(net136),
    .C(_0581_),
    .Y(_1187_));
 sky130_fd_sc_hd__o31ai_4 _3156_ (.A1(net136),
    .A2(_1804_),
    .A3(_0547_),
    .B1(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__a2bb2oi_1 _3157_ (.A1_N(_0645_),
    .A2_N(_0978_),
    .B1(_0648_),
    .B2(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__a21o_1 _3158_ (.A1(_1189_),
    .A2(_1186_),
    .B1(_1790_),
    .X(_1190_));
 sky130_fd_sc_hd__nand3_1 _3159_ (.A(_1189_),
    .B(_1186_),
    .C(_1790_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand2_1 _3160_ (.A(_1190_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__inv_2 _3161_ (.A(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__o2111ai_2 _3162_ (.A1(net136),
    .A2(_0514_),
    .B1(_0991_),
    .C1(\count[4] ),
    .D1(_1801_),
    .Y(_1194_));
 sky130_fd_sc_hd__a31oi_1 _3163_ (.A1(_0534_),
    .A2(net136),
    .A3(_0525_),
    .B1(_0649_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand4_1 _3164_ (.A(_1802_),
    .B(_1803_),
    .C(_0470_),
    .D(_0482_),
    .Y(_1196_));
 sky130_fd_sc_hd__a21oi_1 _3165_ (.A1(net135),
    .A2(_1196_),
    .B1(_1195_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand3_1 _3166_ (.A(\acc[39] ),
    .B(_1197_),
    .C(_1194_),
    .Y(_1198_));
 sky130_fd_sc_hd__a21o_1 _3167_ (.A1(_1197_),
    .A2(_1194_),
    .B1(\acc[39] ),
    .X(_1199_));
 sky130_fd_sc_hd__nand2_1 _3168_ (.A(_1198_),
    .B(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nand4_1 _3169_ (.A(_1190_),
    .B(_1191_),
    .C(_1198_),
    .D(_1199_),
    .Y(_1201_));
 sky130_fd_sc_hd__nor2_1 _3170_ (.A(_1185_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__o211ai_2 _3171_ (.A1(net136),
    .A2(_0793_),
    .B1(_1067_),
    .C1(_0544_),
    .Y(_1203_));
 sky130_fd_sc_hd__a2111o_1 _3172_ (.A1(_0480_),
    .A2(_0481_),
    .B1(_0645_),
    .C1(net137),
    .D1(net136),
    .X(_1204_));
 sky130_fd_sc_hd__nand3_2 _3173_ (.A(_0795_),
    .B(_0796_),
    .C(net136),
    .Y(_1205_));
 sky130_fd_sc_hd__o2111ai_4 _3174_ (.A1(net136),
    .A2(_0787_),
    .B1(_1205_),
    .C1(_1802_),
    .D1(_1801_),
    .Y(_1206_));
 sky130_fd_sc_hd__a31o_2 _3175_ (.A1(_1203_),
    .A2(_1204_),
    .A3(_1206_),
    .B1(_1793_),
    .X(_1207_));
 sky130_fd_sc_hd__and4_1 _3176_ (.A(_1793_),
    .B(_1203_),
    .C(_1204_),
    .D(_1206_),
    .X(_1208_));
 sky130_fd_sc_hd__nand4_2 _3177_ (.A(_1793_),
    .B(_1203_),
    .C(_1204_),
    .D(_1206_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2_1 _3178_ (.A(_1207_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__nand3_2 _3179_ (.A(_0820_),
    .B(\count[3] ),
    .C(_0819_),
    .Y(_1211_));
 sky130_fd_sc_hd__o211ai_4 _3180_ (.A1(_0547_),
    .A2(\count[2] ),
    .B1(_1803_),
    .C1(_0834_),
    .Y(_1212_));
 sky130_fd_sc_hd__nand4_4 _3181_ (.A(_1801_),
    .B(_1802_),
    .C(_1211_),
    .D(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__nand4_4 _3182_ (.A(_1801_),
    .B(_1051_),
    .C(_1052_),
    .D(\count[4] ),
    .Y(_1214_));
 sky130_fd_sc_hd__o211ai_2 _3183_ (.A1(_0645_),
    .A2(_1057_),
    .B1(_1213_),
    .C1(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_2 _3184_ (.A(_1215_),
    .B(\acc[34] ),
    .Y(_1216_));
 sky130_fd_sc_hd__o2111ai_4 _3185_ (.A1(_0645_),
    .A2(_1057_),
    .B1(_1213_),
    .C1(_1214_),
    .D1(_1794_),
    .Y(_1217_));
 sky130_fd_sc_hd__nand2_1 _3186_ (.A(_1216_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__and4_1 _3187_ (.A(_1207_),
    .B(_1209_),
    .C(_1216_),
    .D(_1217_),
    .X(_1219_));
 sky130_fd_sc_hd__nand4_2 _3188_ (.A(_1207_),
    .B(_1209_),
    .C(_1216_),
    .D(_1217_),
    .Y(_1220_));
 sky130_fd_sc_hd__nand4_2 _3189_ (.A(_1801_),
    .B(_1040_),
    .C(_1041_),
    .D(\count[4] ),
    .Y(_1221_));
 sky130_fd_sc_hd__nand3_1 _3190_ (.A(_0886_),
    .B(_0887_),
    .C(\count[3] ),
    .Y(_1222_));
 sky130_fd_sc_hd__o211ai_2 _3191_ (.A1(net137),
    .A2(_0727_),
    .B1(_0878_),
    .C1(_1803_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand3_1 _3192_ (.A(_1222_),
    .B(_1223_),
    .C(_0648_),
    .Y(_1224_));
 sky130_fd_sc_hd__o211ai_4 _3193_ (.A1(_0645_),
    .A2(_1046_),
    .B1(_1221_),
    .C1(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__xnor2_2 _3194_ (.A(\acc[32] ),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__inv_2 _3195_ (.A(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__nand3_1 _3196_ (.A(_0853_),
    .B(_0854_),
    .C(net136),
    .Y(_1228_));
 sky130_fd_sc_hd__o211ai_2 _3197_ (.A1(_0719_),
    .A2(\count[2] ),
    .B1(_1803_),
    .C1(_0867_),
    .Y(_1229_));
 sky130_fd_sc_hd__nand3_1 _3198_ (.A(_1228_),
    .B(_1229_),
    .C(_0648_),
    .Y(_1230_));
 sky130_fd_sc_hd__nand3_1 _3199_ (.A(_1031_),
    .B(_0544_),
    .C(_1030_),
    .Y(_1231_));
 sky130_fd_sc_hd__o311a_2 _3200_ (.A1(_1801_),
    .A2(\count[4] ),
    .A3(_1029_),
    .B1(_1230_),
    .C1(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__nand2_1 _3201_ (.A(_1232_),
    .B(_1795_),
    .Y(_1233_));
 sky130_fd_sc_hd__xor2_2 _3202_ (.A(\acc[33] ),
    .B(_1232_),
    .X(_1234_));
 sky130_fd_sc_hd__nor2_1 _3203_ (.A(_1226_),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__nor4_1 _3204_ (.A(_1210_),
    .B(_1218_),
    .C(_1226_),
    .D(_1234_),
    .Y(_1236_));
 sky130_fd_sc_hd__and3_1 _3205_ (.A(_1202_),
    .B(_1219_),
    .C(_1235_),
    .X(_1237_));
 sky130_fd_sc_hd__nand3_1 _3206_ (.A(_1202_),
    .B(_1219_),
    .C(_1235_),
    .Y(_1238_));
 sky130_fd_sc_hd__a31o_1 _3207_ (.A1(_1163_),
    .A2(_1164_),
    .A3(_0972_),
    .B1(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__nand2_1 _3208_ (.A(_1190_),
    .B(_1198_),
    .Y(_1240_));
 sky130_fd_sc_hd__a22o_1 _3209_ (.A1(_1180_),
    .A2(\acc[36] ),
    .B1(\acc[37] ),
    .B2(_1171_),
    .X(_1241_));
 sky130_fd_sc_hd__a21o_1 _3210_ (.A1(_1174_),
    .A2(_1182_),
    .B1(_1172_),
    .X(_1242_));
 sky130_fd_sc_hd__o2bb2ai_1 _3211_ (.A1_N(_1225_),
    .A2_N(\acc[32] ),
    .B1(_1795_),
    .B2(_1232_),
    .Y(_1243_));
 sky130_fd_sc_hd__nand2_1 _3212_ (.A(_1233_),
    .B(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__o221ai_4 _3213_ (.A1(_1208_),
    .A2(_1216_),
    .B1(_1220_),
    .B2(_1244_),
    .C1(_1207_),
    .Y(_1245_));
 sky130_fd_sc_hd__o2bb2ai_1 _3214_ (.A1_N(_1199_),
    .A2_N(_1240_),
    .B1(_1242_),
    .B2(_1201_),
    .Y(_1246_));
 sky130_fd_sc_hd__a21oi_2 _3215_ (.A1(_1245_),
    .A2(_1202_),
    .B1(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__o21ai_1 _3216_ (.A1(_0924_),
    .A2(_1247_),
    .B1(_0914_),
    .Y(_1248_));
 sky130_fd_sc_hd__nor2_1 _3217_ (.A(_0924_),
    .B(_1238_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand3_1 _3218_ (.A(_0923_),
    .B(_1202_),
    .C(_1236_),
    .Y(_1250_));
 sky130_fd_sc_hd__a31oi_1 _3219_ (.A1(_1163_),
    .A2(_1164_),
    .A3(_0972_),
    .B1(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__a21o_1 _3220_ (.A1(_1165_),
    .A2(_1249_),
    .B1(_1248_),
    .X(_1252_));
 sky130_fd_sc_hd__a21oi_1 _3221_ (.A1(_1165_),
    .A2(_1249_),
    .B1(_1248_),
    .Y(_1253_));
 sky130_fd_sc_hd__o211a_1 _3222_ (.A1(net136),
    .A2(_0787_),
    .B1(_1205_),
    .C1(_0544_),
    .X(_1254_));
 sky130_fd_sc_hd__a31o_1 _3223_ (.A1(_1066_),
    .A2(_1070_),
    .A3(net135),
    .B1(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__nor2_1 _3224_ (.A(\acc[51] ),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__a311o_1 _3225_ (.A1(_1066_),
    .A2(_1070_),
    .A3(net135),
    .B1(_1254_),
    .C1(\acc[51] ),
    .X(_1257_));
 sky130_fd_sc_hd__nand2_1 _3226_ (.A(_1255_),
    .B(\acc[51] ),
    .Y(_1258_));
 sky130_fd_sc_hd__nand2_1 _3227_ (.A(_1257_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__and3_1 _3228_ (.A(_1211_),
    .B(_1212_),
    .C(_0544_),
    .X(_1260_));
 sky130_fd_sc_hd__and3_1 _3229_ (.A(_1055_),
    .B(_1058_),
    .C(net135),
    .X(_1261_));
 sky130_fd_sc_hd__o21ai_2 _3230_ (.A1(_1260_),
    .A2(_1261_),
    .B1(\acc[50] ),
    .Y(_1262_));
 sky130_fd_sc_hd__a311o_1 _3231_ (.A1(net135),
    .A2(_1055_),
    .A3(_1058_),
    .B1(_1260_),
    .C1(\acc[50] ),
    .X(_1263_));
 sky130_fd_sc_hd__nand2_1 _3232_ (.A(_1262_),
    .B(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__and4_1 _3233_ (.A(_1257_),
    .B(_1258_),
    .C(_1262_),
    .D(_1263_),
    .X(_1265_));
 sky130_fd_sc_hd__o211ai_2 _3234_ (.A1(_1802_),
    .A2(_1028_),
    .B1(net135),
    .C1(_1034_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand4_2 _3235_ (.A(_1801_),
    .B(_1228_),
    .C(_1229_),
    .D(\count[4] ),
    .Y(_1267_));
 sky130_fd_sc_hd__a21boi_2 _3236_ (.A1(_1266_),
    .A2(_1267_),
    .B1_N(\acc[49] ),
    .Y(_1268_));
 sky130_fd_sc_hd__nand3b_1 _3237_ (.A_N(\acc[49] ),
    .B(_1266_),
    .C(_1267_),
    .Y(_1269_));
 sky130_fd_sc_hd__and2b_1 _3238_ (.A_N(_1268_),
    .B(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__o21a_1 _3239_ (.A1(_1802_),
    .A2(_1045_),
    .B1(net135),
    .X(_1271_));
 sky130_fd_sc_hd__a32o_1 _3240_ (.A1(_0544_),
    .A2(_1222_),
    .A3(_1223_),
    .B1(_1044_),
    .B2(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__and2_1 _3241_ (.A(_1272_),
    .B(\acc[48] ),
    .X(_1273_));
 sky130_fd_sc_hd__xnor2_1 _3242_ (.A(\acc[48] ),
    .B(_1272_),
    .Y(_1274_));
 sky130_fd_sc_hd__nor3b_2 _3243_ (.A(_1268_),
    .B(_1274_),
    .C_N(_1269_),
    .Y(_1275_));
 sky130_fd_sc_hd__and4_1 _3244_ (.A(_0525_),
    .B(_0534_),
    .C(_0544_),
    .D(net136),
    .X(_1276_));
 sky130_fd_sc_hd__a31o_1 _3245_ (.A1(_0992_),
    .A2(net135),
    .A3(_0989_),
    .B1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__nand2_1 _3246_ (.A(_1277_),
    .B(\acc[55] ),
    .Y(_1278_));
 sky130_fd_sc_hd__a311o_1 _3247_ (.A1(_0992_),
    .A2(net135),
    .A3(_0989_),
    .B1(_1276_),
    .C1(\acc[55] ),
    .X(_1279_));
 sky130_fd_sc_hd__nand2_1 _3248_ (.A(_1278_),
    .B(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__a32oi_4 _3249_ (.A1(_0982_),
    .A2(net135),
    .A3(_0979_),
    .B1(_1188_),
    .B2(_0544_),
    .Y(_1281_));
 sky130_fd_sc_hd__nand2b_1 _3250_ (.A_N(_1281_),
    .B(\acc[54] ),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2b_1 _3251_ (.A_N(\acc[54] ),
    .B(_1281_),
    .Y(_1283_));
 sky130_fd_sc_hd__nand2_1 _3252_ (.A(_1282_),
    .B(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__inv_2 _3253_ (.A(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__nand4_1 _3254_ (.A(_1801_),
    .B(_1167_),
    .C(\count[4] ),
    .D(_1166_),
    .Y(_1286_));
 sky130_fd_sc_hd__o211ai_2 _3255_ (.A1(_1802_),
    .A2(_1014_),
    .B1(net135),
    .C1(_1020_),
    .Y(_1287_));
 sky130_fd_sc_hd__a21boi_1 _3256_ (.A1(_1286_),
    .A2(_1287_),
    .B1_N(\acc[53] ),
    .Y(_1288_));
 sky130_fd_sc_hd__and3b_1 _3257_ (.A_N(\acc[53] ),
    .B(_1286_),
    .C(_1287_),
    .X(_1289_));
 sky130_fd_sc_hd__nor2_1 _3258_ (.A(_1288_),
    .B(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__or2_1 _3259_ (.A(_1288_),
    .B(_1289_),
    .X(_1291_));
 sky130_fd_sc_hd__o32ai_4 _3260_ (.A1(_0545_),
    .A2(_1175_),
    .A3(_1176_),
    .B1(_1007_),
    .B2(_1801_),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _3261_ (.A(_1292_),
    .B(\acc[52] ),
    .Y(_1293_));
 sky130_fd_sc_hd__xnor2_2 _3262_ (.A(\acc[52] ),
    .B(_1292_),
    .Y(_1294_));
 sky130_fd_sc_hd__or3_1 _3263_ (.A(_1288_),
    .B(_1289_),
    .C(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__nor4_1 _3264_ (.A(_1280_),
    .B(_1284_),
    .C(_1291_),
    .D(_1294_),
    .Y(_1296_));
 sky130_fd_sc_hd__and3_1 _3265_ (.A(_1265_),
    .B(_1275_),
    .C(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__nand3_1 _3266_ (.A(_1265_),
    .B(_1275_),
    .C(_1296_),
    .Y(_1298_));
 sky130_fd_sc_hd__o21bai_1 _3267_ (.A1(_1248_),
    .A2(_1251_),
    .B1_N(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__a21oi_1 _3268_ (.A1(_1273_),
    .A2(_1269_),
    .B1(_1268_),
    .Y(_1300_));
 sky130_fd_sc_hd__o21a_1 _3269_ (.A1(_1256_),
    .A2(_1262_),
    .B1(_1258_),
    .X(_1301_));
 sky130_fd_sc_hd__o31ai_2 _3270_ (.A1(_1259_),
    .A2(_1264_),
    .A3(_1300_),
    .B1(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__o21ba_1 _3271_ (.A1(_1293_),
    .A2(_1289_),
    .B1_N(_1288_),
    .X(_1303_));
 sky130_fd_sc_hd__and4bb_1 _3272_ (.A_N(_1284_),
    .B_N(_1303_),
    .C(_1278_),
    .D(_1279_),
    .X(_1304_));
 sky130_fd_sc_hd__and3b_1 _3273_ (.A_N(_1281_),
    .B(\acc[54] ),
    .C(_1279_),
    .X(_1305_));
 sky130_fd_sc_hd__a21o_1 _3274_ (.A1(\acc[55] ),
    .A2(_1277_),
    .B1(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__a211oi_1 _3275_ (.A1(_1296_),
    .A2(_1302_),
    .B1(_1306_),
    .C1(_1304_),
    .Y(_1307_));
 sky130_fd_sc_hd__a211o_1 _3276_ (.A1(_1296_),
    .A2(_1302_),
    .B1(_1306_),
    .C1(_1304_),
    .X(_1308_));
 sky130_fd_sc_hd__a21oi_2 _3277_ (.A1(_1252_),
    .A2(_1297_),
    .B1(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__o2111a_1 _3278_ (.A1(\count[2] ),
    .A2(_0728_),
    .B1(_0877_),
    .C1(_0544_),
    .D1(net136),
    .X(_1310_));
 sky130_fd_sc_hd__a31o_1 _3279_ (.A1(_0965_),
    .A2(_0966_),
    .A3(net135),
    .B1(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__nand2_2 _3280_ (.A(_1311_),
    .B(\acc[56] ),
    .Y(_1312_));
 sky130_fd_sc_hd__a311o_1 _3281_ (.A1(_0965_),
    .A2(_0966_),
    .A3(net135),
    .B1(_1310_),
    .C1(\acc[56] ),
    .X(_1313_));
 sky130_fd_sc_hd__nand2_2 _3282_ (.A(_1312_),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__a32o_1 _3283_ (.A1(_0962_),
    .A2(_0963_),
    .A3(net135),
    .B1(_0544_),
    .B2(_0869_),
    .X(_1315_));
 sky130_fd_sc_hd__nor2_1 _3284_ (.A(\acc[57] ),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2_1 _3285_ (.A(_1315_),
    .B(\acc[57] ),
    .Y(_1317_));
 sky130_fd_sc_hd__nand2b_1 _3286_ (.A_N(_1316_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__and3_1 _3287_ (.A(_0836_),
    .B(_0544_),
    .C(net136),
    .X(_1319_));
 sky130_fd_sc_hd__a31o_1 _3288_ (.A1(net135),
    .A2(_0953_),
    .A3(_0954_),
    .B1(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__nand2_1 _3289_ (.A(_1320_),
    .B(\acc[58] ),
    .Y(_1321_));
 sky130_fd_sc_hd__xor2_1 _3290_ (.A(\acc[58] ),
    .B(_1320_),
    .X(_1322_));
 sky130_fd_sc_hd__xnor2_1 _3291_ (.A(\acc[58] ),
    .B(_1320_),
    .Y(_1323_));
 sky130_fd_sc_hd__a32o_1 _3292_ (.A1(net136),
    .A2(_0544_),
    .A3(_0787_),
    .B1(_0949_),
    .B2(net135),
    .X(_1324_));
 sky130_fd_sc_hd__nor2_1 _3293_ (.A(\acc[59] ),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _3294_ (.A(_1324_),
    .B(\acc[59] ),
    .Y(_1326_));
 sky130_fd_sc_hd__nand2b_1 _3295_ (.A_N(_1325_),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__or4_1 _3296_ (.A(_1314_),
    .B(_1318_),
    .C(_1323_),
    .D(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__a21oi_1 _3297_ (.A1(_1299_),
    .A2(_1307_),
    .B1(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__a2111o_1 _3298_ (.A1(_1312_),
    .A2(_1317_),
    .B1(_1323_),
    .C1(_1316_),
    .D1(_1327_),
    .X(_1330_));
 sky130_fd_sc_hd__a21o_1 _3299_ (.A1(_1321_),
    .A2(_1326_),
    .B1(_1325_),
    .X(_1331_));
 sky130_fd_sc_hd__nand2_1 _3300_ (.A(_1330_),
    .B(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__and3_1 _3301_ (.A(_0728_),
    .B(_0548_),
    .C(_0544_),
    .X(_1333_));
 sky130_fd_sc_hd__a31o_1 _3302_ (.A1(_0926_),
    .A2(_0927_),
    .A3(net135),
    .B1(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__nand2_1 _3303_ (.A(_1334_),
    .B(\acc[60] ),
    .Y(_1335_));
 sky130_fd_sc_hd__xor2_1 _3304_ (.A(\acc[60] ),
    .B(_1334_),
    .X(_1336_));
 sky130_fd_sc_hd__a32o_1 _3305_ (.A1(_0930_),
    .A2(net135),
    .A3(_0929_),
    .B1(_0544_),
    .B2(_0720_),
    .X(_1337_));
 sky130_fd_sc_hd__nor2_1 _3306_ (.A(\acc[61] ),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _3307_ (.A(_1337_),
    .B(\acc[61] ),
    .Y(_1339_));
 sky130_fd_sc_hd__and2b_1 _3308_ (.A_N(_1338_),
    .B(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__inv_2 _3309_ (.A(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _3310_ (.A(_1336_),
    .B(_1340_),
    .Y(_1342_));
 sky130_fd_sc_hd__o21bai_1 _3311_ (.A1(_1332_),
    .A2(_1329_),
    .B1_N(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__o21a_1 _3312_ (.A1(_1335_),
    .A2(_1338_),
    .B1(_1339_),
    .X(_1344_));
 sky130_fd_sc_hd__nor2_1 _3313_ (.A(\acc[62] ),
    .B(_0640_),
    .Y(_1345_));
 sky130_fd_sc_hd__or2_1 _3314_ (.A(\acc[62] ),
    .B(_0640_),
    .X(_1346_));
 sky130_fd_sc_hd__and2_1 _3315_ (.A(\acc[62] ),
    .B(_0640_),
    .X(_1347_));
 sky130_fd_sc_hd__nand2_1 _3316_ (.A(\acc[62] ),
    .B(_0640_),
    .Y(_1348_));
 sky130_fd_sc_hd__a22oi_1 _3317_ (.A1(_1346_),
    .A2(_1348_),
    .B1(_1343_),
    .B2(_1344_),
    .Y(_1349_));
 sky130_fd_sc_hd__o2bb2ai_1 _3318_ (.A1_N(_1344_),
    .A2_N(_1343_),
    .B1(_1347_),
    .B2(_1345_),
    .Y(_1350_));
 sky130_fd_sc_hd__o22ai_1 _3319_ (.A1(_0541_),
    .A2(_0542_),
    .B1(_0642_),
    .B2(_1349_),
    .Y(_1351_));
 sky130_fd_sc_hd__nand3_1 _3320_ (.A(_1350_),
    .B(_0543_),
    .C(_0643_),
    .Y(_1352_));
 sky130_fd_sc_hd__and3_4 _3321_ (.A(\m[0] ),
    .B(_1922_),
    .C(_1801_),
    .X(_1353_));
 sky130_fd_sc_hd__or3b_4 _3322_ (.A(net135),
    .B(_1923_),
    .C_N(\m[0] ),
    .X(_1354_));
 sky130_fd_sc_hd__a31o_1 _3323_ (.A1(_1351_),
    .A2(_1352_),
    .A3(_1353_),
    .B1(_0438_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _3324_ (.A(net133),
    .B(\acc[62] ),
    .Y(_1355_));
 sky130_fd_sc_hd__and4_1 _3325_ (.A(_1343_),
    .B(_1344_),
    .C(_1346_),
    .D(_1348_),
    .X(_1356_));
 sky130_fd_sc_hd__o31ai_1 _3326_ (.A1(_1349_),
    .A2(_1354_),
    .A3(_1356_),
    .B1(_1355_),
    .Y(_0338_));
 sky130_fd_sc_hd__o21ai_1 _3327_ (.A1(_1332_),
    .A2(_1329_),
    .B1(_1336_),
    .Y(_1357_));
 sky130_fd_sc_hd__a21oi_1 _3328_ (.A1(_1335_),
    .A2(_1357_),
    .B1(_1341_),
    .Y(_1358_));
 sky130_fd_sc_hd__a31o_1 _3329_ (.A1(_1335_),
    .A2(_1341_),
    .A3(_1357_),
    .B1(_1354_),
    .X(_1359_));
 sky130_fd_sc_hd__o2bb2ai_1 _3330_ (.A1_N(\acc[61] ),
    .A2_N(net133),
    .B1(_1358_),
    .B2(_1359_),
    .Y(_0337_));
 sky130_fd_sc_hd__o311a_1 _3331_ (.A1(_1332_),
    .A2(_1336_),
    .A3(_1329_),
    .B1(_1353_),
    .C1(_1357_),
    .X(_1360_));
 sky130_fd_sc_hd__a21o_1 _3332_ (.A1(\acc[60] ),
    .A2(net133),
    .B1(_1360_),
    .X(_0336_));
 sky130_fd_sc_hd__o211ai_2 _3333_ (.A1(_1314_),
    .A2(_1309_),
    .B1(_1312_),
    .C1(_1317_),
    .Y(_1361_));
 sky130_fd_sc_hd__o21ai_1 _3334_ (.A1(\acc[57] ),
    .A2(_1315_),
    .B1(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__o211ai_2 _3335_ (.A1(\acc[57] ),
    .A2(_1315_),
    .B1(_1322_),
    .C1(_1361_),
    .Y(_1363_));
 sky130_fd_sc_hd__a21oi_1 _3336_ (.A1(_1321_),
    .A2(_1363_),
    .B1(_1327_),
    .Y(_1364_));
 sky130_fd_sc_hd__a31o_1 _3337_ (.A1(_1321_),
    .A2(_1327_),
    .A3(_1363_),
    .B1(_1354_),
    .X(_1365_));
 sky130_fd_sc_hd__o2bb2ai_1 _3338_ (.A1_N(\acc[59] ),
    .A2_N(net133),
    .B1(_1364_),
    .B2(_1365_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _3339_ (.A(_1323_),
    .B(_1362_),
    .Y(_1366_));
 sky130_fd_sc_hd__a32o_1 _3340_ (.A1(_1366_),
    .A2(_1353_),
    .A3(_1363_),
    .B1(net133),
    .B2(\acc[58] ),
    .X(_0334_));
 sky130_fd_sc_hd__o21ai_1 _3341_ (.A1(_1314_),
    .A2(_1309_),
    .B1(_1312_),
    .Y(_1367_));
 sky130_fd_sc_hd__o211ai_1 _3342_ (.A1(_1314_),
    .A2(_1309_),
    .B1(_1312_),
    .C1(_1318_),
    .Y(_1368_));
 sky130_fd_sc_hd__nand3b_1 _3343_ (.A_N(_1316_),
    .B(_1317_),
    .C(_1367_),
    .Y(_1369_));
 sky130_fd_sc_hd__a32o_1 _3344_ (.A1(_1368_),
    .A2(_1369_),
    .A3(_1353_),
    .B1(net133),
    .B2(\acc[57] ),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _3345_ (.A(_1309_),
    .B(_1314_),
    .Y(_1370_));
 sky130_fd_sc_hd__o211a_1 _3346_ (.A1(_1314_),
    .A2(_1309_),
    .B1(_1924_),
    .C1(\m[0] ),
    .X(_1371_));
 sky130_fd_sc_hd__a22o_1 _3347_ (.A1(\acc[56] ),
    .A2(net133),
    .B1(_1371_),
    .B2(_1370_),
    .X(_0332_));
 sky130_fd_sc_hd__nor2_1 _3348_ (.A(_1253_),
    .B(_1274_),
    .Y(_1372_));
 sky130_fd_sc_hd__a221oi_2 _3349_ (.A1(_1273_),
    .A2(_1269_),
    .B1(_1252_),
    .B2(_1275_),
    .C1(_1268_),
    .Y(_1373_));
 sky130_fd_sc_hd__a31oi_2 _3350_ (.A1(_1252_),
    .A2(_1265_),
    .A3(_1275_),
    .B1(_1302_),
    .Y(_1374_));
 sky130_fd_sc_hd__o21ai_1 _3351_ (.A1(_1295_),
    .A2(_1374_),
    .B1(_1303_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_1 _3352_ (.A(_1375_),
    .B(_1285_),
    .Y(_1376_));
 sky130_fd_sc_hd__a21oi_1 _3353_ (.A1(_1282_),
    .A2(_1376_),
    .B1(_1280_),
    .Y(_1377_));
 sky130_fd_sc_hd__a31o_1 _3354_ (.A1(_1280_),
    .A2(_1282_),
    .A3(_1376_),
    .B1(_1354_),
    .X(_1378_));
 sky130_fd_sc_hd__o2bb2ai_1 _3355_ (.A1_N(\acc[55] ),
    .A2_N(net133),
    .B1(_1377_),
    .B2(_1378_),
    .Y(_0331_));
 sky130_fd_sc_hd__or2_1 _3356_ (.A(_1285_),
    .B(_1375_),
    .X(_1379_));
 sky130_fd_sc_hd__a32o_1 _3357_ (.A1(_1379_),
    .A2(_1353_),
    .A3(_1376_),
    .B1(net133),
    .B2(\acc[54] ),
    .X(_0330_));
 sky130_fd_sc_hd__or2_1 _3358_ (.A(_1294_),
    .B(_1374_),
    .X(_1380_));
 sky130_fd_sc_hd__o21ai_1 _3359_ (.A1(_1294_),
    .A2(_1374_),
    .B1(_1293_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _3360_ (.A(_1381_),
    .B(_1290_),
    .Y(_1382_));
 sky130_fd_sc_hd__or2_1 _3361_ (.A(_1290_),
    .B(_1381_),
    .X(_1383_));
 sky130_fd_sc_hd__a32o_1 _3362_ (.A1(_1383_),
    .A2(_1353_),
    .A3(_1382_),
    .B1(net133),
    .B2(\acc[53] ),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _3363_ (.A(_1374_),
    .B(_1294_),
    .Y(_1384_));
 sky130_fd_sc_hd__a32o_1 _3364_ (.A1(_1380_),
    .A2(_1384_),
    .A3(_1353_),
    .B1(net133),
    .B2(\acc[52] ),
    .X(_0328_));
 sky130_fd_sc_hd__o21a_1 _3365_ (.A1(_1264_),
    .A2(_1373_),
    .B1(_1262_),
    .X(_1385_));
 sky130_fd_sc_hd__o211a_1 _3366_ (.A1(_1264_),
    .A2(_1373_),
    .B1(_1259_),
    .C1(_1262_),
    .X(_1386_));
 sky130_fd_sc_hd__o21ai_1 _3367_ (.A1(_1259_),
    .A2(_1385_),
    .B1(_1353_),
    .Y(_1387_));
 sky130_fd_sc_hd__a2bb2o_1 _3368_ (.A1_N(_1386_),
    .A2_N(_1387_),
    .B1(\acc[51] ),
    .B2(net133),
    .X(_0327_));
 sky130_fd_sc_hd__nand2_1 _3369_ (.A(_1373_),
    .B(_1264_),
    .Y(_1388_));
 sky130_fd_sc_hd__o211a_1 _3370_ (.A1(_1264_),
    .A2(_1373_),
    .B1(\m[0] ),
    .C1(_1924_),
    .X(_1389_));
 sky130_fd_sc_hd__a22o_1 _3371_ (.A1(\acc[50] ),
    .A2(net133),
    .B1(_1389_),
    .B2(_1388_),
    .X(_0326_));
 sky130_fd_sc_hd__o21ai_1 _3372_ (.A1(_1273_),
    .A2(_1372_),
    .B1(_1270_),
    .Y(_1390_));
 sky130_fd_sc_hd__or3_1 _3373_ (.A(_1270_),
    .B(_1273_),
    .C(_1372_),
    .X(_1391_));
 sky130_fd_sc_hd__a32o_1 _3374_ (.A1(_1391_),
    .A2(_1353_),
    .A3(_1390_),
    .B1(net133),
    .B2(\acc[49] ),
    .X(_0325_));
 sky130_fd_sc_hd__a21o_1 _3375_ (.A1(_1253_),
    .A2(_1274_),
    .B1(_1354_),
    .X(_1392_));
 sky130_fd_sc_hd__a2bb2o_1 _3376_ (.A1_N(_1372_),
    .A2_N(_1392_),
    .B1(\acc[48] ),
    .B2(net133),
    .X(_0324_));
 sky130_fd_sc_hd__a21boi_2 _3377_ (.A1(_1165_),
    .A2(_1237_),
    .B1_N(_1247_),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2_1 _3378_ (.A(_1239_),
    .B(_1247_),
    .Y(_1394_));
 sky130_fd_sc_hd__o21bai_1 _3379_ (.A1(_0922_),
    .A2(_1393_),
    .B1_N(_0906_),
    .Y(_1395_));
 sky130_fd_sc_hd__nand2_1 _3380_ (.A(_1395_),
    .B(_0910_),
    .Y(_1396_));
 sky130_fd_sc_hd__nand3_1 _3381_ (.A(_0725_),
    .B(_1395_),
    .C(_0910_),
    .Y(_1397_));
 sky130_fd_sc_hd__a21oi_1 _3382_ (.A1(_1397_),
    .A2(_0786_),
    .B1(_0662_),
    .Y(_1398_));
 sky130_fd_sc_hd__o211ai_1 _3383_ (.A1(_0657_),
    .A2(_1398_),
    .B1(_0658_),
    .C1(_0650_),
    .Y(_1399_));
 sky130_fd_sc_hd__a32o_1 _3384_ (.A1(\acc[46] ),
    .A2(_0655_),
    .A3(_0654_),
    .B1(_0650_),
    .B2(_0658_),
    .X(_1400_));
 sky130_fd_sc_hd__o211a_1 _3385_ (.A1(_1400_),
    .A2(_1398_),
    .B1(_1924_),
    .C1(\m[0] ),
    .X(_1401_));
 sky130_fd_sc_hd__a22o_1 _3386_ (.A1(\acc[47] ),
    .A2(net132),
    .B1(_1401_),
    .B2(_1399_),
    .X(_0323_));
 sky130_fd_sc_hd__a311oi_1 _3387_ (.A1(_0662_),
    .A2(_0786_),
    .A3(_1397_),
    .B1(_1354_),
    .C1(_1398_),
    .Y(_1402_));
 sky130_fd_sc_hd__a21o_1 _3388_ (.A1(\acc[46] ),
    .A2(net132),
    .B1(_1402_),
    .X(_0322_));
 sky130_fd_sc_hd__a221o_1 _3389_ (.A1(_0724_),
    .A2(_0725_),
    .B1(_1395_),
    .B2(_0910_),
    .C1(_0784_),
    .X(_1403_));
 sky130_fd_sc_hd__a21o_1 _3390_ (.A1(_0785_),
    .A2(_1396_),
    .B1(_0908_),
    .X(_1404_));
 sky130_fd_sc_hd__a32o_1 _3391_ (.A1(_1404_),
    .A2(_1353_),
    .A3(_1403_),
    .B1(net132),
    .B2(\acc[45] ),
    .X(_0321_));
 sky130_fd_sc_hd__a311o_1 _3392_ (.A1(_1394_),
    .A2(_0921_),
    .A3(_0846_),
    .B1(_0910_),
    .C1(_0906_),
    .X(_1405_));
 sky130_fd_sc_hd__a32o_1 _3393_ (.A1(_1405_),
    .A2(_1353_),
    .A3(_1396_),
    .B1(net132),
    .B2(\acc[44] ),
    .X(_0320_));
 sky130_fd_sc_hd__o32a_1 _3394_ (.A1(_1789_),
    .A2(_0899_),
    .A3(_0901_),
    .B1(_0920_),
    .B2(_1393_),
    .X(_1406_));
 sky130_fd_sc_hd__a211o_1 _3395_ (.A1(_1406_),
    .A2(_0874_),
    .B1(_0845_),
    .C1(_0875_),
    .X(_1407_));
 sky130_fd_sc_hd__a21oi_1 _3396_ (.A1(_0843_),
    .A2(_1407_),
    .B1(_0813_),
    .Y(_1408_));
 sky130_fd_sc_hd__a31o_1 _3397_ (.A1(_0813_),
    .A2(_0843_),
    .A3(_1407_),
    .B1(_1354_),
    .X(_1409_));
 sky130_fd_sc_hd__o2bb2ai_1 _3398_ (.A1_N(\acc[43] ),
    .A2_N(net132),
    .B1(_1408_),
    .B2(_1409_),
    .Y(_0319_));
 sky130_fd_sc_hd__o311ai_1 _3399_ (.A1(_0875_),
    .A2(_0920_),
    .A3(_1393_),
    .B1(_0905_),
    .C1(_0845_),
    .Y(_1410_));
 sky130_fd_sc_hd__a32o_1 _3400_ (.A1(_1407_),
    .A2(_1410_),
    .A3(_1353_),
    .B1(net132),
    .B2(\acc[42] ),
    .X(_0318_));
 sky130_fd_sc_hd__a221o_1 _3401_ (.A1(\acc[40] ),
    .A2(_0902_),
    .B1(_1394_),
    .B2(_0919_),
    .C1(_0915_),
    .X(_1411_));
 sky130_fd_sc_hd__or3_1 _3402_ (.A(_0873_),
    .B(_0875_),
    .C(_1406_),
    .X(_1412_));
 sky130_fd_sc_hd__a32o_1 _3403_ (.A1(_1412_),
    .A2(_1353_),
    .A3(_1411_),
    .B1(net132),
    .B2(\acc[41] ),
    .X(_0317_));
 sky130_fd_sc_hd__and3_1 _3404_ (.A(_0920_),
    .B(_1239_),
    .C(_1247_),
    .X(_1413_));
 sky130_fd_sc_hd__o21ai_1 _3405_ (.A1(_0920_),
    .A2(_1393_),
    .B1(_1353_),
    .Y(_1414_));
 sky130_fd_sc_hd__a2bb2o_1 _3406_ (.A1_N(_1413_),
    .A2_N(_1414_),
    .B1(\acc[40] ),
    .B2(net132),
    .X(_0316_));
 sky130_fd_sc_hd__a21oi_1 _3407_ (.A1(_1165_),
    .A2(_1236_),
    .B1(_1245_),
    .Y(_1415_));
 sky130_fd_sc_hd__nor2_1 _3408_ (.A(_1184_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__o211a_1 _3409_ (.A1(_1184_),
    .A2(_1415_),
    .B1(_1174_),
    .C1(_1182_),
    .X(_1417_));
 sky130_fd_sc_hd__o221ai_4 _3410_ (.A1(\acc[37] ),
    .A2(_1171_),
    .B1(_1241_),
    .B2(_1416_),
    .C1(_1193_),
    .Y(_1418_));
 sky130_fd_sc_hd__a21oi_1 _3411_ (.A1(_1190_),
    .A2(_1418_),
    .B1(_1200_),
    .Y(_1419_));
 sky130_fd_sc_hd__a31o_1 _3412_ (.A1(_1190_),
    .A2(_1200_),
    .A3(_1418_),
    .B1(_1354_),
    .X(_1420_));
 sky130_fd_sc_hd__a2bb2o_1 _3413_ (.A1_N(_1419_),
    .A2_N(_1420_),
    .B1(\acc[39] ),
    .B2(net132),
    .X(_0315_));
 sky130_fd_sc_hd__o21ai_1 _3414_ (.A1(_1172_),
    .A2(_1417_),
    .B1(_1192_),
    .Y(_1421_));
 sky130_fd_sc_hd__a32o_1 _3415_ (.A1(_1421_),
    .A2(_1353_),
    .A3(_1418_),
    .B1(net132),
    .B2(\acc[38] ),
    .X(_0314_));
 sky130_fd_sc_hd__a221o_1 _3416_ (.A1(_1173_),
    .A2(_1174_),
    .B1(_1180_),
    .B2(\acc[36] ),
    .C1(_1416_),
    .X(_1422_));
 sky130_fd_sc_hd__o211ai_1 _3417_ (.A1(_1181_),
    .A2(_1416_),
    .B1(_1173_),
    .C1(_1174_),
    .Y(_1423_));
 sky130_fd_sc_hd__a32o_1 _3418_ (.A1(_1423_),
    .A2(_1353_),
    .A3(_1422_),
    .B1(net132),
    .B2(\acc[37] ),
    .X(_0313_));
 sky130_fd_sc_hd__a221o_1 _3419_ (.A1(_1182_),
    .A2(_1183_),
    .B1(_1165_),
    .B2(_1236_),
    .C1(_1245_),
    .X(_1424_));
 sky130_fd_sc_hd__o211a_1 _3420_ (.A1(_1184_),
    .A2(_1415_),
    .B1(\m[0] ),
    .C1(_1924_),
    .X(_1425_));
 sky130_fd_sc_hd__a22o_1 _3421_ (.A1(\acc[36] ),
    .A2(net132),
    .B1(_1425_),
    .B2(_1424_),
    .X(_0312_));
 sky130_fd_sc_hd__a31o_1 _3422_ (.A1(_1163_),
    .A2(_1164_),
    .A3(_0972_),
    .B1(_1226_),
    .X(_1426_));
 sky130_fd_sc_hd__a311o_1 _3423_ (.A1(_1163_),
    .A2(_1164_),
    .A3(_0972_),
    .B1(_1226_),
    .C1(_1234_),
    .X(_1427_));
 sky130_fd_sc_hd__a21oi_1 _3424_ (.A1(_1244_),
    .A2(_1427_),
    .B1(_1218_),
    .Y(_1428_));
 sky130_fd_sc_hd__inv_2 _3425_ (.A(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__a21o_1 _3426_ (.A1(_1216_),
    .A2(_1429_),
    .B1(_1210_),
    .X(_1430_));
 sky130_fd_sc_hd__a221o_1 _3427_ (.A1(_1207_),
    .A2(_1209_),
    .B1(_1215_),
    .B2(\acc[34] ),
    .C1(_1428_),
    .X(_1431_));
 sky130_fd_sc_hd__a32o_1 _3428_ (.A1(_1430_),
    .A2(_1431_),
    .A3(_1353_),
    .B1(net133),
    .B2(\acc[35] ),
    .X(_0311_));
 sky130_fd_sc_hd__nand3_1 _3429_ (.A(_1218_),
    .B(_1244_),
    .C(_1427_),
    .Y(_1432_));
 sky130_fd_sc_hd__a32o_1 _3430_ (.A1(_1429_),
    .A2(_1432_),
    .A3(_1353_),
    .B1(net133),
    .B2(\acc[34] ),
    .X(_0310_));
 sky130_fd_sc_hd__a22oi_1 _3431_ (.A1(\acc[32] ),
    .A2(_1225_),
    .B1(_1165_),
    .B2(_1227_),
    .Y(_1433_));
 sky130_fd_sc_hd__nand2_1 _3432_ (.A(_1433_),
    .B(_1234_),
    .Y(_1434_));
 sky130_fd_sc_hd__o211a_1 _3433_ (.A1(_1234_),
    .A2(_1433_),
    .B1(\m[0] ),
    .C1(_1924_),
    .X(_1435_));
 sky130_fd_sc_hd__a22o_1 _3434_ (.A1(\acc[33] ),
    .A2(net133),
    .B1(_1435_),
    .B2(_1434_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _3435_ (.A(_1227_),
    .B(_1165_),
    .X(_1436_));
 sky130_fd_sc_hd__a32o_1 _3436_ (.A1(_1436_),
    .A2(_1353_),
    .A3(_1426_),
    .B1(net133),
    .B2(\acc[32] ),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_1 _3437_ (.A(_0974_),
    .B(_1162_),
    .Y(_1437_));
 sky130_fd_sc_hd__o21bai_1 _3438_ (.A1(_0974_),
    .A2(_1162_),
    .B1_N(_0969_),
    .Y(_1438_));
 sky130_fd_sc_hd__nand3_1 _3439_ (.A(_1438_),
    .B(_0960_),
    .C(_0964_),
    .Y(_1439_));
 sky130_fd_sc_hd__a21oi_1 _3440_ (.A1(_1439_),
    .A2(_0957_),
    .B1(_0942_),
    .Y(_1440_));
 sky130_fd_sc_hd__a21o_1 _3441_ (.A1(_1439_),
    .A2(_0957_),
    .B1(_0942_),
    .X(_1441_));
 sky130_fd_sc_hd__a41o_1 _3442_ (.A1(\acc[28] ),
    .A2(_1801_),
    .A3(_0926_),
    .A4(_0927_),
    .B1(_1440_),
    .X(_1442_));
 sky130_fd_sc_hd__o21ai_1 _3443_ (.A1(_0932_),
    .A2(_1440_),
    .B1(_0934_),
    .Y(_1443_));
 sky130_fd_sc_hd__o2111ai_1 _3444_ (.A1(_0932_),
    .A2(_1440_),
    .B1(_0936_),
    .C1(_0934_),
    .D1(_0933_),
    .Y(_1444_));
 sky130_fd_sc_hd__a21o_1 _3445_ (.A1(_0936_),
    .A2(_1444_),
    .B1(_0939_),
    .X(_1445_));
 sky130_fd_sc_hd__o211ai_1 _3446_ (.A1(_0940_),
    .A2(_1443_),
    .B1(_0936_),
    .C1(_0939_),
    .Y(_1446_));
 sky130_fd_sc_hd__a32o_1 _3447_ (.A1(_1445_),
    .A2(_1446_),
    .A3(_1353_),
    .B1(_0437_),
    .B2(\acc[31] ),
    .X(_0307_));
 sky130_fd_sc_hd__o21ai_1 _3448_ (.A1(_0940_),
    .A2(_1443_),
    .B1(_1353_),
    .Y(_1447_));
 sky130_fd_sc_hd__a21oi_1 _3449_ (.A1(_0940_),
    .A2(_1443_),
    .B1(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__a21o_1 _3450_ (.A1(\acc[30] ),
    .A2(_0437_),
    .B1(_1448_),
    .X(_0306_));
 sky130_fd_sc_hd__nand3_1 _3451_ (.A(_0931_),
    .B(_0934_),
    .C(_1442_),
    .Y(_1449_));
 sky130_fd_sc_hd__a21o_1 _3452_ (.A1(_0931_),
    .A2(_0934_),
    .B1(_1442_),
    .X(_1450_));
 sky130_fd_sc_hd__a32o_1 _3453_ (.A1(_1450_),
    .A2(_1353_),
    .A3(_1449_),
    .B1(_0437_),
    .B2(\acc[29] ),
    .X(_0305_));
 sky130_fd_sc_hd__o211ai_1 _3454_ (.A1(_0951_),
    .A2(_0956_),
    .B1(_1439_),
    .C1(_0942_),
    .Y(_1451_));
 sky130_fd_sc_hd__a32o_1 _3455_ (.A1(_1441_),
    .A2(_1451_),
    .A3(_1353_),
    .B1(net133),
    .B2(\acc[28] ),
    .X(_0304_));
 sky130_fd_sc_hd__o2111ai_2 _3456_ (.A1(_0969_),
    .A2(_1437_),
    .B1(_0955_),
    .C1(_0959_),
    .D1(_0964_),
    .Y(_1452_));
 sky130_fd_sc_hd__a21oi_1 _3457_ (.A1(_0955_),
    .A2(_1452_),
    .B1(_0958_),
    .Y(_1453_));
 sky130_fd_sc_hd__a31o_1 _3458_ (.A1(_0955_),
    .A2(_0958_),
    .A3(_1452_),
    .B1(_1354_),
    .X(_1454_));
 sky130_fd_sc_hd__a2bb2o_1 _3459_ (.A1_N(_1453_),
    .A2_N(_1454_),
    .B1(\acc[27] ),
    .B2(net133),
    .X(_0303_));
 sky130_fd_sc_hd__a22o_1 _3460_ (.A1(_0955_),
    .A2(_0959_),
    .B1(_0964_),
    .B2(_1438_),
    .X(_1455_));
 sky130_fd_sc_hd__a32o_1 _3461_ (.A1(_1455_),
    .A2(_1353_),
    .A3(_1452_),
    .B1(net133),
    .B2(\acc[26] ),
    .X(_0302_));
 sky130_fd_sc_hd__a41o_1 _3462_ (.A1(\acc[24] ),
    .A2(_1801_),
    .A3(_0965_),
    .A4(_0966_),
    .B1(_1437_),
    .X(_1456_));
 sky130_fd_sc_hd__xnor2_1 _3463_ (.A(_0975_),
    .B(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__a32o_1 _3464_ (.A1(\m[0] ),
    .A2(_1924_),
    .A3(_1457_),
    .B1(net133),
    .B2(\acc[25] ),
    .X(_0301_));
 sky130_fd_sc_hd__or4b_1 _3465_ (.A(net135),
    .B(_1923_),
    .C(_1437_),
    .D_N(\m[0] ),
    .X(_1458_));
 sky130_fd_sc_hd__a21oi_1 _3466_ (.A1(_0974_),
    .A2(_1162_),
    .B1(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__a21o_1 _3467_ (.A1(\acc[24] ),
    .A2(net133),
    .B1(_1459_),
    .X(_0300_));
 sky130_fd_sc_hd__a31o_1 _3468_ (.A1(_1159_),
    .A2(_1160_),
    .A3(_1106_),
    .B1(_1087_),
    .X(_1460_));
 sky130_fd_sc_hd__a21oi_2 _3469_ (.A1(_1460_),
    .A2(_1078_),
    .B1(_1013_),
    .Y(_1461_));
 sky130_fd_sc_hd__o31a_1 _3470_ (.A1(_1008_),
    .A2(_1021_),
    .A3(_1461_),
    .B1(_1024_),
    .X(_1462_));
 sky130_fd_sc_hd__o311a_1 _3471_ (.A1(_1008_),
    .A2(_1021_),
    .A3(_1461_),
    .B1(_1024_),
    .C1(_0987_),
    .X(_1463_));
 sky130_fd_sc_hd__or3_1 _3472_ (.A(_0985_),
    .B(_0997_),
    .C(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__o21ai_1 _3473_ (.A1(_0985_),
    .A2(_1463_),
    .B1(_0997_),
    .Y(_1465_));
 sky130_fd_sc_hd__a32o_1 _3474_ (.A1(_1464_),
    .A2(_1465_),
    .A3(_1353_),
    .B1(net133),
    .B2(\acc[23] ),
    .X(_0299_));
 sky130_fd_sc_hd__a21o_1 _3475_ (.A1(_0984_),
    .A2(_0986_),
    .B1(_1462_),
    .X(_1466_));
 sky130_fd_sc_hd__a21oi_1 _3476_ (.A1(_0987_),
    .A2(_1462_),
    .B1(_1354_),
    .Y(_1467_));
 sky130_fd_sc_hd__a22o_1 _3477_ (.A1(\acc[22] ),
    .A2(net133),
    .B1(_1467_),
    .B2(_1466_),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_1 _3478_ (.A1(_1008_),
    .A2(_1461_),
    .B1(_1025_),
    .Y(_1468_));
 sky130_fd_sc_hd__or3_1 _3479_ (.A(_1008_),
    .B(_1025_),
    .C(_1461_),
    .X(_1469_));
 sky130_fd_sc_hd__a32o_1 _3480_ (.A1(_1469_),
    .A2(_1353_),
    .A3(_1468_),
    .B1(net133),
    .B2(\acc[21] ),
    .X(_0297_));
 sky130_fd_sc_hd__and3_1 _3481_ (.A(_1013_),
    .B(_1460_),
    .C(_1078_),
    .X(_1470_));
 sky130_fd_sc_hd__or4b_1 _3482_ (.A(net135),
    .B(_1923_),
    .C(_1461_),
    .D_N(\m[0] ),
    .X(_1471_));
 sky130_fd_sc_hd__a2bb2o_1 _3483_ (.A1_N(_1470_),
    .A2_N(_1471_),
    .B1(\acc[20] ),
    .B2(net133),
    .X(_0296_));
 sky130_fd_sc_hd__a311o_1 _3484_ (.A1(_1159_),
    .A2(_1160_),
    .A3(_1106_),
    .B1(_1083_),
    .C1(_1048_),
    .X(_1472_));
 sky130_fd_sc_hd__a211o_1 _3485_ (.A1(_1161_),
    .A2(_1084_),
    .B1(_1048_),
    .C1(_1038_),
    .X(_1473_));
 sky130_fd_sc_hd__a31o_1 _3486_ (.A1(_1037_),
    .A2(_1061_),
    .A3(_1473_),
    .B1(_1062_),
    .X(_1474_));
 sky130_fd_sc_hd__a311o_1 _3487_ (.A1(_1037_),
    .A2(_1061_),
    .A3(_1473_),
    .B1(_1076_),
    .C1(_1062_),
    .X(_1475_));
 sky130_fd_sc_hd__or3b_1 _3488_ (.A(_1072_),
    .B(_1074_),
    .C_N(_1474_),
    .X(_1476_));
 sky130_fd_sc_hd__a32o_1 _3489_ (.A1(_1475_),
    .A2(_1476_),
    .A3(_1353_),
    .B1(net133),
    .B2(\acc[19] ),
    .X(_0295_));
 sky130_fd_sc_hd__or4b_1 _3490_ (.A(_1036_),
    .B(_1060_),
    .C(_1062_),
    .D_N(_1473_),
    .X(_1477_));
 sky130_fd_sc_hd__a311o_1 _3491_ (.A1(_1085_),
    .A2(_1086_),
    .A3(_1161_),
    .B1(_1064_),
    .C1(_1050_),
    .X(_1478_));
 sky130_fd_sc_hd__a32o_1 _3492_ (.A1(_1477_),
    .A2(_1478_),
    .A3(_1353_),
    .B1(net132),
    .B2(\acc[18] ),
    .X(_0294_));
 sky130_fd_sc_hd__a211o_1 _3493_ (.A1(_1049_),
    .A2(_1472_),
    .B1(_1036_),
    .C1(_1038_),
    .X(_1479_));
 sky130_fd_sc_hd__a211o_1 _3494_ (.A1(_1161_),
    .A2(_1084_),
    .B1(_1048_),
    .C1(_1086_),
    .X(_1480_));
 sky130_fd_sc_hd__a32o_1 _3495_ (.A1(_1479_),
    .A2(_1480_),
    .A3(_1353_),
    .B1(net132),
    .B2(\acc[17] ),
    .X(_0293_));
 sky130_fd_sc_hd__a21o_1 _3496_ (.A1(_1049_),
    .A2(_1084_),
    .B1(_1161_),
    .X(_1481_));
 sky130_fd_sc_hd__a32o_1 _3497_ (.A1(_1481_),
    .A2(_1353_),
    .A3(_1472_),
    .B1(net132),
    .B2(\acc[16] ),
    .X(_0292_));
 sky130_fd_sc_hd__a21o_1 _3498_ (.A1(_1153_),
    .A2(_1157_),
    .B1(_1097_),
    .X(_1482_));
 sky130_fd_sc_hd__a31o_1 _3499_ (.A1(_1096_),
    .A2(_1100_),
    .A3(_1482_),
    .B1(_1098_),
    .X(_1483_));
 sky130_fd_sc_hd__o21ai_1 _3500_ (.A1(_1093_),
    .A2(_1483_),
    .B1(_1091_),
    .Y(_1484_));
 sky130_fd_sc_hd__nand3_1 _3501_ (.A(_1089_),
    .B(_1090_),
    .C(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__a21o_1 _3502_ (.A1(_1089_),
    .A2(_1090_),
    .B1(_1484_),
    .X(_1486_));
 sky130_fd_sc_hd__a32o_1 _3503_ (.A1(_1486_),
    .A2(_1353_),
    .A3(_1485_),
    .B1(net132),
    .B2(\acc[15] ),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _3504_ (.A(_1093_),
    .B(_1483_),
    .Y(_1487_));
 sky130_fd_sc_hd__o211a_1 _3505_ (.A1(_1093_),
    .A2(_1483_),
    .B1(\m[0] ),
    .C1(_1924_),
    .X(_1488_));
 sky130_fd_sc_hd__a22o_1 _3506_ (.A1(\acc[14] ),
    .A2(net132),
    .B1(_1488_),
    .B2(_1487_),
    .X(_0290_));
 sky130_fd_sc_hd__a21o_1 _3507_ (.A1(_1096_),
    .A2(_1482_),
    .B1(_1101_),
    .X(_1489_));
 sky130_fd_sc_hd__nand3_1 _3508_ (.A(_1096_),
    .B(_1101_),
    .C(_1482_),
    .Y(_1490_));
 sky130_fd_sc_hd__a32o_1 _3509_ (.A1(_1489_),
    .A2(_1490_),
    .A3(_1353_),
    .B1(net132),
    .B2(\acc[13] ),
    .X(_0289_));
 sky130_fd_sc_hd__a221o_1 _3510_ (.A1(_1095_),
    .A2(_1096_),
    .B1(_1137_),
    .B2(_1152_),
    .C1(_1158_),
    .X(_1491_));
 sky130_fd_sc_hd__a32o_1 _3511_ (.A1(_1482_),
    .A2(_1491_),
    .A3(_1353_),
    .B1(net132),
    .B2(\acc[12] ),
    .X(_0288_));
 sky130_fd_sc_hd__a31o_1 _3512_ (.A1(_1137_),
    .A2(_1146_),
    .A3(_1147_),
    .B1(_1154_),
    .X(_1492_));
 sky130_fd_sc_hd__and3_1 _3513_ (.A(_1492_),
    .B(_1144_),
    .C(_1148_),
    .X(_1493_));
 sky130_fd_sc_hd__o211ai_1 _3514_ (.A1(_1142_),
    .A2(_1493_),
    .B1(_1139_),
    .C1(_1140_),
    .Y(_1494_));
 sky130_fd_sc_hd__a211o_1 _3515_ (.A1(_1139_),
    .A2(_1140_),
    .B1(_1142_),
    .C1(_1493_),
    .X(_1495_));
 sky130_fd_sc_hd__a32o_1 _3516_ (.A1(_1495_),
    .A2(_1353_),
    .A3(_1494_),
    .B1(net132),
    .B2(\acc[11] ),
    .X(_0287_));
 sky130_fd_sc_hd__a21oi_1 _3517_ (.A1(_1148_),
    .A2(_1492_),
    .B1(_1144_),
    .Y(_1496_));
 sky130_fd_sc_hd__or4b_1 _3518_ (.A(net135),
    .B(_1923_),
    .C(_1496_),
    .D_N(\m[0] ),
    .X(_1497_));
 sky130_fd_sc_hd__a2bb2o_1 _3519_ (.A1_N(_1493_),
    .A2_N(_1497_),
    .B1(\acc[10] ),
    .B2(net132),
    .X(_0286_));
 sky130_fd_sc_hd__a21bo_1 _3520_ (.A1(_1137_),
    .A2(_1146_),
    .B1_N(_1147_),
    .X(_1498_));
 sky130_fd_sc_hd__xnor2_1 _3521_ (.A(_1150_),
    .B(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__a32o_1 _3522_ (.A1(\m[0] ),
    .A2(_1924_),
    .A3(_1499_),
    .B1(net132),
    .B2(\acc[9] ),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_1 _3523_ (.A1(_1146_),
    .A2(_1147_),
    .B1(_1137_),
    .Y(_1500_));
 sky130_fd_sc_hd__a31o_1 _3524_ (.A1(_1137_),
    .A2(_1146_),
    .A3(_1147_),
    .B1(_1354_),
    .X(_1501_));
 sky130_fd_sc_hd__a2bb2o_1 _3525_ (.A1_N(_1500_),
    .A2_N(_1501_),
    .B1(\acc[8] ),
    .B2(net132),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _3526_ (.A(_1130_),
    .B(_1134_),
    .X(_1502_));
 sky130_fd_sc_hd__o21a_1 _3527_ (.A1(_0978_),
    .A2(_1131_),
    .B1(_1135_),
    .X(_1503_));
 sky130_fd_sc_hd__nand2_1 _3528_ (.A(_1128_),
    .B(_1129_),
    .Y(_1504_));
 sky130_fd_sc_hd__o211a_1 _3529_ (.A1(_0978_),
    .A2(_1131_),
    .B1(_1135_),
    .C1(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__o21ai_1 _3530_ (.A1(_1132_),
    .A2(_1505_),
    .B1(_1502_),
    .Y(_1506_));
 sky130_fd_sc_hd__or3_1 _3531_ (.A(_1132_),
    .B(_1502_),
    .C(_1505_),
    .X(_1507_));
 sky130_fd_sc_hd__a32o_1 _3532_ (.A1(_1507_),
    .A2(_1353_),
    .A3(_1506_),
    .B1(net132),
    .B2(\acc[7] ),
    .X(_0283_));
 sky130_fd_sc_hd__o21ai_1 _3533_ (.A1(_1503_),
    .A2(_1504_),
    .B1(_1353_),
    .Y(_1508_));
 sky130_fd_sc_hd__a2bb2o_1 _3534_ (.A1_N(_1505_),
    .A2_N(_1508_),
    .B1(\acc[6] ),
    .B2(net132),
    .X(_0282_));
 sky130_fd_sc_hd__a22o_1 _3535_ (.A1(_1108_),
    .A2(_1122_),
    .B1(_1125_),
    .B2(_1126_),
    .X(_1509_));
 sky130_fd_sc_hd__nand4_1 _3536_ (.A(_1108_),
    .B(_1122_),
    .C(_1125_),
    .D(_1126_),
    .Y(_1510_));
 sky130_fd_sc_hd__a32o_1 _3537_ (.A1(_1509_),
    .A2(_1510_),
    .A3(_1353_),
    .B1(net132),
    .B2(\acc[5] ),
    .X(_0281_));
 sky130_fd_sc_hd__a211o_1 _3538_ (.A1(_1111_),
    .A2(_1121_),
    .B1(_1109_),
    .C1(_1110_),
    .X(_1511_));
 sky130_fd_sc_hd__a32o_1 _3539_ (.A1(_1122_),
    .A2(_1511_),
    .A3(_1353_),
    .B1(\acc[4] ),
    .B2(net132),
    .X(_0280_));
 sky130_fd_sc_hd__o31a_1 _3540_ (.A1(net135),
    .A2(\count[4] ),
    .A3(_1112_),
    .B1(_1111_),
    .X(_1512_));
 sky130_fd_sc_hd__xor2_1 _3541_ (.A(_1120_),
    .B(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__a32o_1 _3542_ (.A1(\m[0] ),
    .A2(_1924_),
    .A3(_1513_),
    .B1(net132),
    .B2(\acc[3] ),
    .X(_0279_));
 sky130_fd_sc_hd__a21o_1 _3543_ (.A1(_1113_),
    .A2(_1114_),
    .B1(_1118_),
    .X(_1514_));
 sky130_fd_sc_hd__nand3_1 _3544_ (.A(_1118_),
    .B(_1114_),
    .C(_1113_),
    .Y(_1515_));
 sky130_fd_sc_hd__a32o_1 _3545_ (.A1(_1515_),
    .A2(_1353_),
    .A3(_1514_),
    .B1(net132),
    .B2(\acc[2] ),
    .X(_0278_));
 sky130_fd_sc_hd__a31o_1 _3546_ (.A1(\acc[1] ),
    .A2(_0648_),
    .A3(_1028_),
    .B1(_1115_),
    .X(_1516_));
 sky130_fd_sc_hd__nand2_1 _3547_ (.A(_1116_),
    .B(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__a311o_1 _3548_ (.A1(\acc[1] ),
    .A2(_0648_),
    .A3(_1028_),
    .B1(_1115_),
    .C1(_1116_),
    .X(_1518_));
 sky130_fd_sc_hd__a32o_1 _3549_ (.A1(_1517_),
    .A2(_1518_),
    .A3(_1353_),
    .B1(net132),
    .B2(\acc[1] ),
    .X(_0277_));
 sky130_fd_sc_hd__a31oi_1 _3550_ (.A1(\acc[0] ),
    .A2(_0897_),
    .A3(_1107_),
    .B1(_1923_),
    .Y(_1519_));
 sky130_fd_sc_hd__and4b_1 _3551_ (.A_N(net132),
    .B(_0648_),
    .C(_0897_),
    .D(_1803_),
    .X(_1520_));
 sky130_fd_sc_hd__o22a_1 _3552_ (.A1(_1519_),
    .A2(net132),
    .B1(\acc[0] ),
    .B2(_1520_),
    .X(_0276_));
 sky130_fd_sc_hd__nor2_1 _3553_ (.A(_1801_),
    .B(_1923_),
    .Y(_0275_));
 sky130_fd_sc_hd__and2b_4 _3554_ (.A_N(\state[0] ),
    .B(\state[1] ),
    .X(_1521_));
 sky130_fd_sc_hd__nand2b_4 _3555_ (.A_N(\state[0] ),
    .B(\state[1] ),
    .Y(_1522_));
 sky130_fd_sc_hd__a21o_1 _3556_ (.A1(_1816_),
    .A2(net67),
    .B1(_1521_),
    .X(_0273_));
 sky130_fd_sc_hd__or4_1 _3557_ (.A(\acc[39] ),
    .B(\acc[38] ),
    .C(\acc[37] ),
    .D(\acc[36] ),
    .X(_1523_));
 sky130_fd_sc_hd__nor2_1 _3558_ (.A(\acc[7] ),
    .B(\acc[6] ),
    .Y(_1524_));
 sky130_fd_sc_hd__nor3_1 _3559_ (.A(\acc[2] ),
    .B(\acc[1] ),
    .C(\acc[0] ),
    .Y(_1525_));
 sky130_fd_sc_hd__or3_1 _3560_ (.A(\acc[2] ),
    .B(\acc[1] ),
    .C(\acc[0] ),
    .X(_1526_));
 sky130_fd_sc_hd__or4_1 _3561_ (.A(\acc[3] ),
    .B(\acc[2] ),
    .C(\acc[1] ),
    .D(\acc[0] ),
    .X(_1527_));
 sky130_fd_sc_hd__nor2_1 _3562_ (.A(\acc[4] ),
    .B(\acc[3] ),
    .Y(_1528_));
 sky130_fd_sc_hd__or3_1 _3563_ (.A(\acc[4] ),
    .B(\acc[3] ),
    .C(_1526_),
    .X(_1529_));
 sky130_fd_sc_hd__or4_1 _3564_ (.A(\acc[5] ),
    .B(\acc[4] ),
    .C(\acc[3] ),
    .D(_1526_),
    .X(_1530_));
 sky130_fd_sc_hd__nand4_2 _3565_ (.A(_1525_),
    .B(_1799_),
    .C(_1524_),
    .D(_1528_),
    .Y(_1531_));
 sky130_fd_sc_hd__or4_1 _3566_ (.A(\acc[8] ),
    .B(\acc[7] ),
    .C(\acc[6] ),
    .D(_1530_),
    .X(_1532_));
 sky130_fd_sc_hd__nor2_1 _3567_ (.A(\acc[10] ),
    .B(\acc[9] ),
    .Y(_1533_));
 sky130_fd_sc_hd__or4_1 _3568_ (.A(\acc[10] ),
    .B(\acc[9] ),
    .C(\acc[8] ),
    .D(_1531_),
    .X(_1534_));
 sky130_fd_sc_hd__nor2_1 _3569_ (.A(\acc[12] ),
    .B(\acc[11] ),
    .Y(_1535_));
 sky130_fd_sc_hd__nand4b_2 _3570_ (.A_N(_1531_),
    .B(_1533_),
    .C(_1535_),
    .D(_1798_),
    .Y(_1536_));
 sky130_fd_sc_hd__or2_1 _3571_ (.A(\acc[14] ),
    .B(\acc[13] ),
    .X(_1537_));
 sky130_fd_sc_hd__or4_2 _3572_ (.A(\acc[12] ),
    .B(_1537_),
    .C(\acc[11] ),
    .D(_1534_),
    .X(_1538_));
 sky130_fd_sc_hd__or3_1 _3573_ (.A(\acc[18] ),
    .B(\acc[17] ),
    .C(\acc[16] ),
    .X(_1539_));
 sky130_fd_sc_hd__or3_1 _3574_ (.A(\acc[17] ),
    .B(\acc[16] ),
    .C(\acc[15] ),
    .X(_1540_));
 sky130_fd_sc_hd__nor2_1 _3575_ (.A(\acc[19] ),
    .B(\acc[18] ),
    .Y(_1541_));
 sky130_fd_sc_hd__or4_1 _3576_ (.A(\acc[19] ),
    .B(_1539_),
    .C(\acc[15] ),
    .D(_1538_),
    .X(_1542_));
 sky130_fd_sc_hd__nor4_1 _3577_ (.A(_1537_),
    .B(\acc[20] ),
    .C(_1536_),
    .D(_1540_),
    .Y(_1543_));
 sky130_fd_sc_hd__or4b_2 _3578_ (.A(_1540_),
    .B(\acc[20] ),
    .C(_1538_),
    .D_N(_1541_),
    .X(_1544_));
 sky130_fd_sc_hd__nor2_1 _3579_ (.A(\acc[23] ),
    .B(\acc[22] ),
    .Y(_1545_));
 sky130_fd_sc_hd__or4_4 _3580_ (.A(\acc[27] ),
    .B(\acc[26] ),
    .C(\acc[25] ),
    .D(\acc[24] ),
    .X(_1546_));
 sky130_fd_sc_hd__nand4_4 _3581_ (.A(_1543_),
    .B(_1797_),
    .C(_1541_),
    .D(_1545_),
    .Y(_1547_));
 sky130_fd_sc_hd__nor2_1 _3582_ (.A(_1546_),
    .B(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__or2_1 _3583_ (.A(_1546_),
    .B(_1547_),
    .X(_1549_));
 sky130_fd_sc_hd__nor4_2 _3584_ (.A(\acc[31] ),
    .B(\acc[30] ),
    .C(\acc[29] ),
    .D(\acc[28] ),
    .Y(_1550_));
 sky130_fd_sc_hd__or3b_2 _3585_ (.A(_1546_),
    .B(_1547_),
    .C_N(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__nor2_1 _3586_ (.A(\acc[33] ),
    .B(\acc[32] ),
    .Y(_1552_));
 sky130_fd_sc_hd__or3_2 _3587_ (.A(\acc[33] ),
    .B(\acc[32] ),
    .C(_1551_),
    .X(_1553_));
 sky130_fd_sc_hd__or3_2 _3588_ (.A(\acc[35] ),
    .B(\acc[34] ),
    .C(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__nor3_1 _3589_ (.A(\acc[35] ),
    .B(\acc[34] ),
    .C(_1523_),
    .Y(_1555_));
 sky130_fd_sc_hd__and4_1 _3590_ (.A(_1548_),
    .B(_1550_),
    .C(_1552_),
    .D(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__or4b_4 _3591_ (.A(\acc[33] ),
    .B(\acc[32] ),
    .C(_1551_),
    .D_N(_1555_),
    .X(_1557_));
 sky130_fd_sc_hd__or3_2 _3592_ (.A(\acc[42] ),
    .B(\acc[41] ),
    .C(\acc[40] ),
    .X(_1558_));
 sky130_fd_sc_hd__or3_1 _3593_ (.A(_1558_),
    .B(\acc[43] ),
    .C(_1557_),
    .X(_1559_));
 sky130_fd_sc_hd__nor4_1 _3594_ (.A(\acc[47] ),
    .B(\acc[46] ),
    .C(\acc[45] ),
    .D(\acc[44] ),
    .Y(_1560_));
 sky130_fd_sc_hd__nand4b_4 _3595_ (.A_N(_1558_),
    .B(_1788_),
    .C(_1556_),
    .D(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__or4_2 _3596_ (.A(\acc[51] ),
    .B(\acc[50] ),
    .C(\acc[49] ),
    .D(\acc[48] ),
    .X(_1562_));
 sky130_fd_sc_hd__or3_1 _3597_ (.A(_1562_),
    .B(\acc[52] ),
    .C(_1561_),
    .X(_1563_));
 sky130_fd_sc_hd__or3_1 _3598_ (.A(\acc[54] ),
    .B(\acc[53] ),
    .C(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__or4_1 _3599_ (.A(\acc[55] ),
    .B(\acc[53] ),
    .C(\acc[52] ),
    .D(_1562_),
    .X(_1565_));
 sky130_fd_sc_hd__or3_4 _3600_ (.A(_1565_),
    .B(\acc[54] ),
    .C(_1561_),
    .X(_1566_));
 sky130_fd_sc_hd__o31a_1 _3601_ (.A1(\acc[57] ),
    .A2(\acc[56] ),
    .A3(_1566_),
    .B1(net134),
    .X(_1567_));
 sky130_fd_sc_hd__a21oi_1 _3602_ (.A1(\acc[58] ),
    .A2(net134),
    .B1(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__o41a_1 _3603_ (.A1(\acc[58] ),
    .A2(\acc[57] ),
    .A3(\acc[56] ),
    .A4(_1566_),
    .B1(net134),
    .X(_1569_));
 sky130_fd_sc_hd__or4_2 _3604_ (.A(\acc[59] ),
    .B(\acc[58] ),
    .C(\acc[57] ),
    .D(\acc[56] ),
    .X(_1570_));
 sky130_fd_sc_hd__or3_1 _3605_ (.A(_1570_),
    .B(\acc[60] ),
    .C(_1566_),
    .X(_1571_));
 sky130_fd_sc_hd__or4_1 _3606_ (.A(\acc[61] ),
    .B(_1570_),
    .C(\acc[60] ),
    .D(_1566_),
    .X(_1572_));
 sky130_fd_sc_hd__o41a_1 _3607_ (.A1(\acc[61] ),
    .A2(_1570_),
    .A3(\acc[60] ),
    .A4(_1566_),
    .B1(net134),
    .X(_1573_));
 sky130_fd_sc_hd__a211oi_1 _3608_ (.A1(\acc[62] ),
    .A2(net134),
    .B1(\acc[63] ),
    .C1(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__o311a_1 _3609_ (.A1(\acc[62] ),
    .A2(\acc[61] ),
    .A3(_1571_),
    .B1(net134),
    .C1(\acc[63] ),
    .X(_1575_));
 sky130_fd_sc_hd__o21ai_1 _3610_ (.A1(_1574_),
    .A2(_1575_),
    .B1(_1521_),
    .Y(_1576_));
 sky130_fd_sc_hd__o21a_1 _3611_ (.A1(net127),
    .A2(_1521_),
    .B1(_1576_),
    .X(_0272_));
 sky130_fd_sc_hd__a21o_1 _3612_ (.A1(_1572_),
    .A2(net134),
    .B1(\acc[62] ),
    .X(_1577_));
 sky130_fd_sc_hd__nand2_1 _3613_ (.A(_1573_),
    .B(\acc[62] ),
    .Y(_1578_));
 sky130_fd_sc_hd__and3_1 _3614_ (.A(_1577_),
    .B(_1578_),
    .C(_1521_),
    .X(_1579_));
 sky130_fd_sc_hd__a21o_1 _3615_ (.A1(net126),
    .A2(_1522_),
    .B1(_1579_),
    .X(_0271_));
 sky130_fd_sc_hd__a21oi_1 _3616_ (.A1(_1571_),
    .A2(net134),
    .B1(\acc[61] ),
    .Y(_1580_));
 sky130_fd_sc_hd__o311a_1 _3617_ (.A1(_1570_),
    .A2(\acc[60] ),
    .A3(_1566_),
    .B1(net134),
    .C1(\acc[61] ),
    .X(_1581_));
 sky130_fd_sc_hd__o21ai_1 _3618_ (.A1(_1580_),
    .A2(_1581_),
    .B1(_1521_),
    .Y(_1582_));
 sky130_fd_sc_hd__o21a_1 _3619_ (.A1(net125),
    .A2(_1521_),
    .B1(_1582_),
    .X(_0270_));
 sky130_fd_sc_hd__a211o_1 _3620_ (.A1(\acc[59] ),
    .A2(net134),
    .B1(\acc[60] ),
    .C1(_1569_),
    .X(_1583_));
 sky130_fd_sc_hd__o211ai_1 _3621_ (.A1(_1566_),
    .A2(_1570_),
    .B1(\acc[60] ),
    .C1(net134),
    .Y(_1584_));
 sky130_fd_sc_hd__and3_1 _3622_ (.A(_1583_),
    .B(_1584_),
    .C(_1521_),
    .X(_1585_));
 sky130_fd_sc_hd__a21o_1 _3623_ (.A1(net124),
    .A2(_1522_),
    .B1(_1585_),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_1 _3624_ (.A(\acc[59] ),
    .B(_1568_),
    .Y(_1586_));
 sky130_fd_sc_hd__a21o_1 _3625_ (.A1(\acc[59] ),
    .A2(_1568_),
    .B1(_1522_),
    .X(_1587_));
 sky130_fd_sc_hd__o22a_1 _3626_ (.A1(net122),
    .A2(_1521_),
    .B1(_1586_),
    .B2(_1587_),
    .X(_0268_));
 sky130_fd_sc_hd__xor2_1 _3627_ (.A(\acc[58] ),
    .B(_1567_),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_1 _3628_ (.A0(_1588_),
    .A1(net121),
    .S(_1522_),
    .X(_0267_));
 sky130_fd_sc_hd__o31a_1 _3629_ (.A1(\acc[56] ),
    .A2(\acc[55] ),
    .A3(_1564_),
    .B1(net134),
    .X(_1589_));
 sky130_fd_sc_hd__o311a_1 _3630_ (.A1(\acc[56] ),
    .A2(\acc[55] ),
    .A3(_1564_),
    .B1(net134),
    .C1(\acc[57] ),
    .X(_1590_));
 sky130_fd_sc_hd__o21ai_1 _3631_ (.A1(\acc[57] ),
    .A2(_1589_),
    .B1(_1521_),
    .Y(_1591_));
 sky130_fd_sc_hd__a2bb2o_1 _3632_ (.A1_N(_1590_),
    .A2_N(_1591_),
    .B1(net120),
    .B2(_1522_),
    .X(_0266_));
 sky130_fd_sc_hd__and3_1 _3633_ (.A(_1566_),
    .B(net134),
    .C(\acc[56] ),
    .X(_1592_));
 sky130_fd_sc_hd__a21oi_1 _3634_ (.A1(_1566_),
    .A2(net134),
    .B1(\acc[56] ),
    .Y(_1593_));
 sky130_fd_sc_hd__or3_1 _3635_ (.A(_1593_),
    .B(_1522_),
    .C(_1592_),
    .X(_1594_));
 sky130_fd_sc_hd__a21bo_1 _3636_ (.A1(net119),
    .A2(_1522_),
    .B1_N(_1594_),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _3637_ (.A1(_1564_),
    .A2(net134),
    .B1(\acc[55] ),
    .Y(_1595_));
 sky130_fd_sc_hd__a31o_1 _3638_ (.A1(_1564_),
    .A2(net134),
    .A3(\acc[55] ),
    .B1(_1522_),
    .X(_1596_));
 sky130_fd_sc_hd__a2bb2o_1 _3639_ (.A1_N(_1595_),
    .A2_N(_1596_),
    .B1(net118),
    .B2(_1522_),
    .X(_0264_));
 sky130_fd_sc_hd__o21ai_1 _3640_ (.A1(\acc[53] ),
    .A2(_1563_),
    .B1(net134),
    .Y(_1597_));
 sky130_fd_sc_hd__o21ai_1 _3641_ (.A1(\acc[54] ),
    .A2(_1597_),
    .B1(_1521_),
    .Y(_1598_));
 sky130_fd_sc_hd__a21o_1 _3642_ (.A1(\acc[54] ),
    .A2(_1597_),
    .B1(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__o21a_1 _3643_ (.A1(net117),
    .A2(_1521_),
    .B1(_1599_),
    .X(_0263_));
 sky130_fd_sc_hd__o311a_1 _3644_ (.A1(_1562_),
    .A2(\acc[52] ),
    .A3(_1561_),
    .B1(net134),
    .C1(\acc[53] ),
    .X(_1600_));
 sky130_fd_sc_hd__a21oi_1 _3645_ (.A1(_1563_),
    .A2(net134),
    .B1(\acc[53] ),
    .Y(_1601_));
 sky130_fd_sc_hd__or3_1 _3646_ (.A(_1522_),
    .B(_1600_),
    .C(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__a21bo_1 _3647_ (.A1(net116),
    .A2(_1522_),
    .B1_N(_1602_),
    .X(_0262_));
 sky130_fd_sc_hd__o21a_1 _3648_ (.A1(_1561_),
    .A2(_1562_),
    .B1(net134),
    .X(_1603_));
 sky130_fd_sc_hd__o211a_1 _3649_ (.A1(_1561_),
    .A2(_1562_),
    .B1(\acc[52] ),
    .C1(net134),
    .X(_1604_));
 sky130_fd_sc_hd__nor2_1 _3650_ (.A(\acc[52] ),
    .B(_1603_),
    .Y(_1605_));
 sky130_fd_sc_hd__o21ai_1 _3651_ (.A1(_1604_),
    .A2(_1605_),
    .B1(_1521_),
    .Y(_1606_));
 sky130_fd_sc_hd__o21a_1 _3652_ (.A1(net115),
    .A2(_1521_),
    .B1(_1606_),
    .X(_0261_));
 sky130_fd_sc_hd__o31a_1 _3653_ (.A1(\acc[49] ),
    .A2(\acc[48] ),
    .A3(_1561_),
    .B1(net134),
    .X(_1607_));
 sky130_fd_sc_hd__a21oi_1 _3654_ (.A1(\acc[50] ),
    .A2(net134),
    .B1(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__nand2_1 _3655_ (.A(_1608_),
    .B(\acc[51] ),
    .Y(_1609_));
 sky130_fd_sc_hd__o21a_1 _3656_ (.A1(\acc[51] ),
    .A2(_1608_),
    .B1(_1521_),
    .X(_1610_));
 sky130_fd_sc_hd__o2bb2a_1 _3657_ (.A1_N(_1609_),
    .A2_N(_1610_),
    .B1(net114),
    .B2(_1521_),
    .X(_0260_));
 sky130_fd_sc_hd__o311a_1 _3658_ (.A1(\acc[49] ),
    .A2(\acc[48] ),
    .A3(_1561_),
    .B1(net134),
    .C1(\acc[50] ),
    .X(_1611_));
 sky130_fd_sc_hd__o21ai_1 _3659_ (.A1(\acc[50] ),
    .A2(_1607_),
    .B1(_1521_),
    .Y(_1612_));
 sky130_fd_sc_hd__a2bb2o_1 _3660_ (.A1_N(_1611_),
    .A2_N(_1612_),
    .B1(net113),
    .B2(_1522_),
    .X(_0259_));
 sky130_fd_sc_hd__o21a_1 _3661_ (.A1(\acc[48] ),
    .A2(_1561_),
    .B1(net134),
    .X(_1613_));
 sky130_fd_sc_hd__o211a_1 _3662_ (.A1(\acc[48] ),
    .A2(_1561_),
    .B1(net134),
    .C1(\acc[49] ),
    .X(_1614_));
 sky130_fd_sc_hd__o21ai_1 _3663_ (.A1(\acc[49] ),
    .A2(_1613_),
    .B1(_1521_),
    .Y(_1615_));
 sky130_fd_sc_hd__a2bb2o_1 _3664_ (.A1_N(_1614_),
    .A2_N(_1615_),
    .B1(net111),
    .B2(_1522_),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _3665_ (.A(_1561_),
    .B(net134),
    .C(\acc[48] ),
    .X(_1616_));
 sky130_fd_sc_hd__a21oi_1 _3666_ (.A1(_1561_),
    .A2(net134),
    .B1(\acc[48] ),
    .Y(_1617_));
 sky130_fd_sc_hd__or3_1 _3667_ (.A(_1617_),
    .B(_1522_),
    .C(_1616_),
    .X(_1618_));
 sky130_fd_sc_hd__a21bo_1 _3668_ (.A1(net110),
    .A2(_1522_),
    .B1_N(_1618_),
    .X(_0257_));
 sky130_fd_sc_hd__or4_1 _3669_ (.A(\acc[46] ),
    .B(\acc[45] ),
    .C(\acc[44] ),
    .D(_1559_),
    .X(_1619_));
 sky130_fd_sc_hd__o41a_1 _3670_ (.A1(\acc[44] ),
    .A2(_1558_),
    .A3(\acc[43] ),
    .A4(_1557_),
    .B1(net134),
    .X(_1620_));
 sky130_fd_sc_hd__a21oi_1 _3671_ (.A1(_1619_),
    .A2(net134),
    .B1(\acc[47] ),
    .Y(_1621_));
 sky130_fd_sc_hd__and3_1 _3672_ (.A(_1619_),
    .B(net134),
    .C(\acc[47] ),
    .X(_1622_));
 sky130_fd_sc_hd__nand2_1 _3673_ (.A(_1522_),
    .B(net109),
    .Y(_1623_));
 sky130_fd_sc_hd__o31ai_1 _3674_ (.A1(_1522_),
    .A2(_1621_),
    .A3(_1622_),
    .B1(_1623_),
    .Y(_0256_));
 sky130_fd_sc_hd__a211o_1 _3675_ (.A1(\acc[45] ),
    .A2(net134),
    .B1(\acc[46] ),
    .C1(_1620_),
    .X(_1624_));
 sky130_fd_sc_hd__o311a_1 _3676_ (.A1(\acc[45] ),
    .A2(\acc[44] ),
    .A3(_1559_),
    .B1(net134),
    .C1(\acc[46] ),
    .X(_1625_));
 sky130_fd_sc_hd__and3b_1 _3677_ (.A_N(_1625_),
    .B(_1521_),
    .C(_1624_),
    .X(_1626_));
 sky130_fd_sc_hd__a21o_1 _3678_ (.A1(net108),
    .A2(_1522_),
    .B1(_1626_),
    .X(_0255_));
 sky130_fd_sc_hd__o211a_1 _3679_ (.A1(\acc[44] ),
    .A2(_1559_),
    .B1(net134),
    .C1(\acc[45] ),
    .X(_1627_));
 sky130_fd_sc_hd__nor2_1 _3680_ (.A(\acc[45] ),
    .B(_1620_),
    .Y(_1628_));
 sky130_fd_sc_hd__o21ai_1 _3681_ (.A1(_1627_),
    .A2(_1628_),
    .B1(_1521_),
    .Y(_1629_));
 sky130_fd_sc_hd__o21a_1 _3682_ (.A1(net107),
    .A2(_1521_),
    .B1(_1629_),
    .X(_0254_));
 sky130_fd_sc_hd__o311a_1 _3683_ (.A1(_1558_),
    .A2(\acc[43] ),
    .A3(_1557_),
    .B1(net134),
    .C1(\acc[44] ),
    .X(_1630_));
 sky130_fd_sc_hd__a21oi_1 _3684_ (.A1(_1559_),
    .A2(net134),
    .B1(\acc[44] ),
    .Y(_1631_));
 sky130_fd_sc_hd__o21ai_1 _3685_ (.A1(_1630_),
    .A2(_1631_),
    .B1(_1521_),
    .Y(_1632_));
 sky130_fd_sc_hd__o21a_1 _3686_ (.A1(net106),
    .A2(_1521_),
    .B1(_1632_),
    .X(_0253_));
 sky130_fd_sc_hd__o31a_1 _3687_ (.A1(_1523_),
    .A2(_1554_),
    .A3(_1558_),
    .B1(net134),
    .X(_1633_));
 sky130_fd_sc_hd__o311a_1 _3688_ (.A1(_1523_),
    .A2(_1554_),
    .A3(_1558_),
    .B1(net134),
    .C1(_1788_),
    .X(_1634_));
 sky130_fd_sc_hd__o21ai_1 _3689_ (.A1(_1788_),
    .A2(_1633_),
    .B1(_1521_),
    .Y(_1635_));
 sky130_fd_sc_hd__o22a_1 _3690_ (.A1(net105),
    .A2(_1521_),
    .B1(_1635_),
    .B2(_1634_),
    .X(_0252_));
 sky130_fd_sc_hd__o31ai_1 _3691_ (.A1(\acc[41] ),
    .A2(\acc[40] ),
    .A3(_1557_),
    .B1(net134),
    .Y(_1636_));
 sky130_fd_sc_hd__o21ai_1 _3692_ (.A1(\acc[42] ),
    .A2(_1636_),
    .B1(_1521_),
    .Y(_1637_));
 sky130_fd_sc_hd__a21o_1 _3693_ (.A1(\acc[42] ),
    .A2(_1636_),
    .B1(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__o21a_1 _3694_ (.A1(net104),
    .A2(_1521_),
    .B1(_1638_),
    .X(_0251_));
 sky130_fd_sc_hd__o21ai_1 _3695_ (.A1(\acc[40] ),
    .A2(_1557_),
    .B1(net134),
    .Y(_1639_));
 sky130_fd_sc_hd__nor2_1 _3696_ (.A(\acc[41] ),
    .B(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__a21o_1 _3697_ (.A1(\acc[41] ),
    .A2(_1639_),
    .B1(_1522_),
    .X(_1641_));
 sky130_fd_sc_hd__o22a_1 _3698_ (.A1(net103),
    .A2(_1521_),
    .B1(_1640_),
    .B2(_1641_),
    .X(_0250_));
 sky130_fd_sc_hd__and3_1 _3699_ (.A(_1557_),
    .B(net134),
    .C(\acc[40] ),
    .X(_1642_));
 sky130_fd_sc_hd__a21oi_1 _3700_ (.A1(_1557_),
    .A2(net134),
    .B1(\acc[40] ),
    .Y(_1643_));
 sky130_fd_sc_hd__or3_1 _3701_ (.A(_1643_),
    .B(_1522_),
    .C(_1642_),
    .X(_1644_));
 sky130_fd_sc_hd__a21bo_1 _3702_ (.A1(net102),
    .A2(_1522_),
    .B1_N(_1644_),
    .X(_0249_));
 sky130_fd_sc_hd__o41ai_1 _3703_ (.A1(\acc[38] ),
    .A2(\acc[37] ),
    .A3(\acc[36] ),
    .A4(_1554_),
    .B1(net134),
    .Y(_1645_));
 sky130_fd_sc_hd__nor2_1 _3704_ (.A(\acc[39] ),
    .B(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__a21o_1 _3705_ (.A1(\acc[39] ),
    .A2(_1645_),
    .B1(_1522_),
    .X(_1647_));
 sky130_fd_sc_hd__o22a_1 _3706_ (.A1(net100),
    .A2(_1521_),
    .B1(_1646_),
    .B2(_1647_),
    .X(_0248_));
 sky130_fd_sc_hd__or3_1 _3707_ (.A(\acc[37] ),
    .B(\acc[36] ),
    .C(_1554_),
    .X(_1648_));
 sky130_fd_sc_hd__o311a_1 _3708_ (.A1(\acc[37] ),
    .A2(\acc[36] ),
    .A3(_1554_),
    .B1(net134),
    .C1(\acc[38] ),
    .X(_1649_));
 sky130_fd_sc_hd__a21oi_1 _3709_ (.A1(_1648_),
    .A2(net134),
    .B1(\acc[38] ),
    .Y(_1650_));
 sky130_fd_sc_hd__nand2_1 _3710_ (.A(_1522_),
    .B(net99),
    .Y(_1651_));
 sky130_fd_sc_hd__o31ai_1 _3711_ (.A1(_1522_),
    .A2(_1649_),
    .A3(_1650_),
    .B1(_1651_),
    .Y(_0247_));
 sky130_fd_sc_hd__o41a_1 _3712_ (.A1(\acc[36] ),
    .A2(\acc[35] ),
    .A3(\acc[34] ),
    .A4(_1553_),
    .B1(net134),
    .X(_1652_));
 sky130_fd_sc_hd__nor2_1 _3713_ (.A(\acc[37] ),
    .B(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__o211a_1 _3714_ (.A1(\acc[36] ),
    .A2(_1554_),
    .B1(net134),
    .C1(\acc[37] ),
    .X(_1654_));
 sky130_fd_sc_hd__o21ai_1 _3715_ (.A1(_1653_),
    .A2(_1654_),
    .B1(_1521_),
    .Y(_1655_));
 sky130_fd_sc_hd__o21a_1 _3716_ (.A1(net98),
    .A2(_1521_),
    .B1(_1655_),
    .X(_0246_));
 sky130_fd_sc_hd__o311a_1 _3717_ (.A1(\acc[35] ),
    .A2(\acc[34] ),
    .A3(_1553_),
    .B1(net134),
    .C1(\acc[36] ),
    .X(_1656_));
 sky130_fd_sc_hd__a21oi_1 _3718_ (.A1(_1554_),
    .A2(net134),
    .B1(\acc[36] ),
    .Y(_1657_));
 sky130_fd_sc_hd__o21ai_1 _3719_ (.A1(_1656_),
    .A2(_1657_),
    .B1(_1521_),
    .Y(_1658_));
 sky130_fd_sc_hd__o21a_1 _3720_ (.A1(net97),
    .A2(_1521_),
    .B1(_1658_),
    .X(_0245_));
 sky130_fd_sc_hd__o41a_1 _3721_ (.A1(\acc[34] ),
    .A2(\acc[33] ),
    .A3(\acc[32] ),
    .A4(_1551_),
    .B1(net134),
    .X(_1659_));
 sky130_fd_sc_hd__o211a_1 _3722_ (.A1(\acc[34] ),
    .A2(_1553_),
    .B1(net134),
    .C1(\acc[35] ),
    .X(_1660_));
 sky130_fd_sc_hd__o21ai_1 _3723_ (.A1(\acc[35] ),
    .A2(_1659_),
    .B1(_1521_),
    .Y(_1661_));
 sky130_fd_sc_hd__a2bb2o_1 _3724_ (.A1_N(_1660_),
    .A2_N(_1661_),
    .B1(net96),
    .B2(_1522_),
    .X(_0244_));
 sky130_fd_sc_hd__o311a_1 _3725_ (.A1(\acc[33] ),
    .A2(\acc[32] ),
    .A3(_1551_),
    .B1(net134),
    .C1(\acc[34] ),
    .X(_1662_));
 sky130_fd_sc_hd__a21oi_1 _3726_ (.A1(_1553_),
    .A2(net134),
    .B1(\acc[34] ),
    .Y(_1663_));
 sky130_fd_sc_hd__o21ai_1 _3727_ (.A1(_1662_),
    .A2(_1663_),
    .B1(_1521_),
    .Y(_1664_));
 sky130_fd_sc_hd__o21a_1 _3728_ (.A1(net95),
    .A2(_1521_),
    .B1(_1664_),
    .X(_0243_));
 sky130_fd_sc_hd__o21ai_1 _3729_ (.A1(\acc[32] ),
    .A2(_1551_),
    .B1(net134),
    .Y(_1665_));
 sky130_fd_sc_hd__xor2_1 _3730_ (.A(_1795_),
    .B(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _3731_ (.A0(_1666_),
    .A1(net94),
    .S(_1522_),
    .X(_0242_));
 sky130_fd_sc_hd__and3_1 _3732_ (.A(_1551_),
    .B(net134),
    .C(\acc[32] ),
    .X(_1667_));
 sky130_fd_sc_hd__a21oi_1 _3733_ (.A1(_1551_),
    .A2(net134),
    .B1(\acc[32] ),
    .Y(_1668_));
 sky130_fd_sc_hd__o21ai_1 _3734_ (.A1(_1667_),
    .A2(_1668_),
    .B1(_1521_),
    .Y(_1669_));
 sky130_fd_sc_hd__o21a_1 _3735_ (.A1(net93),
    .A2(_1521_),
    .B1(_1669_),
    .X(_0241_));
 sky130_fd_sc_hd__o31a_1 _3736_ (.A1(\acc[29] ),
    .A2(\acc[28] ),
    .A3(_1549_),
    .B1(net134),
    .X(_1670_));
 sky130_fd_sc_hd__a21oi_1 _3737_ (.A1(\acc[30] ),
    .A2(net134),
    .B1(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__o21ai_1 _3738_ (.A1(\acc[31] ),
    .A2(_1671_),
    .B1(_1521_),
    .Y(_1672_));
 sky130_fd_sc_hd__a21o_1 _3739_ (.A1(\acc[31] ),
    .A2(_1671_),
    .B1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__o21a_1 _3740_ (.A1(net92),
    .A2(_1521_),
    .B1(_1673_),
    .X(_0240_));
 sky130_fd_sc_hd__xor2_1 _3741_ (.A(\acc[30] ),
    .B(_1670_),
    .X(_1674_));
 sky130_fd_sc_hd__mux2_1 _3742_ (.A0(_1674_),
    .A1(net91),
    .S(_1522_),
    .X(_0239_));
 sky130_fd_sc_hd__o31a_1 _3743_ (.A1(\acc[28] ),
    .A2(_1546_),
    .A3(_1547_),
    .B1(net134),
    .X(_1675_));
 sky130_fd_sc_hd__nor2_1 _3744_ (.A(\acc[29] ),
    .B(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__o311a_1 _3745_ (.A1(\acc[28] ),
    .A2(_1546_),
    .A3(_1547_),
    .B1(net134),
    .C1(\acc[29] ),
    .X(_1677_));
 sky130_fd_sc_hd__o21ai_1 _3746_ (.A1(_1676_),
    .A2(_1677_),
    .B1(_1521_),
    .Y(_1678_));
 sky130_fd_sc_hd__o21a_1 _3747_ (.A1(net89),
    .A2(_1521_),
    .B1(_1678_),
    .X(_0238_));
 sky130_fd_sc_hd__and3_1 _3748_ (.A(_1549_),
    .B(net134),
    .C(\acc[28] ),
    .X(_1679_));
 sky130_fd_sc_hd__a21oi_1 _3749_ (.A1(_1549_),
    .A2(net134),
    .B1(\acc[28] ),
    .Y(_1680_));
 sky130_fd_sc_hd__o21ai_1 _3750_ (.A1(_1679_),
    .A2(_1680_),
    .B1(_1521_),
    .Y(_1681_));
 sky130_fd_sc_hd__o21a_1 _3751_ (.A1(net88),
    .A2(_1521_),
    .B1(_1681_),
    .X(_0237_));
 sky130_fd_sc_hd__or3_1 _3752_ (.A(\acc[25] ),
    .B(\acc[24] ),
    .C(_1547_),
    .X(_1682_));
 sky130_fd_sc_hd__o41a_2 _3753_ (.A1(\acc[23] ),
    .A2(\acc[22] ),
    .A3(\acc[21] ),
    .A4(_1544_),
    .B1(net134),
    .X(_1683_));
 sky130_fd_sc_hd__o41a_1 _3754_ (.A1(\acc[26] ),
    .A2(\acc[25] ),
    .A3(\acc[24] ),
    .A4(_1547_),
    .B1(net134),
    .X(_1684_));
 sky130_fd_sc_hd__xor2_1 _3755_ (.A(\acc[27] ),
    .B(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__mux2_1 _3756_ (.A0(_1685_),
    .A1(net87),
    .S(_1522_),
    .X(_0236_));
 sky130_fd_sc_hd__o311a_1 _3757_ (.A1(\acc[25] ),
    .A2(\acc[24] ),
    .A3(_1547_),
    .B1(net134),
    .C1(\acc[26] ),
    .X(_1686_));
 sky130_fd_sc_hd__a21oi_1 _3758_ (.A1(_1682_),
    .A2(net134),
    .B1(\acc[26] ),
    .Y(_1687_));
 sky130_fd_sc_hd__or3_1 _3759_ (.A(_1522_),
    .B(_1686_),
    .C(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__a21bo_1 _3760_ (.A1(net86),
    .A2(_1522_),
    .B1_N(_1688_),
    .X(_0235_));
 sky130_fd_sc_hd__a211o_1 _3761_ (.A1(\acc[24] ),
    .A2(net134),
    .B1(_1683_),
    .C1(\acc[25] ),
    .X(_1689_));
 sky130_fd_sc_hd__o211ai_1 _3762_ (.A1(\acc[24] ),
    .A2(_1547_),
    .B1(net134),
    .C1(\acc[25] ),
    .Y(_1690_));
 sky130_fd_sc_hd__and3_1 _3763_ (.A(_1689_),
    .B(_1690_),
    .C(_1521_),
    .X(_1691_));
 sky130_fd_sc_hd__a21o_1 _3764_ (.A1(net85),
    .A2(_1522_),
    .B1(_1691_),
    .X(_0234_));
 sky130_fd_sc_hd__o21ai_1 _3765_ (.A1(\acc[24] ),
    .A2(_1683_),
    .B1(_1521_),
    .Y(_1692_));
 sky130_fd_sc_hd__a21oi_1 _3766_ (.A1(\acc[24] ),
    .A2(_1683_),
    .B1(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__a21o_1 _3767_ (.A1(net84),
    .A2(_1522_),
    .B1(_1693_),
    .X(_0233_));
 sky130_fd_sc_hd__o31a_1 _3768_ (.A1(\acc[22] ),
    .A2(\acc[21] ),
    .A3(_1544_),
    .B1(net134),
    .X(_1694_));
 sky130_fd_sc_hd__xor2_1 _3769_ (.A(\acc[23] ),
    .B(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__mux2_1 _3770_ (.A0(_1695_),
    .A1(net83),
    .S(_1522_),
    .X(_0232_));
 sky130_fd_sc_hd__o21ai_1 _3771_ (.A1(\acc[21] ),
    .A2(_1544_),
    .B1(net134),
    .Y(_1696_));
 sky130_fd_sc_hd__xnor2_1 _3772_ (.A(\acc[22] ),
    .B(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(_1697_),
    .A1(net82),
    .S(_1522_),
    .X(_0231_));
 sky130_fd_sc_hd__a21oi_1 _3774_ (.A1(_1544_),
    .A2(net134),
    .B1(_1797_),
    .Y(_1698_));
 sky130_fd_sc_hd__a31o_1 _3775_ (.A1(_1797_),
    .A2(_1544_),
    .A3(net134),
    .B1(_1522_),
    .X(_1699_));
 sky130_fd_sc_hd__o22a_1 _3776_ (.A1(net81),
    .A2(_1521_),
    .B1(_1698_),
    .B2(_1699_),
    .X(_0230_));
 sky130_fd_sc_hd__and3_1 _3777_ (.A(_1542_),
    .B(net134),
    .C(\acc[20] ),
    .X(_1700_));
 sky130_fd_sc_hd__a21oi_1 _3778_ (.A1(_1542_),
    .A2(net134),
    .B1(\acc[20] ),
    .Y(_1701_));
 sky130_fd_sc_hd__or3_1 _3779_ (.A(_1701_),
    .B(_1522_),
    .C(_1700_),
    .X(_1702_));
 sky130_fd_sc_hd__a21bo_1 _3780_ (.A1(net80),
    .A2(_1522_),
    .B1_N(_1702_),
    .X(_0229_));
 sky130_fd_sc_hd__o31a_1 _3781_ (.A1(_1539_),
    .A2(\acc[15] ),
    .A3(_1538_),
    .B1(net134),
    .X(_1703_));
 sky130_fd_sc_hd__or2_1 _3782_ (.A(\acc[19] ),
    .B(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__a21oi_1 _3783_ (.A1(\acc[19] ),
    .A2(_1703_),
    .B1(_1522_),
    .Y(_1705_));
 sky130_fd_sc_hd__a22o_1 _3784_ (.A1(net78),
    .A2(_1522_),
    .B1(_1704_),
    .B2(_1705_),
    .X(_0228_));
 sky130_fd_sc_hd__o21ai_1 _3785_ (.A1(\acc[15] ),
    .A2(_1538_),
    .B1(net134),
    .Y(_1706_));
 sky130_fd_sc_hd__o31a_1 _3786_ (.A1(_1536_),
    .A2(_1537_),
    .A3(_1540_),
    .B1(net134),
    .X(_1707_));
 sky130_fd_sc_hd__xor2_1 _3787_ (.A(\acc[18] ),
    .B(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__mux2_1 _3788_ (.A0(_1708_),
    .A1(net77),
    .S(_1522_),
    .X(_0227_));
 sky130_fd_sc_hd__o31ai_1 _3789_ (.A1(\acc[16] ),
    .A2(\acc[15] ),
    .A3(_1538_),
    .B1(net134),
    .Y(_1709_));
 sky130_fd_sc_hd__a21oi_1 _3790_ (.A1(\acc[17] ),
    .A2(_1709_),
    .B1(_1522_),
    .Y(_1710_));
 sky130_fd_sc_hd__o21ai_1 _3791_ (.A1(\acc[17] ),
    .A2(_1709_),
    .B1(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__o21a_1 _3792_ (.A1(net76),
    .A2(_1521_),
    .B1(_1711_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _3793_ (.A(net75),
    .B(_1521_),
    .X(_1712_));
 sky130_fd_sc_hd__nor2_1 _3794_ (.A(\acc[16] ),
    .B(_1706_),
    .Y(_1713_));
 sky130_fd_sc_hd__and2_1 _3795_ (.A(_1706_),
    .B(\acc[16] ),
    .X(_1714_));
 sky130_fd_sc_hd__o31a_1 _3796_ (.A1(_1522_),
    .A2(_1713_),
    .A3(_1714_),
    .B1(_1712_),
    .X(_0225_));
 sky130_fd_sc_hd__a21oi_1 _3797_ (.A1(_1538_),
    .A2(net134),
    .B1(\acc[15] ),
    .Y(_1715_));
 sky130_fd_sc_hd__o311a_1 _3798_ (.A1(\acc[14] ),
    .A2(\acc[13] ),
    .A3(_1536_),
    .B1(net134),
    .C1(\acc[15] ),
    .X(_1716_));
 sky130_fd_sc_hd__o21ai_1 _3799_ (.A1(_1715_),
    .A2(_1716_),
    .B1(_1521_),
    .Y(_1717_));
 sky130_fd_sc_hd__o21a_1 _3800_ (.A1(net74),
    .A2(_1521_),
    .B1(_1717_),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _3801_ (.A(_1536_),
    .B(net134),
    .Y(_1718_));
 sky130_fd_sc_hd__nand2_1 _3802_ (.A(\acc[13] ),
    .B(net134),
    .Y(_1719_));
 sky130_fd_sc_hd__and3_1 _3803_ (.A(_1718_),
    .B(_1719_),
    .C(\acc[14] ),
    .X(_1720_));
 sky130_fd_sc_hd__a21oi_1 _3804_ (.A1(_1718_),
    .A2(_1719_),
    .B1(\acc[14] ),
    .Y(_1721_));
 sky130_fd_sc_hd__or2_1 _3805_ (.A(net73),
    .B(_1521_),
    .X(_1722_));
 sky130_fd_sc_hd__o31a_1 _3806_ (.A1(_1721_),
    .A2(_1522_),
    .A3(_1720_),
    .B1(_1722_),
    .X(_0223_));
 sky130_fd_sc_hd__o21ai_1 _3807_ (.A1(\acc[13] ),
    .A2(_1718_),
    .B1(_1521_),
    .Y(_1723_));
 sky130_fd_sc_hd__a21o_1 _3808_ (.A1(\acc[13] ),
    .A2(_1718_),
    .B1(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__o21a_1 _3809_ (.A1(net72),
    .A2(_1521_),
    .B1(_1724_),
    .X(_0222_));
 sky130_fd_sc_hd__o21ai_1 _3810_ (.A1(\acc[11] ),
    .A2(_1534_),
    .B1(sign),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _3811_ (.A(_1725_),
    .B(\acc[12] ),
    .Y(_1726_));
 sky130_fd_sc_hd__o21a_1 _3812_ (.A1(\acc[12] ),
    .A2(_1725_),
    .B1(_1521_),
    .X(_1727_));
 sky130_fd_sc_hd__o2bb2a_1 _3813_ (.A1_N(_1726_),
    .A2_N(_1727_),
    .B1(net71),
    .B2(_1521_),
    .X(_0221_));
 sky130_fd_sc_hd__a21oi_1 _3814_ (.A1(_1534_),
    .A2(sign),
    .B1(\acc[11] ),
    .Y(_1728_));
 sky130_fd_sc_hd__o311a_1 _3815_ (.A1(\acc[10] ),
    .A2(\acc[9] ),
    .A3(_1532_),
    .B1(sign),
    .C1(\acc[11] ),
    .X(_1729_));
 sky130_fd_sc_hd__o21ai_1 _3816_ (.A1(_1728_),
    .A2(_1729_),
    .B1(_1521_),
    .Y(_1730_));
 sky130_fd_sc_hd__o21a_1 _3817_ (.A1(net70),
    .A2(_1521_),
    .B1(_1730_),
    .X(_0220_));
 sky130_fd_sc_hd__o31a_1 _3818_ (.A1(\acc[9] ),
    .A2(\acc[8] ),
    .A3(_1531_),
    .B1(sign),
    .X(_1731_));
 sky130_fd_sc_hd__o311a_1 _3819_ (.A1(\acc[9] ),
    .A2(\acc[8] ),
    .A3(_1531_),
    .B1(sign),
    .C1(\acc[10] ),
    .X(_1732_));
 sky130_fd_sc_hd__o21ai_1 _3820_ (.A1(\acc[10] ),
    .A2(_1731_),
    .B1(_1521_),
    .Y(_1733_));
 sky130_fd_sc_hd__a2bb2o_1 _3821_ (.A1_N(_1732_),
    .A2_N(_1733_),
    .B1(net69),
    .B2(_1522_),
    .X(_0219_));
 sky130_fd_sc_hd__and3_1 _3822_ (.A(_1532_),
    .B(sign),
    .C(\acc[9] ),
    .X(_1734_));
 sky130_fd_sc_hd__a21oi_1 _3823_ (.A1(_1532_),
    .A2(sign),
    .B1(\acc[9] ),
    .Y(_1735_));
 sky130_fd_sc_hd__o21ai_1 _3824_ (.A1(_1734_),
    .A2(_1735_),
    .B1(_1521_),
    .Y(_1736_));
 sky130_fd_sc_hd__o21a_1 _3825_ (.A1(net131),
    .A2(_1521_),
    .B1(_1736_),
    .X(_0218_));
 sky130_fd_sc_hd__a21oi_1 _3826_ (.A1(_1531_),
    .A2(sign),
    .B1(_1798_),
    .Y(_1737_));
 sky130_fd_sc_hd__a31o_1 _3827_ (.A1(_1798_),
    .A2(_1531_),
    .A3(sign),
    .B1(_1522_),
    .X(_1738_));
 sky130_fd_sc_hd__o22a_1 _3828_ (.A1(net130),
    .A2(_1521_),
    .B1(_1737_),
    .B2(_1738_),
    .X(_0217_));
 sky130_fd_sc_hd__o31a_1 _3829_ (.A1(\acc[6] ),
    .A2(\acc[5] ),
    .A3(_1529_),
    .B1(sign),
    .X(_1739_));
 sky130_fd_sc_hd__xor2_1 _3830_ (.A(\acc[7] ),
    .B(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__mux2_1 _3831_ (.A0(_1740_),
    .A1(net129),
    .S(_1522_),
    .X(_0216_));
 sky130_fd_sc_hd__a21oi_1 _3832_ (.A1(_1530_),
    .A2(sign),
    .B1(\acc[6] ),
    .Y(_1741_));
 sky130_fd_sc_hd__o311a_1 _3833_ (.A1(\acc[5] ),
    .A2(\acc[4] ),
    .A3(_1527_),
    .B1(sign),
    .C1(\acc[6] ),
    .X(_1742_));
 sky130_fd_sc_hd__o21ai_1 _3834_ (.A1(_1741_),
    .A2(_1742_),
    .B1(_1521_),
    .Y(_1743_));
 sky130_fd_sc_hd__o21a_1 _3835_ (.A1(net128),
    .A2(_1521_),
    .B1(_1743_),
    .X(_0215_));
 sky130_fd_sc_hd__a21oi_1 _3836_ (.A1(_1529_),
    .A2(sign),
    .B1(_1799_),
    .Y(_1744_));
 sky130_fd_sc_hd__a31o_1 _3837_ (.A1(_1799_),
    .A2(_1529_),
    .A3(sign),
    .B1(_1522_),
    .X(_1745_));
 sky130_fd_sc_hd__o22a_1 _3838_ (.A1(net123),
    .A2(_1521_),
    .B1(_1744_),
    .B2(_1745_),
    .X(_0214_));
 sky130_fd_sc_hd__a21oi_1 _3839_ (.A1(_1527_),
    .A2(sign),
    .B1(\acc[4] ),
    .Y(_1746_));
 sky130_fd_sc_hd__and3_1 _3840_ (.A(_1527_),
    .B(sign),
    .C(\acc[4] ),
    .X(_1747_));
 sky130_fd_sc_hd__o21ai_1 _3841_ (.A1(_1746_),
    .A2(_1747_),
    .B1(_1521_),
    .Y(_1748_));
 sky130_fd_sc_hd__o21a_1 _3842_ (.A1(net112),
    .A2(_1521_),
    .B1(_1748_),
    .X(_0213_));
 sky130_fd_sc_hd__o311a_1 _3843_ (.A1(\acc[2] ),
    .A2(\acc[1] ),
    .A3(\acc[0] ),
    .B1(sign),
    .C1(\acc[3] ),
    .X(_1749_));
 sky130_fd_sc_hd__a21oi_1 _3844_ (.A1(_1526_),
    .A2(sign),
    .B1(\acc[3] ),
    .Y(_1750_));
 sky130_fd_sc_hd__o21ai_1 _3845_ (.A1(_1749_),
    .A2(_1750_),
    .B1(_1521_),
    .Y(_1751_));
 sky130_fd_sc_hd__o21a_1 _3846_ (.A1(net101),
    .A2(_1521_),
    .B1(_1751_),
    .X(_0212_));
 sky130_fd_sc_hd__o21a_1 _3847_ (.A1(\acc[1] ),
    .A2(\acc[0] ),
    .B1(sign),
    .X(_1752_));
 sky130_fd_sc_hd__or2_1 _3848_ (.A(\acc[2] ),
    .B(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__a21oi_1 _3849_ (.A1(\acc[2] ),
    .A2(_1752_),
    .B1(_1522_),
    .Y(_1754_));
 sky130_fd_sc_hd__a22o_1 _3850_ (.A1(net90),
    .A2(_1522_),
    .B1(_1753_),
    .B2(_1754_),
    .X(_0211_));
 sky130_fd_sc_hd__and3_1 _3851_ (.A(\acc[1] ),
    .B(\acc[0] ),
    .C(sign),
    .X(_1755_));
 sky130_fd_sc_hd__a21oi_1 _3852_ (.A1(\acc[0] ),
    .A2(sign),
    .B1(\acc[1] ),
    .Y(_1756_));
 sky130_fd_sc_hd__o21ai_1 _3853_ (.A1(_1755_),
    .A2(_1756_),
    .B1(_1521_),
    .Y(_1757_));
 sky130_fd_sc_hd__o21a_1 _3854_ (.A1(net79),
    .A2(_1521_),
    .B1(_1757_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _3855_ (.A0(net68),
    .A1(\acc[0] ),
    .S(_1521_),
    .X(_0209_));
 sky130_fd_sc_hd__xor2_1 _3856_ (.A(net57),
    .B(net25),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _3857_ (.A0(net134),
    .A1(_1758_),
    .S(_1817_),
    .X(_0208_));
 sky130_fd_sc_hd__a32o_1 _3858_ (.A1(_1922_),
    .A2(_0544_),
    .A3(_0549_),
    .B1(_1818_),
    .B2(\count[5] ),
    .X(_0207_));
 sky130_fd_sc_hd__o21ai_1 _3859_ (.A1(_1923_),
    .A2(_0549_),
    .B1(_0274_),
    .Y(_1759_));
 sky130_fd_sc_hd__and3_1 _3860_ (.A(_1922_),
    .B(_0549_),
    .C(_0648_),
    .X(_1760_));
 sky130_fd_sc_hd__a21o_1 _3861_ (.A1(\count[4] ),
    .A2(_1759_),
    .B1(_1760_),
    .X(_0206_));
 sky130_fd_sc_hd__and4_1 _3862_ (.A(_0274_),
    .B(\count[0] ),
    .C(\count[1] ),
    .D(\count[2] ),
    .X(_1761_));
 sky130_fd_sc_hd__o21a_1 _3863_ (.A1(net136),
    .A2(_1761_),
    .B1(_1759_),
    .X(_0205_));
 sky130_fd_sc_hd__a2bb2o_1 _3864_ (.A1_N(_1817_),
    .A2_N(_1924_),
    .B1(_0546_),
    .B2(_1922_),
    .X(_1762_));
 sky130_fd_sc_hd__a32o_1 _3865_ (.A1(_1801_),
    .A2(_1922_),
    .A3(_0835_),
    .B1(_1762_),
    .B2(\count[2] ),
    .X(_0204_));
 sky130_fd_sc_hd__o21a_1 _3866_ (.A1(_1817_),
    .A2(_1924_),
    .B1(\count[0] ),
    .X(_1763_));
 sky130_fd_sc_hd__o21a_1 _3867_ (.A1(\count[1] ),
    .A2(_1763_),
    .B1(_1762_),
    .X(_0203_));
 sky130_fd_sc_hd__o21ba_1 _3868_ (.A1(\count[0] ),
    .A2(_1924_),
    .B1_N(_1763_),
    .X(_0202_));
 sky130_fd_sc_hd__inv_2 _3869_ (.A(net65),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _3870_ (.A(net65),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _3871_ (.A(net65),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _3872_ (.A(net65),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _3873_ (.A(net65),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _3874_ (.A(net65),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _3875_ (.A(net141),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _3876_ (.A(net141),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _3877_ (.A(net141),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _3878_ (.A(net141),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _3879_ (.A(net141),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _3880_ (.A(net141),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _3881_ (.A(net141),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _3882_ (.A(net141),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _3883_ (.A(net141),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _3884_ (.A(net141),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _3885_ (.A(net141),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _3886_ (.A(net141),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _3887_ (.A(net141),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _3888_ (.A(net141),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _3889_ (.A(net141),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _3890_ (.A(net141),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _3891_ (.A(net141),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _3892_ (.A(net141),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _3893_ (.A(net141),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _3894_ (.A(net141),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _3895_ (.A(net141),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _3896_ (.A(net141),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _3897_ (.A(net141),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _3898_ (.A(net141),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _3899_ (.A(net141),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _3900_ (.A(net65),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _3901_ (.A(net65),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _3902_ (.A(net65),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _3903_ (.A(net65),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _3904_ (.A(net65),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _3905_ (.A(net65),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _3906_ (.A(net65),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _3907_ (.A(net141),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _3908_ (.A(net141),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _3909_ (.A(net141),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _3910_ (.A(net141),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _3911_ (.A(net141),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _3912_ (.A(net141),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _3913_ (.A(net141),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _3914_ (.A(net141),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _3915_ (.A(net141),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _3916_ (.A(net141),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _3917_ (.A(net141),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _3918_ (.A(net141),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _3919_ (.A(net141),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _3920_ (.A(net141),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _3921_ (.A(net141),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _3922_ (.A(net141),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _3923_ (.A(net141),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _3924_ (.A(net141),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _3925_ (.A(net141),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _3926_ (.A(net141),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _3927_ (.A(net141),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _3928_ (.A(net141),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _3929_ (.A(net141),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _3930_ (.A(net141),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _3931_ (.A(net141),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _3932_ (.A(net141),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _3933_ (.A(net141),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _3934_ (.A(net141),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _3935_ (.A(net141),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _3936_ (.A(net141),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _3937_ (.A(net65),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _3938_ (.A(net65),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _3939_ (.A(net65),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _3940_ (.A(net65),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _3941_ (.A(net65),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _3942_ (.A(net141),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _3943_ (.A(net141),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _3944_ (.A(net141),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _3945_ (.A(net141),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _3946_ (.A(net141),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _3947_ (.A(net141),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _3948_ (.A(net141),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _3949_ (.A(net141),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _3950_ (.A(net141),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _3951_ (.A(net141),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _3952_ (.A(net141),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _3953_ (.A(net141),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _3954_ (.A(net141),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _3955_ (.A(net141),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _3956_ (.A(net141),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _3957_ (.A(net141),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _3958_ (.A(net141),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _3959_ (.A(net141),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _3960_ (.A(net141),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _3961_ (.A(net141),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _3962_ (.A(net141),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _3963_ (.A(net141),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _3964_ (.A(net141),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _3965_ (.A(net141),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _3966_ (.A(net65),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _3967_ (.A(net65),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _3968_ (.A(net65),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _3969_ (.A(net65),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _3970_ (.A(net65),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _3971_ (.A(net65),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _3972_ (.A(net65),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _3973_ (.A(net65),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _3974_ (.A(net141),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _3975_ (.A(net141),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _3976_ (.A(net141),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _3977_ (.A(net141),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _3978_ (.A(net141),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _3979_ (.A(net141),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _3980_ (.A(net141),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _3981_ (.A(net141),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _3982_ (.A(net141),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _3983_ (.A(net65),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _3984_ (.A(net141),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _3985_ (.A(net141),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _3986_ (.A(net141),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _3987_ (.A(net141),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _3988_ (.A(net141),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _3989_ (.A(net141),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _3990_ (.A(net141),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _3991_ (.A(net141),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _3992_ (.A(net141),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _3993_ (.A(net141),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _3994_ (.A(net141),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _3995_ (.A(net141),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _3996_ (.A(net141),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _3997_ (.A(net141),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _3998_ (.A(net65),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _3999_ (.A(net141),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _4000_ (.A(net141),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _4001_ (.A(net141),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _4002_ (.A(net65),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _4003_ (.A(net65),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _4004_ (.A(net65),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _4005_ (.A(net65),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _4006_ (.A(net65),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _4007_ (.A(net65),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _4008_ (.A(net65),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _4009_ (.A(net65),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _4010_ (.A(net65),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _4011_ (.A(net65),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _4012_ (.A(net65),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _4013_ (.A(net65),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _4014_ (.A(net65),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _4015_ (.A(net65),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _4016_ (.A(net65),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _4017_ (.A(net65),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _4018_ (.A(net65),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _4019_ (.A(net65),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _4020_ (.A(net65),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _4021_ (.A(net65),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _4022_ (.A(net65),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _4023_ (.A(net65),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _4024_ (.A(net65),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _4025_ (.A(net65),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _4026_ (.A(net65),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _4027_ (.A(net65),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _4028_ (.A(net65),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _4029_ (.A(net65),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _4030_ (.A(net65),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _4031_ (.A(net65),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _4032_ (.A(net65),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _4033_ (.A(net65),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _4034_ (.A(net65),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _4035_ (.A(net65),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _4036_ (.A(net65),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _4037_ (.A(net65),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _4038_ (.A(net65),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _4039_ (.A(net141),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _4040_ (.A(net65),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _4041_ (.A(net65),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _4042_ (.A(net65),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _4043_ (.A(net65),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _4044_ (.A(net65),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _4045_ (.A(net65),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _4046_ (.A(net65),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _4047_ (.A(net65),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _4048_ (.A(net65),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _4049_ (.A(net65),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _4050_ (.A(net65),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _4051_ (.A(net65),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _4052_ (.A(net65),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _4053_ (.A(net65),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _4054_ (.A(net65),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _4055_ (.A(net65),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _4056_ (.A(net65),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _4057_ (.A(net65),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _4058_ (.A(net65),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _4059_ (.A(net65),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _4060_ (.A(net65),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _4061_ (.A(net65),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _4062_ (.A(net65),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _4063_ (.A(net65),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _4064_ (.A(net65),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _4065_ (.A(net65),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _4066_ (.A(net65),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _4067_ (.A(net65),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _4068_ (.A(net65),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _4069_ (.A(net65),
    .Y(_0201_));
 sky130_fd_sc_hd__dfrtp_4 _4070_ (.CLK(clknet_leaf_23_clk),
    .D(_0202_),
    .RESET_B(_0000_),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4071_ (.CLK(clknet_leaf_23_clk),
    .D(_0203_),
    .RESET_B(_0001_),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4072_ (.CLK(clknet_leaf_23_clk),
    .D(_0204_),
    .RESET_B(_0002_),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4073_ (.CLK(clknet_leaf_1_clk),
    .D(_0205_),
    .RESET_B(_0003_),
    .Q(\count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4074_ (.CLK(clknet_leaf_0_clk),
    .D(_0206_),
    .RESET_B(_0004_),
    .Q(\count[4] ));
 sky130_fd_sc_hd__dfrtp_4 _4075_ (.CLK(clknet_leaf_0_clk),
    .D(_0207_),
    .RESET_B(_0005_),
    .Q(\count[5] ));
 sky130_fd_sc_hd__dfrtp_4 _4076_ (.CLK(clknet_leaf_21_clk),
    .D(_0208_),
    .RESET_B(_0006_),
    .Q(sign));
 sky130_fd_sc_hd__dfrtp_1 _4077_ (.CLK(clknet_leaf_17_clk),
    .D(_0209_),
    .RESET_B(_0007_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _4078_ (.CLK(clknet_leaf_17_clk),
    .D(_0210_),
    .RESET_B(_0008_),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _4079_ (.CLK(clknet_leaf_17_clk),
    .D(_0211_),
    .RESET_B(_0009_),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _4080_ (.CLK(clknet_leaf_17_clk),
    .D(_0212_),
    .RESET_B(_0010_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _4081_ (.CLK(clknet_leaf_16_clk),
    .D(_0213_),
    .RESET_B(_0011_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_1 _4082_ (.CLK(clknet_leaf_16_clk),
    .D(_0214_),
    .RESET_B(_0012_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_1 _4083_ (.CLK(clknet_leaf_16_clk),
    .D(_0215_),
    .RESET_B(_0013_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_1 _4084_ (.CLK(clknet_leaf_16_clk),
    .D(_0216_),
    .RESET_B(_0014_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_1 _4085_ (.CLK(clknet_leaf_14_clk),
    .D(_0217_),
    .RESET_B(_0015_),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_1 _4086_ (.CLK(clknet_leaf_16_clk),
    .D(_0218_),
    .RESET_B(_0016_),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_1 _4087_ (.CLK(clknet_leaf_16_clk),
    .D(_0219_),
    .RESET_B(_0017_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _4088_ (.CLK(clknet_leaf_13_clk),
    .D(_0220_),
    .RESET_B(_0018_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _4089_ (.CLK(clknet_leaf_13_clk),
    .D(_0221_),
    .RESET_B(_0019_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _4090_ (.CLK(clknet_leaf_13_clk),
    .D(_0222_),
    .RESET_B(_0020_),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _4091_ (.CLK(clknet_leaf_13_clk),
    .D(_0223_),
    .RESET_B(_0021_),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _4092_ (.CLK(clknet_leaf_13_clk),
    .D(_0224_),
    .RESET_B(_0022_),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _4093_ (.CLK(clknet_leaf_12_clk),
    .D(_0225_),
    .RESET_B(_0023_),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _4094_ (.CLK(clknet_leaf_13_clk),
    .D(_0226_),
    .RESET_B(_0024_),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _4095_ (.CLK(clknet_leaf_12_clk),
    .D(_0227_),
    .RESET_B(_0025_),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _4096_ (.CLK(clknet_leaf_12_clk),
    .D(_0228_),
    .RESET_B(_0026_),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _4097_ (.CLK(clknet_leaf_12_clk),
    .D(_0229_),
    .RESET_B(_0027_),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _4098_ (.CLK(clknet_leaf_12_clk),
    .D(_0230_),
    .RESET_B(_0028_),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _4099_ (.CLK(clknet_leaf_12_clk),
    .D(_0231_),
    .RESET_B(_0029_),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _4100_ (.CLK(clknet_leaf_11_clk),
    .D(_0232_),
    .RESET_B(_0030_),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _4101_ (.CLK(clknet_leaf_5_clk),
    .D(_0233_),
    .RESET_B(_0031_),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _4102_ (.CLK(clknet_leaf_4_clk),
    .D(_0234_),
    .RESET_B(_0032_),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _4103_ (.CLK(clknet_leaf_3_clk),
    .D(_0235_),
    .RESET_B(_0033_),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _4104_ (.CLK(clknet_leaf_3_clk),
    .D(_0236_),
    .RESET_B(_0034_),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _4105_ (.CLK(clknet_leaf_3_clk),
    .D(_0237_),
    .RESET_B(_0035_),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _4106_ (.CLK(clknet_leaf_3_clk),
    .D(_0238_),
    .RESET_B(_0036_),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _4107_ (.CLK(clknet_leaf_3_clk),
    .D(_0239_),
    .RESET_B(_0037_),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _4108_ (.CLK(clknet_leaf_3_clk),
    .D(_0240_),
    .RESET_B(_0038_),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _4109_ (.CLK(clknet_leaf_10_clk),
    .D(_0241_),
    .RESET_B(_0039_),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _4110_ (.CLK(clknet_leaf_10_clk),
    .D(_0242_),
    .RESET_B(_0040_),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _4111_ (.CLK(clknet_leaf_11_clk),
    .D(_0243_),
    .RESET_B(_0041_),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _4112_ (.CLK(clknet_leaf_10_clk),
    .D(_0244_),
    .RESET_B(_0042_),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _4113_ (.CLK(clknet_leaf_11_clk),
    .D(_0245_),
    .RESET_B(_0043_),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _4114_ (.CLK(clknet_leaf_11_clk),
    .D(_0246_),
    .RESET_B(_0044_),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _4115_ (.CLK(clknet_leaf_11_clk),
    .D(_0247_),
    .RESET_B(_0045_),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _4116_ (.CLK(clknet_leaf_11_clk),
    .D(_0248_),
    .RESET_B(_0046_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _4117_ (.CLK(clknet_leaf_6_clk),
    .D(_0249_),
    .RESET_B(_0047_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _4118_ (.CLK(clknet_leaf_6_clk),
    .D(_0250_),
    .RESET_B(_0048_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _4119_ (.CLK(clknet_leaf_6_clk),
    .D(_0251_),
    .RESET_B(_0049_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _4120_ (.CLK(clknet_leaf_11_clk),
    .D(_0252_),
    .RESET_B(_0050_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _4121_ (.CLK(clknet_leaf_7_clk),
    .D(_0253_),
    .RESET_B(_0051_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _4122_ (.CLK(clknet_leaf_7_clk),
    .D(_0254_),
    .RESET_B(_0052_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_1 _4123_ (.CLK(clknet_leaf_7_clk),
    .D(_0255_),
    .RESET_B(_0053_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_1 _4124_ (.CLK(clknet_leaf_10_clk),
    .D(_0256_),
    .RESET_B(_0054_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_1 _4125_ (.CLK(clknet_leaf_10_clk),
    .D(_0257_),
    .RESET_B(_0055_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_1 _4126_ (.CLK(clknet_leaf_10_clk),
    .D(_0258_),
    .RESET_B(_0056_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_1 _4127_ (.CLK(clknet_leaf_10_clk),
    .D(_0259_),
    .RESET_B(_0057_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_1 _4128_ (.CLK(clknet_leaf_7_clk),
    .D(_0260_),
    .RESET_B(_0058_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_1 _4129_ (.CLK(clknet_leaf_7_clk),
    .D(_0261_),
    .RESET_B(_0059_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_1 _4130_ (.CLK(clknet_leaf_7_clk),
    .D(_0262_),
    .RESET_B(_0060_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_1 _4131_ (.CLK(clknet_leaf_6_clk),
    .D(_0263_),
    .RESET_B(_0061_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_1 _4132_ (.CLK(clknet_leaf_6_clk),
    .D(_0264_),
    .RESET_B(_0062_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_1 _4133_ (.CLK(clknet_leaf_6_clk),
    .D(_0265_),
    .RESET_B(_0063_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_1 _4134_ (.CLK(clknet_leaf_6_clk),
    .D(_0266_),
    .RESET_B(_0064_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 _4135_ (.CLK(clknet_leaf_5_clk),
    .D(_0267_),
    .RESET_B(_0065_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_1 _4136_ (.CLK(clknet_leaf_5_clk),
    .D(_0268_),
    .RESET_B(_0066_),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_1 _4137_ (.CLK(clknet_leaf_5_clk),
    .D(_0269_),
    .RESET_B(_0067_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_1 _4138_ (.CLK(clknet_leaf_5_clk),
    .D(_0270_),
    .RESET_B(_0068_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_1 _4139_ (.CLK(clknet_leaf_5_clk),
    .D(_0271_),
    .RESET_B(_0069_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_1 _4140_ (.CLK(clknet_leaf_5_clk),
    .D(_0272_),
    .RESET_B(_0070_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_1 _4141_ (.CLK(clknet_leaf_21_clk),
    .D(_0273_),
    .RESET_B(_0071_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_2 _4142_ (.CLK(clknet_leaf_21_clk),
    .D(_0274_),
    .RESET_B(_0072_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4143_ (.CLK(clknet_leaf_23_clk),
    .D(_0275_),
    .RESET_B(_0073_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4144_ (.CLK(clknet_leaf_17_clk),
    .D(_0276_),
    .RESET_B(_0074_),
    .Q(\acc[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4145_ (.CLK(clknet_leaf_17_clk),
    .D(_0277_),
    .RESET_B(_0075_),
    .Q(\acc[1] ));
 sky130_fd_sc_hd__dfrtp_4 _4146_ (.CLK(clknet_leaf_17_clk),
    .D(_0278_),
    .RESET_B(_0076_),
    .Q(\acc[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4147_ (.CLK(clknet_leaf_17_clk),
    .D(_0279_),
    .RESET_B(_0077_),
    .Q(\acc[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4148_ (.CLK(clknet_leaf_16_clk),
    .D(_0280_),
    .RESET_B(_0078_),
    .Q(\acc[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4149_ (.CLK(clknet_leaf_16_clk),
    .D(_0281_),
    .RESET_B(_0079_),
    .Q(\acc[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4150_ (.CLK(clknet_leaf_16_clk),
    .D(_0282_),
    .RESET_B(_0080_),
    .Q(\acc[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4151_ (.CLK(clknet_leaf_16_clk),
    .D(_0283_),
    .RESET_B(_0081_),
    .Q(\acc[7] ));
 sky130_fd_sc_hd__dfrtp_4 _4152_ (.CLK(clknet_leaf_16_clk),
    .D(_0284_),
    .RESET_B(_0082_),
    .Q(\acc[8] ));
 sky130_fd_sc_hd__dfrtp_4 _4153_ (.CLK(clknet_leaf_16_clk),
    .D(_0285_),
    .RESET_B(_0083_),
    .Q(\acc[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4154_ (.CLK(clknet_leaf_14_clk),
    .D(_0286_),
    .RESET_B(_0084_),
    .Q(\acc[10] ));
 sky130_fd_sc_hd__dfrtp_4 _4155_ (.CLK(clknet_leaf_14_clk),
    .D(_0287_),
    .RESET_B(_0085_),
    .Q(\acc[11] ));
 sky130_fd_sc_hd__dfrtp_4 _4156_ (.CLK(clknet_leaf_13_clk),
    .D(_0288_),
    .RESET_B(_0086_),
    .Q(\acc[12] ));
 sky130_fd_sc_hd__dfrtp_4 _4157_ (.CLK(clknet_leaf_13_clk),
    .D(_0289_),
    .RESET_B(_0087_),
    .Q(\acc[13] ));
 sky130_fd_sc_hd__dfrtp_2 _4158_ (.CLK(clknet_leaf_13_clk),
    .D(_0290_),
    .RESET_B(_0088_),
    .Q(\acc[14] ));
 sky130_fd_sc_hd__dfrtp_4 _4159_ (.CLK(clknet_leaf_15_clk),
    .D(_0291_),
    .RESET_B(_0089_),
    .Q(\acc[15] ));
 sky130_fd_sc_hd__dfrtp_4 _4160_ (.CLK(clknet_leaf_13_clk),
    .D(_0292_),
    .RESET_B(_0090_),
    .Q(\acc[16] ));
 sky130_fd_sc_hd__dfrtp_4 _4161_ (.CLK(clknet_leaf_13_clk),
    .D(_0293_),
    .RESET_B(_0091_),
    .Q(\acc[17] ));
 sky130_fd_sc_hd__dfrtp_4 _4162_ (.CLK(clknet_leaf_12_clk),
    .D(_0294_),
    .RESET_B(_0092_),
    .Q(\acc[18] ));
 sky130_fd_sc_hd__dfrtp_4 _4163_ (.CLK(clknet_leaf_12_clk),
    .D(_0295_),
    .RESET_B(_0093_),
    .Q(\acc[19] ));
 sky130_fd_sc_hd__dfrtp_4 _4164_ (.CLK(clknet_leaf_12_clk),
    .D(_0296_),
    .RESET_B(_0094_),
    .Q(\acc[20] ));
 sky130_fd_sc_hd__dfrtp_4 _4165_ (.CLK(clknet_leaf_11_clk),
    .D(_0297_),
    .RESET_B(_0095_),
    .Q(\acc[21] ));
 sky130_fd_sc_hd__dfrtp_4 _4166_ (.CLK(clknet_leaf_11_clk),
    .D(_0298_),
    .RESET_B(_0096_),
    .Q(\acc[22] ));
 sky130_fd_sc_hd__dfrtp_4 _4167_ (.CLK(clknet_leaf_11_clk),
    .D(_0299_),
    .RESET_B(_0097_),
    .Q(\acc[23] ));
 sky130_fd_sc_hd__dfrtp_4 _4168_ (.CLK(clknet_leaf_2_clk),
    .D(_0300_),
    .RESET_B(_0098_),
    .Q(\acc[24] ));
 sky130_fd_sc_hd__dfrtp_4 _4169_ (.CLK(clknet_leaf_2_clk),
    .D(_0301_),
    .RESET_B(_0099_),
    .Q(\acc[25] ));
 sky130_fd_sc_hd__dfrtp_4 _4170_ (.CLK(clknet_leaf_2_clk),
    .D(_0302_),
    .RESET_B(_0100_),
    .Q(\acc[26] ));
 sky130_fd_sc_hd__dfrtp_4 _4171_ (.CLK(clknet_leaf_2_clk),
    .D(_0303_),
    .RESET_B(_0101_),
    .Q(\acc[27] ));
 sky130_fd_sc_hd__dfrtp_4 _4172_ (.CLK(clknet_leaf_3_clk),
    .D(_0304_),
    .RESET_B(_0102_),
    .Q(\acc[28] ));
 sky130_fd_sc_hd__dfrtp_4 _4173_ (.CLK(clknet_leaf_0_clk),
    .D(_0305_),
    .RESET_B(_0103_),
    .Q(\acc[29] ));
 sky130_fd_sc_hd__dfrtp_4 _4174_ (.CLK(clknet_leaf_0_clk),
    .D(_0306_),
    .RESET_B(_0104_),
    .Q(\acc[30] ));
 sky130_fd_sc_hd__dfrtp_2 _4175_ (.CLK(clknet_leaf_3_clk),
    .D(_0307_),
    .RESET_B(_0105_),
    .Q(\acc[31] ));
 sky130_fd_sc_hd__dfrtp_4 _4176_ (.CLK(clknet_leaf_9_clk),
    .D(_0308_),
    .RESET_B(_0106_),
    .Q(\acc[32] ));
 sky130_fd_sc_hd__dfrtp_4 _4177_ (.CLK(clknet_leaf_11_clk),
    .D(_0309_),
    .RESET_B(_0107_),
    .Q(\acc[33] ));
 sky130_fd_sc_hd__dfrtp_4 _4178_ (.CLK(clknet_leaf_9_clk),
    .D(_0310_),
    .RESET_B(_0108_),
    .Q(\acc[34] ));
 sky130_fd_sc_hd__dfrtp_4 _4179_ (.CLK(clknet_leaf_9_clk),
    .D(_0311_),
    .RESET_B(_0109_),
    .Q(\acc[35] ));
 sky130_fd_sc_hd__dfrtp_4 _4180_ (.CLK(clknet_leaf_15_clk),
    .D(_0312_),
    .RESET_B(_0110_),
    .Q(\acc[36] ));
 sky130_fd_sc_hd__dfrtp_4 _4181_ (.CLK(clknet_leaf_15_clk),
    .D(_0313_),
    .RESET_B(_0111_),
    .Q(\acc[37] ));
 sky130_fd_sc_hd__dfrtp_4 _4182_ (.CLK(clknet_leaf_9_clk),
    .D(_0314_),
    .RESET_B(_0112_),
    .Q(\acc[38] ));
 sky130_fd_sc_hd__dfrtp_2 _4183_ (.CLK(clknet_leaf_15_clk),
    .D(_0315_),
    .RESET_B(_0113_),
    .Q(\acc[39] ));
 sky130_fd_sc_hd__dfrtp_4 _4184_ (.CLK(clknet_leaf_8_clk),
    .D(_0316_),
    .RESET_B(_0114_),
    .Q(\acc[40] ));
 sky130_fd_sc_hd__dfrtp_4 _4185_ (.CLK(clknet_leaf_2_clk),
    .D(_0317_),
    .RESET_B(_0115_),
    .Q(\acc[41] ));
 sky130_fd_sc_hd__dfrtp_4 _4186_ (.CLK(clknet_leaf_8_clk),
    .D(_0318_),
    .RESET_B(_0116_),
    .Q(\acc[42] ));
 sky130_fd_sc_hd__dfrtp_2 _4187_ (.CLK(clknet_leaf_8_clk),
    .D(_0319_),
    .RESET_B(_0117_),
    .Q(\acc[43] ));
 sky130_fd_sc_hd__dfrtp_4 _4188_ (.CLK(clknet_leaf_8_clk),
    .D(_0320_),
    .RESET_B(_0118_),
    .Q(\acc[44] ));
 sky130_fd_sc_hd__dfrtp_4 _4189_ (.CLK(clknet_leaf_8_clk),
    .D(_0321_),
    .RESET_B(_0119_),
    .Q(\acc[45] ));
 sky130_fd_sc_hd__dfrtp_4 _4190_ (.CLK(clknet_leaf_9_clk),
    .D(_0322_),
    .RESET_B(_0120_),
    .Q(\acc[46] ));
 sky130_fd_sc_hd__dfrtp_2 _4191_ (.CLK(clknet_leaf_15_clk),
    .D(_0323_),
    .RESET_B(_0121_),
    .Q(\acc[47] ));
 sky130_fd_sc_hd__dfrtp_4 _4192_ (.CLK(clknet_leaf_10_clk),
    .D(_0324_),
    .RESET_B(_0122_),
    .Q(\acc[48] ));
 sky130_fd_sc_hd__dfrtp_2 _4193_ (.CLK(clknet_leaf_10_clk),
    .D(_0325_),
    .RESET_B(_0123_),
    .Q(\acc[49] ));
 sky130_fd_sc_hd__dfrtp_4 _4194_ (.CLK(clknet_leaf_7_clk),
    .D(_0326_),
    .RESET_B(_0124_),
    .Q(\acc[50] ));
 sky130_fd_sc_hd__dfrtp_2 _4195_ (.CLK(clknet_leaf_7_clk),
    .D(_0327_),
    .RESET_B(_0125_),
    .Q(\acc[51] ));
 sky130_fd_sc_hd__dfrtp_4 _4196_ (.CLK(clknet_leaf_7_clk),
    .D(_0328_),
    .RESET_B(_0126_),
    .Q(\acc[52] ));
 sky130_fd_sc_hd__dfrtp_2 _4197_ (.CLK(clknet_leaf_6_clk),
    .D(_0329_),
    .RESET_B(_0127_),
    .Q(\acc[53] ));
 sky130_fd_sc_hd__dfrtp_2 _4198_ (.CLK(clknet_leaf_6_clk),
    .D(_0330_),
    .RESET_B(_0128_),
    .Q(\acc[54] ));
 sky130_fd_sc_hd__dfrtp_4 _4199_ (.CLK(clknet_leaf_8_clk),
    .D(_0331_),
    .RESET_B(_0129_),
    .Q(\acc[55] ));
 sky130_fd_sc_hd__dfrtp_4 _4200_ (.CLK(clknet_leaf_8_clk),
    .D(_0332_),
    .RESET_B(_0130_),
    .Q(\acc[56] ));
 sky130_fd_sc_hd__dfrtp_4 _4201_ (.CLK(clknet_leaf_6_clk),
    .D(_0333_),
    .RESET_B(_0131_),
    .Q(\acc[57] ));
 sky130_fd_sc_hd__dfrtp_4 _4202_ (.CLK(clknet_leaf_6_clk),
    .D(_0334_),
    .RESET_B(_0132_),
    .Q(\acc[58] ));
 sky130_fd_sc_hd__dfrtp_2 _4203_ (.CLK(clknet_leaf_4_clk),
    .D(_0335_),
    .RESET_B(_0133_),
    .Q(\acc[59] ));
 sky130_fd_sc_hd__dfrtp_4 _4204_ (.CLK(clknet_leaf_4_clk),
    .D(_0336_),
    .RESET_B(_0134_),
    .Q(\acc[60] ));
 sky130_fd_sc_hd__dfrtp_2 _4205_ (.CLK(clknet_leaf_4_clk),
    .D(_0337_),
    .RESET_B(_0135_),
    .Q(\acc[61] ));
 sky130_fd_sc_hd__dfrtp_4 _4206_ (.CLK(clknet_leaf_4_clk),
    .D(_0338_),
    .RESET_B(_0136_),
    .Q(\acc[62] ));
 sky130_fd_sc_hd__dfrtp_1 _4207_ (.CLK(clknet_leaf_3_clk),
    .D(_0339_),
    .RESET_B(_0137_),
    .Q(\acc[63] ));
 sky130_fd_sc_hd__dfrtp_4 _4208_ (.CLK(clknet_leaf_0_clk),
    .D(_0340_),
    .RESET_B(_0138_),
    .Q(\m[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4209_ (.CLK(clknet_leaf_0_clk),
    .D(_0341_),
    .RESET_B(_0139_),
    .Q(\m[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4210_ (.CLK(clknet_leaf_0_clk),
    .D(_0342_),
    .RESET_B(_0140_),
    .Q(\m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4211_ (.CLK(clknet_leaf_0_clk),
    .D(_0343_),
    .RESET_B(_0141_),
    .Q(\m[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4212_ (.CLK(clknet_leaf_0_clk),
    .D(_0344_),
    .RESET_B(_0142_),
    .Q(\m[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4213_ (.CLK(clknet_leaf_0_clk),
    .D(_0345_),
    .RESET_B(_0143_),
    .Q(\m[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4214_ (.CLK(clknet_leaf_23_clk),
    .D(_0346_),
    .RESET_B(_0144_),
    .Q(\m[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4215_ (.CLK(clknet_leaf_23_clk),
    .D(_0347_),
    .RESET_B(_0145_),
    .Q(\m[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4216_ (.CLK(clknet_leaf_23_clk),
    .D(_0348_),
    .RESET_B(_0146_),
    .Q(\m[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4217_ (.CLK(clknet_leaf_23_clk),
    .D(_0349_),
    .RESET_B(_0147_),
    .Q(\m[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4218_ (.CLK(clknet_leaf_23_clk),
    .D(_0350_),
    .RESET_B(_0148_),
    .Q(\m[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4219_ (.CLK(clknet_leaf_23_clk),
    .D(_0351_),
    .RESET_B(_0149_),
    .Q(\m[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4220_ (.CLK(clknet_leaf_23_clk),
    .D(_0352_),
    .RESET_B(_0150_),
    .Q(\m[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4221_ (.CLK(clknet_leaf_23_clk),
    .D(_0353_),
    .RESET_B(_0151_),
    .Q(\m[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4222_ (.CLK(clknet_leaf_23_clk),
    .D(_0354_),
    .RESET_B(_0152_),
    .Q(\m[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4223_ (.CLK(clknet_leaf_23_clk),
    .D(_0355_),
    .RESET_B(_0153_),
    .Q(\m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4224_ (.CLK(clknet_leaf_23_clk),
    .D(_0356_),
    .RESET_B(_0154_),
    .Q(\m[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4225_ (.CLK(clknet_leaf_23_clk),
    .D(_0357_),
    .RESET_B(_0155_),
    .Q(\m[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4226_ (.CLK(clknet_leaf_22_clk),
    .D(_0358_),
    .RESET_B(_0156_),
    .Q(\m[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4227_ (.CLK(clknet_leaf_22_clk),
    .D(_0359_),
    .RESET_B(_0157_),
    .Q(\m[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4228_ (.CLK(clknet_leaf_22_clk),
    .D(_0360_),
    .RESET_B(_0158_),
    .Q(\m[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4229_ (.CLK(clknet_leaf_22_clk),
    .D(_0361_),
    .RESET_B(_0159_),
    .Q(\m[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4230_ (.CLK(clknet_leaf_22_clk),
    .D(_0362_),
    .RESET_B(_0160_),
    .Q(\m[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4231_ (.CLK(clknet_leaf_22_clk),
    .D(_0363_),
    .RESET_B(_0161_),
    .Q(\m[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4232_ (.CLK(clknet_leaf_22_clk),
    .D(_0364_),
    .RESET_B(_0162_),
    .Q(\m[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4233_ (.CLK(clknet_leaf_22_clk),
    .D(_0365_),
    .RESET_B(_0163_),
    .Q(\m[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4234_ (.CLK(clknet_leaf_22_clk),
    .D(_0366_),
    .RESET_B(_0164_),
    .Q(\m[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4235_ (.CLK(clknet_leaf_22_clk),
    .D(_0367_),
    .RESET_B(_0165_),
    .Q(\m[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4236_ (.CLK(clknet_leaf_21_clk),
    .D(_0368_),
    .RESET_B(_0166_),
    .Q(\m[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4237_ (.CLK(clknet_leaf_21_clk),
    .D(_0369_),
    .RESET_B(_0167_),
    .Q(\m[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4238_ (.CLK(clknet_leaf_21_clk),
    .D(_0370_),
    .RESET_B(_0168_),
    .Q(\m[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4239_ (.CLK(clknet_leaf_21_clk),
    .D(_0371_),
    .RESET_B(_0169_),
    .Q(\m[31] ));
 sky130_fd_sc_hd__dfrtp_4 _4240_ (.CLK(clknet_leaf_18_clk),
    .D(_0372_),
    .RESET_B(_0170_),
    .Q(\q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _4241_ (.CLK(clknet_leaf_18_clk),
    .D(_0373_),
    .RESET_B(_0171_),
    .Q(\q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4242_ (.CLK(clknet_leaf_18_clk),
    .D(_0374_),
    .RESET_B(_0172_),
    .Q(\q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _4243_ (.CLK(clknet_leaf_18_clk),
    .D(_0375_),
    .RESET_B(_0173_),
    .Q(\q[3] ));
 sky130_fd_sc_hd__dfrtp_2 _4244_ (.CLK(clknet_leaf_18_clk),
    .D(_0376_),
    .RESET_B(_0174_),
    .Q(\q[4] ));
 sky130_fd_sc_hd__dfrtp_4 _4245_ (.CLK(clknet_leaf_18_clk),
    .D(_0377_),
    .RESET_B(_0175_),
    .Q(\q[5] ));
 sky130_fd_sc_hd__dfrtp_4 _4246_ (.CLK(clknet_leaf_19_clk),
    .D(_0378_),
    .RESET_B(_0176_),
    .Q(\q[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4247_ (.CLK(clknet_leaf_18_clk),
    .D(_0379_),
    .RESET_B(_0177_),
    .Q(\q[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4248_ (.CLK(clknet_leaf_19_clk),
    .D(_0380_),
    .RESET_B(_0178_),
    .Q(\q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4249_ (.CLK(clknet_leaf_18_clk),
    .D(_0381_),
    .RESET_B(_0179_),
    .Q(\q[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4250_ (.CLK(clknet_leaf_19_clk),
    .D(_0382_),
    .RESET_B(_0180_),
    .Q(\q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4251_ (.CLK(clknet_leaf_19_clk),
    .D(_0383_),
    .RESET_B(_0181_),
    .Q(\q[11] ));
 sky130_fd_sc_hd__dfrtp_2 _4252_ (.CLK(clknet_leaf_19_clk),
    .D(_0384_),
    .RESET_B(_0182_),
    .Q(\q[12] ));
 sky130_fd_sc_hd__dfrtp_2 _4253_ (.CLK(clknet_leaf_19_clk),
    .D(_0385_),
    .RESET_B(_0183_),
    .Q(\q[13] ));
 sky130_fd_sc_hd__dfrtp_2 _4254_ (.CLK(clknet_leaf_19_clk),
    .D(_0386_),
    .RESET_B(_0184_),
    .Q(\q[14] ));
 sky130_fd_sc_hd__dfrtp_2 _4255_ (.CLK(clknet_leaf_19_clk),
    .D(_0387_),
    .RESET_B(_0185_),
    .Q(\q[15] ));
 sky130_fd_sc_hd__dfrtp_4 _4256_ (.CLK(clknet_leaf_19_clk),
    .D(_0388_),
    .RESET_B(_0186_),
    .Q(\q[16] ));
 sky130_fd_sc_hd__dfrtp_4 _4257_ (.CLK(clknet_leaf_19_clk),
    .D(_0389_),
    .RESET_B(_0187_),
    .Q(\q[17] ));
 sky130_fd_sc_hd__dfrtp_2 _4258_ (.CLK(clknet_leaf_19_clk),
    .D(_0390_),
    .RESET_B(_0188_),
    .Q(\q[18] ));
 sky130_fd_sc_hd__dfrtp_2 _4259_ (.CLK(clknet_leaf_19_clk),
    .D(_0391_),
    .RESET_B(_0189_),
    .Q(\q[19] ));
 sky130_fd_sc_hd__dfrtp_2 _4260_ (.CLK(clknet_leaf_20_clk),
    .D(_0392_),
    .RESET_B(_0190_),
    .Q(\q[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4261_ (.CLK(clknet_leaf_20_clk),
    .D(_0393_),
    .RESET_B(_0191_),
    .Q(\q[21] ));
 sky130_fd_sc_hd__dfrtp_2 _4262_ (.CLK(clknet_leaf_20_clk),
    .D(_0394_),
    .RESET_B(_0192_),
    .Q(\q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4263_ (.CLK(clknet_leaf_20_clk),
    .D(_0395_),
    .RESET_B(_0193_),
    .Q(\q[23] ));
 sky130_fd_sc_hd__dfrtp_2 _4264_ (.CLK(clknet_leaf_20_clk),
    .D(_0396_),
    .RESET_B(_0194_),
    .Q(\q[24] ));
 sky130_fd_sc_hd__dfrtp_2 _4265_ (.CLK(clknet_leaf_20_clk),
    .D(_0397_),
    .RESET_B(_0195_),
    .Q(\q[25] ));
 sky130_fd_sc_hd__dfrtp_2 _4266_ (.CLK(clknet_leaf_20_clk),
    .D(_0398_),
    .RESET_B(_0196_),
    .Q(\q[26] ));
 sky130_fd_sc_hd__dfrtp_2 _4267_ (.CLK(clknet_leaf_21_clk),
    .D(_0399_),
    .RESET_B(_0197_),
    .Q(\q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4268_ (.CLK(clknet_leaf_1_clk),
    .D(_0400_),
    .RESET_B(_0198_),
    .Q(\q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4269_ (.CLK(clknet_leaf_0_clk),
    .D(_0401_),
    .RESET_B(_0199_),
    .Q(\q[29] ));
 sky130_fd_sc_hd__dfrtp_2 _4270_ (.CLK(clknet_leaf_20_clk),
    .D(_0402_),
    .RESET_B(_0200_),
    .Q(\q[30] ));
 sky130_fd_sc_hd__dfrtp_4 _4271_ (.CLK(clknet_leaf_21_clk),
    .D(_0403_),
    .RESET_B(_0201_),
    .Q(\q[31] ));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(multiplicand[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(multiplicand[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(multiplicand[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(multiplicand[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(multiplicand[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(multiplicand[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(multiplicand[15]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(multiplicand[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(multiplicand[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(multiplicand[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(multiplicand[19]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(multiplicand[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(multiplicand[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(multiplicand[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(multiplicand[22]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(multiplicand[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(multiplicand[24]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(multiplicand[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(multiplicand[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(multiplicand[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(multiplicand[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(multiplicand[29]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(multiplicand[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(multiplicand[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_16 input25 (.A(multiplicand[31]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(multiplicand[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(multiplicand[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(multiplicand[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(multiplicand[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(multiplicand[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(multiplicand[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(multiplicand[9]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(multiplier[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(multiplier[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(multiplier[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(multiplier[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(multiplier[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(multiplier[14]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(multiplier[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(multiplier[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(multiplier[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(multiplier[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(multiplier[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(multiplier[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(multiplier[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(multiplier[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(multiplier[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(multiplier[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(multiplier[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(multiplier[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(multiplier[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(multiplier[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(multiplier[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(multiplier[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(multiplier[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(multiplier[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_6 input57 (.A(multiplier[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(multiplier[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(multiplier[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(multiplier[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(multiplier[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(multiplier[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(multiplier[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(multiplier[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_16 input65 (.A(rst),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(start),
    .X(net66));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(done));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(product[0]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(product[10]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(product[11]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(product[12]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(product[13]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(product[14]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(product[15]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(product[16]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(product[17]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(product[18]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(product[19]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(product[1]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(product[20]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(product[21]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(product[22]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(product[23]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(product[24]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(product[25]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(product[26]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(product[27]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(product[28]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(product[29]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(product[2]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(product[30]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(product[31]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(product[32]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(product[33]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(product[34]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(product[35]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(product[36]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(product[37]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(product[38]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(product[39]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(product[3]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(product[40]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(product[41]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(product[42]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(product[43]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(product[44]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(product[45]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(product[46]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(product[47]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(product[48]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(product[49]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(product[4]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(product[50]));
 sky130_fd_sc_hd__buf_1 output114 (.A(net114),
    .X(product[51]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(product[52]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(product[53]));
 sky130_fd_sc_hd__buf_1 output117 (.A(net117),
    .X(product[54]));
 sky130_fd_sc_hd__buf_1 output118 (.A(net118),
    .X(product[55]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(product[56]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(product[57]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(product[58]));
 sky130_fd_sc_hd__buf_1 output122 (.A(net122),
    .X(product[59]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(product[5]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(product[60]));
 sky130_fd_sc_hd__buf_1 output125 (.A(net125),
    .X(product[61]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(product[62]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(product[63]));
 sky130_fd_sc_hd__buf_1 output128 (.A(net128),
    .X(product[6]));
 sky130_fd_sc_hd__buf_1 output129 (.A(net129),
    .X(product[7]));
 sky130_fd_sc_hd__buf_1 output130 (.A(net130),
    .X(product[8]));
 sky130_fd_sc_hd__buf_1 output131 (.A(net131),
    .X(product[9]));
 sky130_fd_sc_hd__buf_12 max_cap132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_8 max_cap133 (.A(_0437_),
    .X(net133));
 sky130_fd_sc_hd__buf_12 max_cap134 (.A(sign),
    .X(net134));
 sky130_fd_sc_hd__buf_12 max_cap135 (.A(\count[5] ),
    .X(net135));
 sky130_fd_sc_hd__buf_12 max_cap136 (.A(\count[3] ),
    .X(net136));
 sky130_fd_sc_hd__buf_12 max_cap137 (.A(\count[2] ),
    .X(net137));
 sky130_fd_sc_hd__buf_12 max_cap138 (.A(\count[1] ),
    .X(net138));
 sky130_fd_sc_hd__buf_12 max_cap139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_12 max_cap140 (.A(\count[0] ),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_16 max_cap141 (.A(net65),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_1_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_1_0__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__inv_12 clkload2 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__bufinv_16 clkload3 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__inv_6 clkload7 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkinv_4 clkload10 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload11 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_4 clkload12 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__bufinv_16 clkload13 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload14 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__bufinv_16 clkload15 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_4 clkload16 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload17 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload18 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload19 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__inv_6 clkload20 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_4 clkload21 (.A(clknet_leaf_15_clk));
endmodule
