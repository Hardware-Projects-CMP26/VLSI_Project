module dadda_multiplier_32 (product,
    signed_A,
    signed_B);
 output [63:0] product;
 input [31:0] signed_A;
 input [31:0] signed_B;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;

 sky130_fd_sc_hd__clkinv_16 _07585_ (.A(net1),
    .Y(_00288_));
 sky130_fd_sc_hd__clkinv_16 _07586_ (.A(net173),
    .Y(_00299_));
 sky130_fd_sc_hd__inv_16 _07587_ (.A(net33),
    .Y(_00310_));
 sky130_fd_sc_hd__clkinv_16 _07588_ (.A(net25),
    .Y(_00321_));
 sky130_fd_sc_hd__inv_2 _07589_ (.A(net55),
    .Y(_00332_));
 sky130_fd_sc_hd__inv_2 _07590_ (.A(net23),
    .Y(_00343_));
 sky130_fd_sc_hd__inv_2 _07591_ (.A(net58),
    .Y(_00354_));
 sky130_fd_sc_hd__inv_4 _07592_ (.A(net26),
    .Y(_00365_));
 sky130_fd_sc_hd__inv_8 _07593_ (.A(net59),
    .Y(_00376_));
 sky130_fd_sc_hd__inv_2 _07594_ (.A(net27),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_4 _07595_ (.A(net60),
    .Y(_00398_));
 sky130_fd_sc_hd__inv_2 _07596_ (.A(net28),
    .Y(_00408_));
 sky130_fd_sc_hd__inv_2 _07597_ (.A(net61),
    .Y(_00419_));
 sky130_fd_sc_hd__clkinv_4 _07598_ (.A(net29),
    .Y(_00430_));
 sky130_fd_sc_hd__clkinv_4 _07599_ (.A(net62),
    .Y(_00441_));
 sky130_fd_sc_hd__inv_2 _07600_ (.A(net30),
    .Y(_00452_));
 sky130_fd_sc_hd__inv_4 _07601_ (.A(net63),
    .Y(_00463_));
 sky130_fd_sc_hd__inv_2 _07602_ (.A(net64),
    .Y(_00474_));
 sky130_fd_sc_hd__inv_4 _07603_ (.A(net32),
    .Y(_00485_));
 sky130_fd_sc_hd__inv_2 _07604_ (.A(net2),
    .Y(_00496_));
 sky130_fd_sc_hd__inv_2 _07605_ (.A(net35),
    .Y(_00507_));
 sky130_fd_sc_hd__inv_2 _07606_ (.A(net3),
    .Y(_00518_));
 sky130_fd_sc_hd__inv_2 _07607_ (.A(net36),
    .Y(_00529_));
 sky130_fd_sc_hd__inv_4 _07608_ (.A(net4),
    .Y(_00540_));
 sky130_fd_sc_hd__inv_4 _07609_ (.A(net37),
    .Y(_00551_));
 sky130_fd_sc_hd__inv_2 _07610_ (.A(net5),
    .Y(_00561_));
 sky130_fd_sc_hd__clkinv_4 _07611_ (.A(net38),
    .Y(_00572_));
 sky130_fd_sc_hd__inv_2 _07612_ (.A(net39),
    .Y(_00583_));
 sky130_fd_sc_hd__inv_2 _07613_ (.A(net8),
    .Y(_00594_));
 sky130_fd_sc_hd__inv_2 _07614_ (.A(net9),
    .Y(_00605_));
 sky130_fd_sc_hd__inv_2 _07615_ (.A(net42),
    .Y(_00616_));
 sky130_fd_sc_hd__inv_2 _07616_ (.A(net10),
    .Y(_00627_));
 sky130_fd_sc_hd__inv_2 _07617_ (.A(net43),
    .Y(_00638_));
 sky130_fd_sc_hd__inv_2 _07618_ (.A(net11),
    .Y(_00649_));
 sky130_fd_sc_hd__inv_2 _07619_ (.A(net45),
    .Y(_00660_));
 sky130_fd_sc_hd__inv_2 _07620_ (.A(net13),
    .Y(_00671_));
 sky130_fd_sc_hd__inv_4 _07621_ (.A(net46),
    .Y(_00682_));
 sky130_fd_sc_hd__inv_2 _07622_ (.A(net14),
    .Y(_00693_));
 sky130_fd_sc_hd__inv_2 _07623_ (.A(net47),
    .Y(_00704_));
 sky130_fd_sc_hd__inv_2 _07624_ (.A(net15),
    .Y(_00715_));
 sky130_fd_sc_hd__inv_2 _07625_ (.A(net48),
    .Y(_00726_));
 sky130_fd_sc_hd__inv_2 _07626_ (.A(net51),
    .Y(_00736_));
 sky130_fd_sc_hd__inv_2 _07627_ (.A(net20),
    .Y(_00747_));
 sky130_fd_sc_hd__inv_2 _07628_ (.A(net53),
    .Y(_00758_));
 sky130_fd_sc_hd__inv_2 _07629_ (.A(net21),
    .Y(_00769_));
 sky130_fd_sc_hd__inv_2 _07630_ (.A(net54),
    .Y(_00780_));
 sky130_fd_sc_hd__inv_2 _07631_ (.A(net22),
    .Y(_00791_));
 sky130_fd_sc_hd__nor2_2 _07632_ (.A(_00288_),
    .B(_00310_),
    .Y(net65));
 sky130_fd_sc_hd__nor2_8 _07633_ (.A(net174),
    .B(_00299_),
    .Y(_00812_));
 sky130_fd_sc_hd__nor2_8 _07634_ (.A(net173),
    .B(_00321_),
    .Y(_00823_));
 sky130_fd_sc_hd__nor2_8 _07635_ (.A(_00812_),
    .B(_00823_),
    .Y(_00834_));
 sky130_fd_sc_hd__or2_4 _07636_ (.A(_00812_),
    .B(_00823_),
    .X(_00845_));
 sky130_fd_sc_hd__a21boi_4 _07637_ (.A1(net173),
    .A2(net33),
    .B1_N(net44),
    .Y(_00856_));
 sky130_fd_sc_hd__a21bo_2 _07638_ (.A1(net173),
    .A2(net33),
    .B1_N(net44),
    .X(_00867_));
 sky130_fd_sc_hd__and3b_4 _07639_ (.A_N(net44),
    .B(net173),
    .C(net33),
    .X(_00878_));
 sky130_fd_sc_hd__nand3b_4 _07640_ (.A_N(net44),
    .B(net173),
    .C(net33),
    .Y(_00889_));
 sky130_fd_sc_hd__nor2_8 _07641_ (.A(_00856_),
    .B(_00878_),
    .Y(_00900_));
 sky130_fd_sc_hd__nand2_8 _07642_ (.A(_00867_),
    .B(_00889_),
    .Y(_00911_));
 sky130_fd_sc_hd__a21boi_4 _07643_ (.A1(net1),
    .A2(net174),
    .B1_N(net12),
    .Y(_00921_));
 sky130_fd_sc_hd__a21bo_4 _07644_ (.A1(net1),
    .A2(net174),
    .B1_N(net12),
    .X(_00932_));
 sky130_fd_sc_hd__and3b_4 _07645_ (.A_N(net12),
    .B(net174),
    .C(net1),
    .X(_00943_));
 sky130_fd_sc_hd__nand3b_4 _07646_ (.A_N(net12),
    .B(net174),
    .C(net1),
    .Y(_00954_));
 sky130_fd_sc_hd__a21o_2 _07647_ (.A1(net1),
    .A2(net174),
    .B1(net12),
    .X(_00965_));
 sky130_fd_sc_hd__nand3_4 _07648_ (.A(net1),
    .B(net12),
    .C(net174),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_8 _07649_ (.A(_00965_),
    .B(_00976_),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_8 _07650_ (.A(_00932_),
    .B(_00954_),
    .Y(_00998_));
 sky130_fd_sc_hd__or4_2 _07651_ (.A(_00288_),
    .B(_00987_),
    .C(_00310_),
    .D(_00900_),
    .X(_01009_));
 sky130_fd_sc_hd__a32o_1 _07652_ (.A1(net33),
    .A2(_00965_),
    .A3(_00976_),
    .B1(_00911_),
    .B2(net1),
    .X(_01020_));
 sky130_fd_sc_hd__a22oi_1 _07653_ (.A1(net65),
    .A2(_00845_),
    .B1(_01009_),
    .B2(_01020_),
    .Y(_01031_));
 sky130_fd_sc_hd__and4_1 _07654_ (.A(_01009_),
    .B(net65),
    .C(_00845_),
    .D(_01020_),
    .X(_01042_));
 sky130_fd_sc_hd__nor2_1 _07655_ (.A(_01031_),
    .B(_01042_),
    .Y(net76));
 sky130_fd_sc_hd__o22a_1 _07656_ (.A1(_00812_),
    .A2(_00823_),
    .B1(net65),
    .B2(_01020_),
    .X(_01063_));
 sky130_fd_sc_hd__nor2_4 _07657_ (.A(net1),
    .B(net12),
    .Y(_01074_));
 sky130_fd_sc_hd__or2_1 _07658_ (.A(net1),
    .B(net12),
    .X(_01084_));
 sky130_fd_sc_hd__and3_4 _07659_ (.A(_01084_),
    .B(net174),
    .C(_00343_),
    .X(_01095_));
 sky130_fd_sc_hd__or3_4 _07660_ (.A(net23),
    .B(_01074_),
    .C(_00321_),
    .X(_01106_));
 sky130_fd_sc_hd__o21a_4 _07661_ (.A1(_00321_),
    .A2(_01074_),
    .B1(net23),
    .X(_01117_));
 sky130_fd_sc_hd__o21ai_4 _07662_ (.A1(_00321_),
    .A2(_01074_),
    .B1(net23),
    .Y(_01128_));
 sky130_fd_sc_hd__o21ai_4 _07663_ (.A1(net1),
    .A2(net12),
    .B1(net23),
    .Y(_01139_));
 sky130_fd_sc_hd__and3_2 _07664_ (.A(_01084_),
    .B(net23),
    .C(net174),
    .X(_01150_));
 sky130_fd_sc_hd__o21a_1 _07665_ (.A1(_00321_),
    .A2(_01074_),
    .B1(_00343_),
    .X(_01161_));
 sky130_fd_sc_hd__o21ai_4 _07666_ (.A1(_00321_),
    .A2(_01074_),
    .B1(_00343_),
    .Y(_01172_));
 sky130_fd_sc_hd__o21ai_4 _07667_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01172_),
    .Y(_01183_));
 sky130_fd_sc_hd__o21a_4 _07668_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01172_),
    .X(_01194_));
 sky130_fd_sc_hd__o211a_1 _07669_ (.A1(_00321_),
    .A2(_01139_),
    .B1(net33),
    .C1(_01172_),
    .X(_01205_));
 sky130_fd_sc_hd__nor2_8 _07670_ (.A(net44),
    .B(net33),
    .Y(_01216_));
 sky130_fd_sc_hd__o21ai_4 _07671_ (.A1(net44),
    .A2(net33),
    .B1(net173),
    .Y(_01227_));
 sky130_fd_sc_hd__o211a_4 _07672_ (.A1(net44),
    .A2(net33),
    .B1(net173),
    .C1(_00332_),
    .X(_01238_));
 sky130_fd_sc_hd__o21a_4 _07673_ (.A1(_00299_),
    .A2(_01216_),
    .B1(net55),
    .X(_01249_));
 sky130_fd_sc_hd__o21ai_1 _07674_ (.A1(net44),
    .A2(net33),
    .B1(net55),
    .Y(_01259_));
 sky130_fd_sc_hd__o211ai_4 _07675_ (.A1(net44),
    .A2(net33),
    .B1(net55),
    .C1(net173),
    .Y(_01270_));
 sky130_fd_sc_hd__o21ai_4 _07676_ (.A1(_00299_),
    .A2(_01216_),
    .B1(_00332_),
    .Y(_01281_));
 sky130_fd_sc_hd__nand2_8 _07677_ (.A(_01270_),
    .B(_01281_),
    .Y(_01292_));
 sky130_fd_sc_hd__o21a_4 _07678_ (.A1(_00299_),
    .A2(_01259_),
    .B1(_01281_),
    .X(_01303_));
 sky130_fd_sc_hd__nand3_2 _07679_ (.A(_01281_),
    .B(net1),
    .C(_01270_),
    .Y(_01314_));
 sky130_fd_sc_hd__and4_1 _07680_ (.A(_00911_),
    .B(_00998_),
    .C(_01303_),
    .D(net1),
    .X(_01325_));
 sky130_fd_sc_hd__o22a_1 _07681_ (.A1(_00900_),
    .A2(_00987_),
    .B1(_00288_),
    .B2(_01292_),
    .X(_01336_));
 sky130_fd_sc_hd__or4_1 _07682_ (.A(_00310_),
    .B(_01183_),
    .C(_01325_),
    .D(_01336_),
    .X(_01347_));
 sky130_fd_sc_hd__a2bb2o_1 _07683_ (.A1_N(_01325_),
    .A2_N(_01336_),
    .B1(net33),
    .B2(_01194_),
    .X(_01358_));
 sky130_fd_sc_hd__nand2_1 _07684_ (.A(_01347_),
    .B(_01358_),
    .Y(_01369_));
 sky130_fd_sc_hd__xor2_2 _07685_ (.A(_01009_),
    .B(_01369_),
    .X(_01380_));
 sky130_fd_sc_hd__xor2_1 _07686_ (.A(_01063_),
    .B(_01380_),
    .X(net87));
 sky130_fd_sc_hd__or3_1 _07687_ (.A(net65),
    .B(_01020_),
    .C(_01380_),
    .X(_01401_));
 sky130_fd_sc_hd__nor3_4 _07688_ (.A(net1),
    .B(net12),
    .C(net23),
    .Y(_01412_));
 sky130_fd_sc_hd__o311a_4 _07689_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .B1(_00365_),
    .C1(net174),
    .X(_01423_));
 sky130_fd_sc_hd__o311ai_4 _07690_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .B1(_00365_),
    .C1(net174),
    .Y(_01434_));
 sky130_fd_sc_hd__o21a_4 _07691_ (.A1(_00321_),
    .A2(_01412_),
    .B1(net26),
    .X(_01445_));
 sky130_fd_sc_hd__o21ai_4 _07692_ (.A1(_00321_),
    .A2(_01412_),
    .B1(net26),
    .Y(_01455_));
 sky130_fd_sc_hd__o311ai_4 _07693_ (.A1(net1),
    .A2(net12),
    .A3(net23),
    .B1(net26),
    .C1(net174),
    .Y(_01466_));
 sky130_fd_sc_hd__o21ai_4 _07694_ (.A1(_00321_),
    .A2(_01412_),
    .B1(_00365_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_8 _07695_ (.A(_01466_),
    .B(_01477_),
    .Y(_01488_));
 sky130_fd_sc_hd__nand2_8 _07696_ (.A(_01434_),
    .B(_01455_),
    .Y(_01499_));
 sky130_fd_sc_hd__o21ai_1 _07697_ (.A1(_01423_),
    .A2(_01445_),
    .B1(net33),
    .Y(_01510_));
 sky130_fd_sc_hd__nand2_1 _07698_ (.A(net173),
    .B(net55),
    .Y(_01521_));
 sky130_fd_sc_hd__and3_4 _07699_ (.A(_01227_),
    .B(_01521_),
    .C(net58),
    .X(_01532_));
 sky130_fd_sc_hd__nand3_4 _07700_ (.A(_01227_),
    .B(_01521_),
    .C(net58),
    .Y(_01543_));
 sky130_fd_sc_hd__o311a_4 _07701_ (.A1(net44),
    .A2(net33),
    .A3(net55),
    .B1(_00354_),
    .C1(net173),
    .X(_01554_));
 sky130_fd_sc_hd__o311ai_4 _07702_ (.A1(net44),
    .A2(net33),
    .A3(net55),
    .B1(_00354_),
    .C1(net173),
    .Y(_01565_));
 sky130_fd_sc_hd__o311a_4 _07703_ (.A1(net44),
    .A2(net33),
    .A3(net55),
    .B1(net58),
    .C1(net173),
    .X(_01576_));
 sky130_fd_sc_hd__o311ai_4 _07704_ (.A1(net44),
    .A2(net33),
    .A3(net55),
    .B1(net58),
    .C1(net173),
    .Y(_01587_));
 sky130_fd_sc_hd__and3_4 _07705_ (.A(_00354_),
    .B(_01227_),
    .C(_01521_),
    .X(_01598_));
 sky130_fd_sc_hd__o211ai_4 _07706_ (.A1(_00299_),
    .A2(_00332_),
    .B1(_00354_),
    .C1(_01227_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_8 _07707_ (.A(_01587_),
    .B(_01609_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_8 _07708_ (.A(_01543_),
    .B(_01565_),
    .Y(_01631_));
 sky130_fd_sc_hd__a22o_1 _07709_ (.A1(_00932_),
    .A2(_00954_),
    .B1(_01543_),
    .B2(_01565_),
    .X(_01642_));
 sky130_fd_sc_hd__nor2_2 _07710_ (.A(_01314_),
    .B(_01642_),
    .Y(_01652_));
 sky130_fd_sc_hd__or4_1 _07711_ (.A(_00987_),
    .B(_01576_),
    .C(_01598_),
    .D(_01314_),
    .X(_01663_));
 sky130_fd_sc_hd__o32a_1 _07712_ (.A1(_00288_),
    .A2(_01576_),
    .A3(_01598_),
    .B1(_00987_),
    .B2(_01292_),
    .X(_01674_));
 sky130_fd_sc_hd__a32o_1 _07713_ (.A1(_00998_),
    .A2(_01270_),
    .A3(_01281_),
    .B1(_01631_),
    .B2(net1),
    .X(_01685_));
 sky130_fd_sc_hd__o22ai_4 _07714_ (.A1(_00900_),
    .A2(_01183_),
    .B1(_01652_),
    .B2(_01674_),
    .Y(_01696_));
 sky130_fd_sc_hd__inv_2 _07715_ (.A(_01696_),
    .Y(_01707_));
 sky130_fd_sc_hd__and4_1 _07716_ (.A(_00911_),
    .B(_01194_),
    .C(_01663_),
    .D(_01685_),
    .X(_01718_));
 sky130_fd_sc_hd__o2111ai_2 _07717_ (.A1(_01314_),
    .A2(_01642_),
    .B1(_01685_),
    .C1(_01194_),
    .D1(_00911_),
    .Y(_01729_));
 sky130_fd_sc_hd__a21oi_1 _07718_ (.A1(_01696_),
    .A2(_01729_),
    .B1(_01510_),
    .Y(_01740_));
 sky130_fd_sc_hd__o211a_1 _07719_ (.A1(_01488_),
    .A2(_00310_),
    .B1(_01729_),
    .C1(_01696_),
    .X(_01751_));
 sky130_fd_sc_hd__o21a_1 _07720_ (.A1(_01740_),
    .A2(_01751_),
    .B1(_01325_),
    .X(_01762_));
 sky130_fd_sc_hd__nor3_1 _07721_ (.A(_01325_),
    .B(_01740_),
    .C(_01751_),
    .Y(_01773_));
 sky130_fd_sc_hd__nor2_1 _07722_ (.A(_01762_),
    .B(_01773_),
    .Y(_01784_));
 sky130_fd_sc_hd__o2111ai_1 _07723_ (.A1(_01314_),
    .A2(_01205_),
    .B1(_00911_),
    .C1(net65),
    .D1(_00998_),
    .Y(_01795_));
 sky130_fd_sc_hd__o41a_1 _07724_ (.A1(_00310_),
    .A2(_01183_),
    .A3(_01325_),
    .A4(_01336_),
    .B1(_01795_),
    .X(_01806_));
 sky130_fd_sc_hd__xnor2_1 _07725_ (.A(_01784_),
    .B(_01806_),
    .Y(_01817_));
 sky130_fd_sc_hd__o311a_1 _07726_ (.A1(net65),
    .A2(_01020_),
    .A3(_01380_),
    .B1(_01817_),
    .C1(_00845_),
    .X(_01828_));
 sky130_fd_sc_hd__a21oi_1 _07727_ (.A1(_00845_),
    .A2(_01401_),
    .B1(_01817_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _07728_ (.A(_01828_),
    .B(_01839_),
    .Y(net98));
 sky130_fd_sc_hd__or4_2 _07729_ (.A(net65),
    .B(_01020_),
    .C(_01380_),
    .D(_01817_),
    .X(_01860_));
 sky130_fd_sc_hd__nor4_2 _07730_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(net26),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _07731_ (.A(_01412_),
    .B(_00365_),
    .Y(_01881_));
 sky130_fd_sc_hd__o311a_4 _07732_ (.A1(net23),
    .A2(net26),
    .A3(_01084_),
    .B1(_00387_),
    .C1(net174),
    .X(_01892_));
 sky130_fd_sc_hd__a311o_4 _07733_ (.A1(_00343_),
    .A2(_01074_),
    .A3(_00365_),
    .B1(_00321_),
    .C1(net27),
    .X(_01903_));
 sky130_fd_sc_hd__o21a_4 _07734_ (.A1(_00321_),
    .A2(net171),
    .B1(net27),
    .X(_01914_));
 sky130_fd_sc_hd__o21ai_4 _07735_ (.A1(_00321_),
    .A2(net171),
    .B1(net27),
    .Y(_01925_));
 sky130_fd_sc_hd__nand3_4 _07736_ (.A(_01881_),
    .B(net27),
    .C(net174),
    .Y(_01936_));
 sky130_fd_sc_hd__o21ai_4 _07737_ (.A1(_00321_),
    .A2(_01870_),
    .B1(_00387_),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_8 _07738_ (.A(_01936_),
    .B(_01947_),
    .Y(_01958_));
 sky130_fd_sc_hd__nand2_8 _07739_ (.A(_01903_),
    .B(_01925_),
    .Y(_01969_));
 sky130_fd_sc_hd__and3_1 _07740_ (.A(_00911_),
    .B(_01466_),
    .C(_01477_),
    .X(_01980_));
 sky130_fd_sc_hd__o221a_1 _07741_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01238_),
    .B2(_01249_),
    .C1(_01172_),
    .X(_01991_));
 sky130_fd_sc_hd__nor2_8 _07742_ (.A(net55),
    .B(net58),
    .Y(_02002_));
 sky130_fd_sc_hd__nor4_4 _07743_ (.A(net44),
    .B(net33),
    .C(net55),
    .D(net58),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_4 _07744_ (.A(_01216_),
    .B(_02002_),
    .Y(_02024_));
 sky130_fd_sc_hd__a311oi_1 _07745_ (.A1(_00332_),
    .A2(_01216_),
    .A3(_00354_),
    .B1(_00299_),
    .C1(net59),
    .Y(_02035_));
 sky130_fd_sc_hd__a211o_4 _07746_ (.A1(_01216_),
    .A2(_02002_),
    .B1(_00299_),
    .C1(net59),
    .X(_02046_));
 sky130_fd_sc_hd__a21oi_4 _07747_ (.A1(_02024_),
    .A2(net173),
    .B1(_00376_),
    .Y(_02057_));
 sky130_fd_sc_hd__o21bai_4 _07748_ (.A1(_00299_),
    .A2(_02013_),
    .B1_N(_00376_),
    .Y(_02068_));
 sky130_fd_sc_hd__a211oi_4 _07749_ (.A1(_01216_),
    .A2(_02002_),
    .B1(_00299_),
    .C1(_00376_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand3_4 _07750_ (.A(_02024_),
    .B(net59),
    .C(net173),
    .Y(_02089_));
 sky130_fd_sc_hd__a21oi_4 _07751_ (.A1(_02024_),
    .A2(net173),
    .B1(net59),
    .Y(_02100_));
 sky130_fd_sc_hd__o21bai_4 _07752_ (.A1(_00299_),
    .A2(_02013_),
    .B1_N(net59),
    .Y(_02111_));
 sky130_fd_sc_hd__nand2_8 _07753_ (.A(_02089_),
    .B(_02111_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_8 _07754_ (.A(_02046_),
    .B(_02068_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand3_1 _07755_ (.A(_02111_),
    .B(net1),
    .C(_02089_),
    .Y(_02144_));
 sky130_fd_sc_hd__a32oi_4 _07756_ (.A1(_02111_),
    .A2(net1),
    .A3(_02089_),
    .B1(_00998_),
    .B2(_01631_),
    .Y(_02155_));
 sky130_fd_sc_hd__o21ai_2 _07757_ (.A1(_00987_),
    .A2(_01620_),
    .B1(_02144_),
    .Y(_02166_));
 sky130_fd_sc_hd__and3_4 _07758_ (.A(_00965_),
    .B(_00976_),
    .C(net1),
    .X(_02177_));
 sky130_fd_sc_hd__o21ai_4 _07759_ (.A1(net172),
    .A2(_00943_),
    .B1(net1),
    .Y(_02188_));
 sky130_fd_sc_hd__and3_2 _07760_ (.A(_01631_),
    .B(_02089_),
    .C(_02111_),
    .X(_02199_));
 sky130_fd_sc_hd__a22o_4 _07761_ (.A1(_01543_),
    .A2(_01565_),
    .B1(_02046_),
    .B2(_02068_),
    .X(_02210_));
 sky130_fd_sc_hd__and4_2 _07762_ (.A(_02177_),
    .B(_02111_),
    .C(_02089_),
    .D(_01631_),
    .X(_02221_));
 sky130_fd_sc_hd__nand4_2 _07763_ (.A(_02177_),
    .B(_02111_),
    .C(_02089_),
    .D(_01631_),
    .Y(_02232_));
 sky130_fd_sc_hd__a22oi_1 _07764_ (.A1(_01194_),
    .A2(_01303_),
    .B1(_02166_),
    .B2(_02232_),
    .Y(_02243_));
 sky130_fd_sc_hd__o22ai_4 _07765_ (.A1(_01183_),
    .A2(_01292_),
    .B1(_02155_),
    .B2(_02221_),
    .Y(_02254_));
 sky130_fd_sc_hd__o311a_1 _07766_ (.A1(_01620_),
    .A2(_02188_),
    .A3(_02122_),
    .B1(_01991_),
    .C1(_02166_),
    .X(_02265_));
 sky130_fd_sc_hd__o2111ai_2 _07767_ (.A1(_02188_),
    .A2(_02210_),
    .B1(_01194_),
    .C1(_01303_),
    .D1(_02166_),
    .Y(_02276_));
 sky130_fd_sc_hd__o2111ai_2 _07768_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_01499_),
    .C1(_02254_),
    .D1(_02276_),
    .Y(_02287_));
 sky130_fd_sc_hd__o22ai_1 _07769_ (.A1(_00900_),
    .A2(_01488_),
    .B1(_02243_),
    .B2(_02265_),
    .Y(_02298_));
 sky130_fd_sc_hd__o21ai_1 _07770_ (.A1(_02243_),
    .A2(_02265_),
    .B1(_01980_),
    .Y(_02309_));
 sky130_fd_sc_hd__o211ai_1 _07771_ (.A1(_00900_),
    .A2(_01488_),
    .B1(_02254_),
    .C1(_02276_),
    .Y(_02320_));
 sky130_fd_sc_hd__nand3_2 _07772_ (.A(_02287_),
    .B(_02298_),
    .C(_01652_),
    .Y(_02331_));
 sky130_fd_sc_hd__and3_1 _07773_ (.A(_01663_),
    .B(_02309_),
    .C(_02320_),
    .X(_02342_));
 sky130_fd_sc_hd__nand3_1 _07774_ (.A(_01663_),
    .B(_02309_),
    .C(_02320_),
    .Y(_02352_));
 sky130_fd_sc_hd__and4_1 _07775_ (.A(_01969_),
    .B(_02331_),
    .C(_02352_),
    .D(net33),
    .X(_02363_));
 sky130_fd_sc_hd__nand4_2 _07776_ (.A(_01969_),
    .B(_02331_),
    .C(_02352_),
    .D(net33),
    .Y(_02374_));
 sky130_fd_sc_hd__o2bb2ai_2 _07777_ (.A1_N(_02331_),
    .A2_N(_02352_),
    .B1(_00310_),
    .B2(_01958_),
    .Y(_02385_));
 sky130_fd_sc_hd__o41a_1 _07778_ (.A1(_00900_),
    .A2(_01183_),
    .A3(_01652_),
    .A4(_01674_),
    .B1(_01510_),
    .X(_02396_));
 sky130_fd_sc_hd__and3_1 _07779_ (.A(_01696_),
    .B(net33),
    .C(_01499_),
    .X(_02407_));
 sky130_fd_sc_hd__a31o_1 _07780_ (.A1(_01696_),
    .A2(net33),
    .A3(_01499_),
    .B1(_01718_),
    .X(_02418_));
 sky130_fd_sc_hd__a21oi_1 _07781_ (.A1(_02374_),
    .A2(_02385_),
    .B1(_02418_),
    .Y(_02429_));
 sky130_fd_sc_hd__o2bb2ai_1 _07782_ (.A1_N(_02374_),
    .A2_N(_02385_),
    .B1(_02396_),
    .B2(_01707_),
    .Y(_02440_));
 sky130_fd_sc_hd__o21bai_2 _07783_ (.A1(_01773_),
    .A2(_01806_),
    .B1_N(_01762_),
    .Y(_02451_));
 sky130_fd_sc_hd__o21ai_1 _07784_ (.A1(_01718_),
    .A2(_02407_),
    .B1(_02385_),
    .Y(_02462_));
 sky130_fd_sc_hd__and3_1 _07785_ (.A(_02374_),
    .B(_02385_),
    .C(_02418_),
    .X(_02473_));
 sky130_fd_sc_hd__a31oi_2 _07786_ (.A1(_02374_),
    .A2(_02385_),
    .A3(_02418_),
    .B1(_02451_),
    .Y(_02484_));
 sky130_fd_sc_hd__o21ai_1 _07787_ (.A1(_02429_),
    .A2(_02473_),
    .B1(_02451_),
    .Y(_02495_));
 sky130_fd_sc_hd__a21bo_1 _07788_ (.A1(_02440_),
    .A2(_02484_),
    .B1_N(_02495_),
    .X(_02506_));
 sky130_fd_sc_hd__a21oi_1 _07789_ (.A1(_00845_),
    .A2(_01860_),
    .B1(_02506_),
    .Y(_02517_));
 sky130_fd_sc_hd__and3_1 _07790_ (.A(_00845_),
    .B(_01860_),
    .C(_02506_),
    .X(_02528_));
 sky130_fd_sc_hd__nor2_1 _07791_ (.A(_02517_),
    .B(_02528_),
    .Y(net109));
 sky130_fd_sc_hd__o21ai_1 _07792_ (.A1(_01860_),
    .A2(_02506_),
    .B1(_00845_),
    .Y(_02549_));
 sky130_fd_sc_hd__o21a_1 _07793_ (.A1(_00310_),
    .A2(_01958_),
    .B1(_02331_),
    .X(_02560_));
 sky130_fd_sc_hd__nor2_1 _07794_ (.A(_02342_),
    .B(_02560_),
    .Y(_02571_));
 sky130_fd_sc_hd__nand4_1 _07795_ (.A(_01074_),
    .B(_00387_),
    .C(_00365_),
    .D(_00343_),
    .Y(_02581_));
 sky130_fd_sc_hd__a311o_4 _07796_ (.A1(_01412_),
    .A2(_00387_),
    .A3(_00365_),
    .B1(_00321_),
    .C1(net28),
    .X(_02592_));
 sky130_fd_sc_hd__a21o_2 _07797_ (.A1(_02581_),
    .A2(net174),
    .B1(_00408_),
    .X(_02603_));
 sky130_fd_sc_hd__a311o_4 _07798_ (.A1(_01412_),
    .A2(_00387_),
    .A3(_00365_),
    .B1(_00321_),
    .C1(_00408_),
    .X(_02614_));
 sky130_fd_sc_hd__a21o_4 _07799_ (.A1(_02581_),
    .A2(net174),
    .B1(net28),
    .X(_02625_));
 sky130_fd_sc_hd__nand2_8 _07800_ (.A(_02614_),
    .B(_02625_),
    .Y(_02636_));
 sky130_fd_sc_hd__nand2_8 _07801_ (.A(_02592_),
    .B(_02603_),
    .Y(_02647_));
 sky130_fd_sc_hd__a21o_1 _07802_ (.A1(_02592_),
    .A2(_02603_),
    .B1(_00310_),
    .X(_02658_));
 sky130_fd_sc_hd__a31o_1 _07803_ (.A1(_02166_),
    .A2(_02232_),
    .A3(_01991_),
    .B1(_01980_),
    .X(_02669_));
 sky130_fd_sc_hd__and3_1 _07804_ (.A(_00911_),
    .B(_01499_),
    .C(_02254_),
    .X(_02680_));
 sky130_fd_sc_hd__a31o_1 _07805_ (.A1(_00911_),
    .A2(_01499_),
    .A3(_02254_),
    .B1(_02265_),
    .X(_02691_));
 sky130_fd_sc_hd__a32oi_4 _07806_ (.A1(_00911_),
    .A2(_01936_),
    .A3(_01947_),
    .B1(_01303_),
    .B2(_01499_),
    .Y(_02702_));
 sky130_fd_sc_hd__nor4_4 _07807_ (.A(_00900_),
    .B(_01292_),
    .C(_01488_),
    .D(_01958_),
    .Y(_02713_));
 sky130_fd_sc_hd__a31oi_2 _07808_ (.A1(_01303_),
    .A2(_01969_),
    .A3(_01980_),
    .B1(_02702_),
    .Y(_02724_));
 sky130_fd_sc_hd__o221a_1 _07809_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01532_),
    .B2(_01554_),
    .C1(_01172_),
    .X(_02735_));
 sky130_fd_sc_hd__o211ai_2 _07810_ (.A1(_00921_),
    .A2(_00943_),
    .B1(_02089_),
    .C1(_02111_),
    .Y(_02746_));
 sky130_fd_sc_hd__nand3_4 _07811_ (.A(_01216_),
    .B(_02002_),
    .C(_00376_),
    .Y(_02757_));
 sky130_fd_sc_hd__a31oi_1 _07812_ (.A1(_01216_),
    .A2(_02002_),
    .A3(_00376_),
    .B1(_00299_),
    .Y(_02768_));
 sky130_fd_sc_hd__a31o_2 _07813_ (.A1(_01216_),
    .A2(_02002_),
    .A3(_00376_),
    .B1(_00299_),
    .X(_02779_));
 sky130_fd_sc_hd__a311oi_4 _07814_ (.A1(_01216_),
    .A2(_02002_),
    .A3(_00376_),
    .B1(net60),
    .C1(_00299_),
    .Y(_02790_));
 sky130_fd_sc_hd__a21oi_4 _07815_ (.A1(_02757_),
    .A2(net173),
    .B1(_00398_),
    .Y(_02800_));
 sky130_fd_sc_hd__a311oi_4 _07816_ (.A1(_01216_),
    .A2(_02002_),
    .A3(_00376_),
    .B1(_00398_),
    .C1(_00299_),
    .Y(_02811_));
 sky130_fd_sc_hd__o211ai_4 _07817_ (.A1(net59),
    .A2(_02024_),
    .B1(net60),
    .C1(net173),
    .Y(_02822_));
 sky130_fd_sc_hd__a21oi_4 _07818_ (.A1(_02757_),
    .A2(net173),
    .B1(net60),
    .Y(_02833_));
 sky130_fd_sc_hd__a21o_1 _07819_ (.A1(_02757_),
    .A2(net173),
    .B1(net60),
    .X(_02844_));
 sky130_fd_sc_hd__nor2_4 _07820_ (.A(net169),
    .B(_02800_),
    .Y(_02855_));
 sky130_fd_sc_hd__nor2_8 _07821_ (.A(_02811_),
    .B(_02833_),
    .Y(_02866_));
 sky130_fd_sc_hd__o21ai_2 _07822_ (.A1(net60),
    .A2(_02768_),
    .B1(net1),
    .Y(_02877_));
 sky130_fd_sc_hd__nand3_1 _07823_ (.A(_02844_),
    .B(net1),
    .C(_02822_),
    .Y(_02888_));
 sky130_fd_sc_hd__and3_2 _07824_ (.A(_02133_),
    .B(_02822_),
    .C(_02844_),
    .X(_02899_));
 sky130_fd_sc_hd__o2bb2ai_4 _07825_ (.A1_N(_02046_),
    .A2_N(_02068_),
    .B1(net169),
    .B2(_02800_),
    .Y(_02910_));
 sky130_fd_sc_hd__o32a_1 _07826_ (.A1(_00987_),
    .A2(_02079_),
    .A3(_02100_),
    .B1(net167),
    .B2(_02877_),
    .X(_02921_));
 sky130_fd_sc_hd__o32ai_4 _07827_ (.A1(_00987_),
    .A2(_02079_),
    .A3(_02100_),
    .B1(net167),
    .B2(_02877_),
    .Y(_02932_));
 sky130_fd_sc_hd__o21ai_2 _07828_ (.A1(_02188_),
    .A2(_02910_),
    .B1(_02932_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand2_1 _07829_ (.A(_02943_),
    .B(_02735_),
    .Y(_02954_));
 sky130_fd_sc_hd__o22ai_4 _07830_ (.A1(net165),
    .A2(_01620_),
    .B1(_02746_),
    .B2(_02888_),
    .Y(_02965_));
 sky130_fd_sc_hd__o221a_1 _07831_ (.A1(net165),
    .A2(_01620_),
    .B1(_02188_),
    .B2(_02910_),
    .C1(_02932_),
    .X(_02976_));
 sky130_fd_sc_hd__o41ai_2 _07832_ (.A1(_01150_),
    .A2(_01161_),
    .A3(_01576_),
    .A4(_01598_),
    .B1(_02943_),
    .Y(_02987_));
 sky130_fd_sc_hd__o2111ai_4 _07833_ (.A1(_02188_),
    .A2(_02910_),
    .B1(_02932_),
    .C1(_01631_),
    .D1(_01194_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand3_4 _07834_ (.A(_02987_),
    .B(_02998_),
    .C(_02724_),
    .Y(_03009_));
 sky130_fd_sc_hd__o2bb2ai_2 _07835_ (.A1_N(_02735_),
    .A2_N(_02943_),
    .B1(_02702_),
    .B2(_02713_),
    .Y(_03020_));
 sky130_fd_sc_hd__o221ai_4 _07836_ (.A1(_02702_),
    .A2(_02713_),
    .B1(_02921_),
    .B2(_02965_),
    .C1(_02954_),
    .Y(_03030_));
 sky130_fd_sc_hd__o2bb2ai_2 _07837_ (.A1_N(_03009_),
    .A2_N(_03030_),
    .B1(_02188_),
    .B2(_02210_),
    .Y(_03041_));
 sky130_fd_sc_hd__o211ai_4 _07838_ (.A1(_02976_),
    .A2(_03020_),
    .B1(_03009_),
    .C1(_02221_),
    .Y(_03052_));
 sky130_fd_sc_hd__a21o_1 _07839_ (.A1(_03009_),
    .A2(_03030_),
    .B1(_02232_),
    .X(_03063_));
 sky130_fd_sc_hd__o211ai_1 _07840_ (.A1(_02188_),
    .A2(_02210_),
    .B1(_03009_),
    .C1(_03030_),
    .Y(_03074_));
 sky130_fd_sc_hd__a22oi_4 _07841_ (.A1(_02254_),
    .A2(_02669_),
    .B1(_03041_),
    .B2(_03052_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand3b_1 _07842_ (.A_N(_02691_),
    .B(_03063_),
    .C(_03074_),
    .Y(_03096_));
 sky130_fd_sc_hd__o211a_1 _07843_ (.A1(_02265_),
    .A2(_02680_),
    .B1(_03041_),
    .C1(_03052_),
    .X(_03107_));
 sky130_fd_sc_hd__a31oi_1 _07844_ (.A1(_03041_),
    .A2(_03052_),
    .A3(_02691_),
    .B1(_02658_),
    .Y(_03118_));
 sky130_fd_sc_hd__nor3_2 _07845_ (.A(_02658_),
    .B(_03085_),
    .C(_03107_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_1 _07846_ (.A(_03118_),
    .B(_03096_),
    .Y(_03140_));
 sky130_fd_sc_hd__o22a_1 _07847_ (.A1(_00310_),
    .A2(_02636_),
    .B1(_03085_),
    .B2(_03107_),
    .X(_03151_));
 sky130_fd_sc_hd__o22ai_2 _07848_ (.A1(_00310_),
    .A2(_02636_),
    .B1(_03085_),
    .B2(_03107_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand2_1 _07849_ (.A(_03162_),
    .B(_02571_),
    .Y(_03173_));
 sky130_fd_sc_hd__nand3_1 _07850_ (.A(_03162_),
    .B(_02571_),
    .C(_03140_),
    .Y(_03184_));
 sky130_fd_sc_hd__a2bb2oi_1 _07851_ (.A1_N(_02342_),
    .A2_N(_02560_),
    .B1(_03140_),
    .B2(_03162_),
    .Y(_03195_));
 sky130_fd_sc_hd__o22ai_2 _07852_ (.A1(_02342_),
    .A2(_02560_),
    .B1(_03129_),
    .B2(_03151_),
    .Y(_03206_));
 sky130_fd_sc_hd__o21ai_1 _07853_ (.A1(_03129_),
    .A2(_03173_),
    .B1(_03206_),
    .Y(_03217_));
 sky130_fd_sc_hd__a2bb2oi_2 _07854_ (.A1_N(_02462_),
    .A2_N(_02363_),
    .B1(_02451_),
    .B2(_02440_),
    .Y(_03228_));
 sky130_fd_sc_hd__xor2_2 _07855_ (.A(_03217_),
    .B(_03228_),
    .X(_03239_));
 sky130_fd_sc_hd__xnor2_1 _07856_ (.A(_02549_),
    .B(_03239_),
    .Y(net120));
 sky130_fd_sc_hd__o32a_1 _07857_ (.A1(_01860_),
    .A2(_02506_),
    .A3(_03239_),
    .B1(_00823_),
    .B2(_00812_),
    .X(_03259_));
 sky130_fd_sc_hd__o21ai_1 _07858_ (.A1(_02429_),
    .A2(_02484_),
    .B1(_03184_),
    .Y(_03270_));
 sky130_fd_sc_hd__o32a_1 _07859_ (.A1(_02429_),
    .A2(_02484_),
    .A3(_03195_),
    .B1(_03173_),
    .B2(_03129_),
    .X(_03281_));
 sky130_fd_sc_hd__a31o_2 _07860_ (.A1(_03096_),
    .A2(net33),
    .A3(_02647_),
    .B1(_03107_),
    .X(_03292_));
 sky130_fd_sc_hd__inv_2 _07861_ (.A(_03292_),
    .Y(_03303_));
 sky130_fd_sc_hd__a21oi_1 _07862_ (.A1(_02932_),
    .A2(_02965_),
    .B1(_02713_),
    .Y(_03314_));
 sky130_fd_sc_hd__a32o_1 _07863_ (.A1(_01303_),
    .A2(_01980_),
    .A3(_01969_),
    .B1(_02965_),
    .B2(_02932_),
    .X(_03325_));
 sky130_fd_sc_hd__and3_2 _07864_ (.A(_02713_),
    .B(_02932_),
    .C(_02965_),
    .X(_03336_));
 sky130_fd_sc_hd__nand3_1 _07865_ (.A(_02713_),
    .B(_02932_),
    .C(_02965_),
    .Y(_03347_));
 sky130_fd_sc_hd__nand2_1 _07866_ (.A(_03325_),
    .B(_03347_),
    .Y(_03358_));
 sky130_fd_sc_hd__o21ai_1 _07867_ (.A1(_01095_),
    .A2(_01117_),
    .B1(_02111_),
    .Y(_03369_));
 sky130_fd_sc_hd__o221a_2 _07868_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_02035_),
    .B2(_02057_),
    .C1(_01172_),
    .X(_03380_));
 sky130_fd_sc_hd__a22oi_4 _07869_ (.A1(_00932_),
    .A2(_00954_),
    .B1(_02779_),
    .B2(_00398_),
    .Y(_03391_));
 sky130_fd_sc_hd__o211ai_2 _07870_ (.A1(_00921_),
    .A2(_00943_),
    .B1(_02822_),
    .C1(_02844_),
    .Y(_03402_));
 sky130_fd_sc_hd__nand4_4 _07871_ (.A(_01216_),
    .B(_02002_),
    .C(_00376_),
    .D(_00398_),
    .Y(_03413_));
 sky130_fd_sc_hd__a41o_1 _07872_ (.A1(_01216_),
    .A2(_02002_),
    .A3(_00376_),
    .A4(_00398_),
    .B1(_00299_),
    .X(_03424_));
 sky130_fd_sc_hd__o311a_4 _07873_ (.A1(net59),
    .A2(net60),
    .A3(_02024_),
    .B1(_00419_),
    .C1(net173),
    .X(_03435_));
 sky130_fd_sc_hd__a311o_2 _07874_ (.A1(_02013_),
    .A2(_00398_),
    .A3(_00376_),
    .B1(_00299_),
    .C1(net61),
    .X(_03446_));
 sky130_fd_sc_hd__a21oi_4 _07875_ (.A1(_03413_),
    .A2(net173),
    .B1(_00419_),
    .Y(_03457_));
 sky130_fd_sc_hd__a21o_1 _07876_ (.A1(_03413_),
    .A2(net173),
    .B1(_00419_),
    .X(_03468_));
 sky130_fd_sc_hd__a21oi_4 _07877_ (.A1(_03413_),
    .A2(net173),
    .B1(net61),
    .Y(_03479_));
 sky130_fd_sc_hd__a21o_4 _07878_ (.A1(_03413_),
    .A2(net173),
    .B1(net61),
    .X(_03490_));
 sky130_fd_sc_hd__a41oi_4 _07879_ (.A1(_01216_),
    .A2(_02002_),
    .A3(_00376_),
    .A4(_00398_),
    .B1(_00419_),
    .Y(_03501_));
 sky130_fd_sc_hd__nand2_8 _07880_ (.A(_03413_),
    .B(net61),
    .Y(_03511_));
 sky130_fd_sc_hd__o311a_4 _07881_ (.A1(net59),
    .A2(net60),
    .A3(_02024_),
    .B1(net61),
    .C1(net173),
    .X(_03522_));
 sky130_fd_sc_hd__o211ai_4 _07882_ (.A1(net60),
    .A2(_02757_),
    .B1(net61),
    .C1(net173),
    .Y(_03533_));
 sky130_fd_sc_hd__o21ai_4 _07883_ (.A1(_00299_),
    .A2(_03511_),
    .B1(_03490_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21oi_4 _07884_ (.A1(net173),
    .A2(_03501_),
    .B1(_03479_),
    .Y(_03555_));
 sky130_fd_sc_hd__nand3_2 _07885_ (.A(_03490_),
    .B(_03533_),
    .C(net1),
    .Y(_03566_));
 sky130_fd_sc_hd__nand4_4 _07886_ (.A(_03391_),
    .B(_03490_),
    .C(_03533_),
    .D(_02822_),
    .Y(_03577_));
 sky130_fd_sc_hd__nor2_2 _07887_ (.A(_03402_),
    .B(_03566_),
    .Y(_03588_));
 sky130_fd_sc_hd__o2111ai_4 _07888_ (.A1(_00398_),
    .A2(_02779_),
    .B1(_03391_),
    .C1(net1),
    .D1(net157),
    .Y(_03599_));
 sky130_fd_sc_hd__a32oi_4 _07889_ (.A1(_03490_),
    .A2(_03533_),
    .A3(net1),
    .B1(_03391_),
    .B2(_02822_),
    .Y(_03610_));
 sky130_fd_sc_hd__o31ai_4 _07890_ (.A1(_00987_),
    .A2(net167),
    .A3(_02833_),
    .B1(_03566_),
    .Y(_03621_));
 sky130_fd_sc_hd__a22oi_4 _07891_ (.A1(_01194_),
    .A2(_02133_),
    .B1(_03599_),
    .B2(_03621_),
    .Y(_03632_));
 sky130_fd_sc_hd__o22ai_4 _07892_ (.A1(_03369_),
    .A2(_02079_),
    .B1(_03610_),
    .B2(_03588_),
    .Y(_03643_));
 sky130_fd_sc_hd__o21a_1 _07893_ (.A1(_03402_),
    .A2(_03566_),
    .B1(_03380_),
    .X(_03654_));
 sky130_fd_sc_hd__o211a_1 _07894_ (.A1(_00288_),
    .A2(_03577_),
    .B1(_03380_),
    .C1(_03621_),
    .X(_03665_));
 sky130_fd_sc_hd__o211ai_2 _07895_ (.A1(_00288_),
    .A2(_03577_),
    .B1(_03380_),
    .C1(_03621_),
    .Y(_03676_));
 sky130_fd_sc_hd__a22o_1 _07896_ (.A1(_01434_),
    .A2(_01455_),
    .B1(_01543_),
    .B2(_01565_),
    .X(_03687_));
 sky130_fd_sc_hd__a22oi_2 _07897_ (.A1(_01499_),
    .A2(_01631_),
    .B1(_03643_),
    .B2(_03676_),
    .Y(_03698_));
 sky130_fd_sc_hd__o22ai_2 _07898_ (.A1(_01488_),
    .A2(_01620_),
    .B1(_03632_),
    .B2(_03665_),
    .Y(_03709_));
 sky130_fd_sc_hd__a211oi_2 _07899_ (.A1(_03654_),
    .A2(_03621_),
    .B1(_03687_),
    .C1(_03632_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand3b_1 _07900_ (.A_N(_03687_),
    .B(_03676_),
    .C(_03643_),
    .Y(_03731_));
 sky130_fd_sc_hd__o22ai_2 _07901_ (.A1(_03314_),
    .A2(_03336_),
    .B1(_03698_),
    .B2(_03720_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand4_2 _07902_ (.A(_03325_),
    .B(_03347_),
    .C(_03709_),
    .D(_03731_),
    .Y(_03753_));
 sky130_fd_sc_hd__o21bai_1 _07903_ (.A1(_03698_),
    .A2(_03720_),
    .B1_N(_03358_),
    .Y(_03763_));
 sky130_fd_sc_hd__o211ai_1 _07904_ (.A1(_03314_),
    .A2(_03336_),
    .B1(_03709_),
    .C1(_03731_),
    .Y(_03774_));
 sky130_fd_sc_hd__a2bb2oi_1 _07905_ (.A1_N(_02976_),
    .A2_N(_03020_),
    .B1(_03009_),
    .B2(_02232_),
    .Y(_03785_));
 sky130_fd_sc_hd__a2bb2o_1 _07906_ (.A1_N(_02976_),
    .A2_N(_03020_),
    .B1(_03009_),
    .B2(_02232_),
    .X(_03796_));
 sky130_fd_sc_hd__nand3_4 _07907_ (.A(_03742_),
    .B(_03753_),
    .C(_03785_),
    .Y(_03807_));
 sky130_fd_sc_hd__and3_2 _07908_ (.A(_03763_),
    .B(_03774_),
    .C(_03796_),
    .X(_03818_));
 sky130_fd_sc_hd__nand3_2 _07909_ (.A(_03763_),
    .B(_03774_),
    .C(_03796_),
    .Y(_03829_));
 sky130_fd_sc_hd__nor2_4 _07910_ (.A(net27),
    .B(net28),
    .Y(_03840_));
 sky130_fd_sc_hd__nand4_2 _07911_ (.A(_01074_),
    .B(_03840_),
    .C(_00343_),
    .D(_00365_),
    .Y(_03851_));
 sky130_fd_sc_hd__a311o_4 _07912_ (.A1(_01412_),
    .A2(_03840_),
    .A3(_00365_),
    .B1(net29),
    .C1(_00321_),
    .X(_03862_));
 sky130_fd_sc_hd__a21o_2 _07913_ (.A1(_03851_),
    .A2(net174),
    .B1(_00430_),
    .X(_03873_));
 sky130_fd_sc_hd__a21o_1 _07914_ (.A1(_03851_),
    .A2(net174),
    .B1(net29),
    .X(_03884_));
 sky130_fd_sc_hd__a311o_2 _07915_ (.A1(_01412_),
    .A2(_03840_),
    .A3(_00365_),
    .B1(_00430_),
    .C1(_00321_),
    .X(_03895_));
 sky130_fd_sc_hd__nand2_8 _07916_ (.A(_03884_),
    .B(_03895_),
    .Y(_03906_));
 sky130_fd_sc_hd__nand2_8 _07917_ (.A(_03862_),
    .B(_03873_),
    .Y(_03917_));
 sky130_fd_sc_hd__a21o_1 _07918_ (.A1(_03862_),
    .A2(_03873_),
    .B1(_00310_),
    .X(_03928_));
 sky130_fd_sc_hd__o22a_1 _07919_ (.A1(_01292_),
    .A2(_01958_),
    .B1(_02636_),
    .B2(_00900_),
    .X(_03939_));
 sky130_fd_sc_hd__a32o_1 _07920_ (.A1(_00911_),
    .A2(_02614_),
    .A3(_02625_),
    .B1(_01303_),
    .B2(_01969_),
    .X(_03950_));
 sky130_fd_sc_hd__nand4_2 _07921_ (.A(_00911_),
    .B(_01303_),
    .C(_01969_),
    .D(_02647_),
    .Y(_03961_));
 sky130_fd_sc_hd__o2bb2a_1 _07922_ (.A1_N(_03950_),
    .A2_N(_03961_),
    .B1(_00310_),
    .B2(_03906_),
    .X(_03972_));
 sky130_fd_sc_hd__and4_1 _07923_ (.A(_03950_),
    .B(net33),
    .C(_03917_),
    .D(_03961_),
    .X(_03983_));
 sky130_fd_sc_hd__a21oi_1 _07924_ (.A1(_03950_),
    .A2(_03961_),
    .B1(_03928_),
    .Y(_03993_));
 sky130_fd_sc_hd__and3_1 _07925_ (.A(_03928_),
    .B(_03950_),
    .C(_03961_),
    .X(_04004_));
 sky130_fd_sc_hd__nor2_1 _07926_ (.A(_03993_),
    .B(_04004_),
    .Y(_04015_));
 sky130_fd_sc_hd__o211ai_1 _07927_ (.A1(_03972_),
    .A2(_03983_),
    .B1(_03807_),
    .C1(_03829_),
    .Y(_04026_));
 sky130_fd_sc_hd__o2bb2ai_1 _07928_ (.A1_N(_03807_),
    .A2_N(_03829_),
    .B1(_03993_),
    .B2(_04004_),
    .Y(_04037_));
 sky130_fd_sc_hd__o211ai_2 _07929_ (.A1(_03993_),
    .A2(_04004_),
    .B1(_03807_),
    .C1(_03829_),
    .Y(_04048_));
 sky130_fd_sc_hd__a21bo_1 _07930_ (.A1(_03807_),
    .A2(_03829_),
    .B1_N(_04015_),
    .X(_04059_));
 sky130_fd_sc_hd__nand2_1 _07931_ (.A(_04048_),
    .B(_04059_),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_2 _07932_ (.A(_04026_),
    .B(_04037_),
    .Y(_04081_));
 sky130_fd_sc_hd__a311o_1 _07933_ (.A1(net33),
    .A2(_02647_),
    .A3(_03096_),
    .B1(_03107_),
    .C1(_04081_),
    .X(_04092_));
 sky130_fd_sc_hd__nand3_2 _07934_ (.A(_04059_),
    .B(_03292_),
    .C(_04048_),
    .Y(_04103_));
 sky130_fd_sc_hd__a21oi_1 _07935_ (.A1(_04092_),
    .A2(_04103_),
    .B1(_03281_),
    .Y(_04114_));
 sky130_fd_sc_hd__o2111ai_1 _07936_ (.A1(_03228_),
    .A2(_03195_),
    .B1(_03184_),
    .C1(_04103_),
    .D1(_04092_),
    .Y(_04125_));
 sky130_fd_sc_hd__and2b_1 _07937_ (.A_N(_04114_),
    .B(_04125_),
    .X(_04136_));
 sky130_fd_sc_hd__xnor2_1 _07938_ (.A(_03259_),
    .B(_04136_),
    .Y(net125));
 sky130_fd_sc_hd__nor4b_2 _07939_ (.A(_01860_),
    .B(_02506_),
    .C(_03239_),
    .D_N(_04136_),
    .Y(_04157_));
 sky130_fd_sc_hd__o21a_1 _07940_ (.A1(_03972_),
    .A2(_03983_),
    .B1(_03807_),
    .X(_04168_));
 sky130_fd_sc_hd__o21ai_4 _07941_ (.A1(_04015_),
    .A2(_03818_),
    .B1(_03807_),
    .Y(_04179_));
 sky130_fd_sc_hd__nand4_4 _07942_ (.A(_01412_),
    .B(_03840_),
    .C(_00365_),
    .D(_00430_),
    .Y(_04190_));
 sky130_fd_sc_hd__a311o_4 _07943_ (.A1(net171),
    .A2(_03840_),
    .A3(_00430_),
    .B1(net30),
    .C1(_00321_),
    .X(_04201_));
 sky130_fd_sc_hd__a21o_4 _07944_ (.A1(_04190_),
    .A2(net174),
    .B1(_00452_),
    .X(_04212_));
 sky130_fd_sc_hd__a311o_4 _07945_ (.A1(net171),
    .A2(_03840_),
    .A3(_00430_),
    .B1(_00452_),
    .C1(_00321_),
    .X(_04222_));
 sky130_fd_sc_hd__a21o_4 _07946_ (.A1(_04190_),
    .A2(net174),
    .B1(net30),
    .X(_04233_));
 sky130_fd_sc_hd__nand2_8 _07947_ (.A(_04222_),
    .B(_04233_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_8 _07948_ (.A(_04201_),
    .B(_04212_),
    .Y(_04255_));
 sky130_fd_sc_hd__and4_2 _07949_ (.A(_00911_),
    .B(_01303_),
    .C(_02647_),
    .D(_03917_),
    .X(_04266_));
 sky130_fd_sc_hd__o22a_1 _07950_ (.A1(_01292_),
    .A2(_02636_),
    .B1(_03906_),
    .B2(_00900_),
    .X(_04277_));
 sky130_fd_sc_hd__a32o_1 _07951_ (.A1(_01303_),
    .A2(_02614_),
    .A3(_02625_),
    .B1(_03917_),
    .B2(_00911_),
    .X(_04288_));
 sky130_fd_sc_hd__o22a_2 _07952_ (.A1(_04244_),
    .A2(_00310_),
    .B1(_04277_),
    .B2(_04266_),
    .X(_04299_));
 sky130_fd_sc_hd__and4b_2 _07953_ (.A_N(_04266_),
    .B(net33),
    .C(_04255_),
    .D(_04288_),
    .X(_04310_));
 sky130_fd_sc_hd__o211a_1 _07954_ (.A1(_04266_),
    .A2(_04277_),
    .B1(net33),
    .C1(_04255_),
    .X(_04321_));
 sky130_fd_sc_hd__a311oi_4 _07955_ (.A1(net33),
    .A2(_04222_),
    .A3(_04233_),
    .B1(_04266_),
    .C1(_04277_),
    .Y(_04332_));
 sky130_fd_sc_hd__and3_2 _07956_ (.A(_03325_),
    .B(_03709_),
    .C(_03731_),
    .X(_04343_));
 sky130_fd_sc_hd__o31a_1 _07957_ (.A1(_03314_),
    .A2(_03698_),
    .A3(_03720_),
    .B1(_03347_),
    .X(_04354_));
 sky130_fd_sc_hd__o21ai_1 _07958_ (.A1(_00310_),
    .A2(_03906_),
    .B1(_03961_),
    .Y(_04365_));
 sky130_fd_sc_hd__a21oi_1 _07959_ (.A1(_03928_),
    .A2(_03961_),
    .B1(_03939_),
    .Y(_04376_));
 sky130_fd_sc_hd__o21ai_1 _07960_ (.A1(_01488_),
    .A2(_01620_),
    .B1(_03676_),
    .Y(_04387_));
 sky130_fd_sc_hd__nand3_2 _07961_ (.A(_03643_),
    .B(_04376_),
    .C(_04387_),
    .Y(_04398_));
 sky130_fd_sc_hd__inv_2 _07962_ (.A(_04398_),
    .Y(_04409_));
 sky130_fd_sc_hd__o2bb2ai_2 _07963_ (.A1_N(_03950_),
    .A2_N(_04365_),
    .B1(_03687_),
    .B2(_03632_),
    .Y(_04420_));
 sky130_fd_sc_hd__a31o_1 _07964_ (.A1(_03380_),
    .A2(_03599_),
    .A3(_03621_),
    .B1(_04420_),
    .X(_04430_));
 sky130_fd_sc_hd__o21a_1 _07965_ (.A1(_03665_),
    .A2(_04420_),
    .B1(_04398_),
    .X(_04441_));
 sky130_fd_sc_hd__o21ai_2 _07966_ (.A1(_03665_),
    .A2(_04420_),
    .B1(_04398_),
    .Y(_04452_));
 sky130_fd_sc_hd__and3_1 _07967_ (.A(_01631_),
    .B(_01936_),
    .C(_01947_),
    .X(_04463_));
 sky130_fd_sc_hd__nand4_4 _07968_ (.A(_01587_),
    .B(_01609_),
    .C(_01936_),
    .D(_01947_),
    .Y(_04474_));
 sky130_fd_sc_hd__o32a_1 _07969_ (.A1(_01488_),
    .A2(_02079_),
    .A3(_02100_),
    .B1(_01620_),
    .B2(_01958_),
    .X(_04485_));
 sky130_fd_sc_hd__o21ai_1 _07970_ (.A1(_01488_),
    .A2(_02122_),
    .B1(_04474_),
    .Y(_04496_));
 sky130_fd_sc_hd__and4_1 _07971_ (.A(_01499_),
    .B(_01631_),
    .C(_01969_),
    .D(_02133_),
    .X(_04507_));
 sky130_fd_sc_hd__nand4_2 _07972_ (.A(_01499_),
    .B(_01631_),
    .C(_01969_),
    .D(_02133_),
    .Y(_04518_));
 sky130_fd_sc_hd__o31a_1 _07973_ (.A1(_01958_),
    .A2(_02122_),
    .A3(_03687_),
    .B1(_04496_),
    .X(_04529_));
 sky130_fd_sc_hd__nand2_2 _07974_ (.A(_04496_),
    .B(_04518_),
    .Y(_04540_));
 sky130_fd_sc_hd__o221a_1 _07975_ (.A1(_00321_),
    .A2(_01139_),
    .B1(net169),
    .B2(_02800_),
    .C1(_01172_),
    .X(_04551_));
 sky130_fd_sc_hd__or4_1 _07976_ (.A(_01150_),
    .B(_01161_),
    .C(net167),
    .D(_02833_),
    .X(_04562_));
 sky130_fd_sc_hd__a22oi_4 _07977_ (.A1(_00932_),
    .A2(_00954_),
    .B1(_03424_),
    .B2(_00419_),
    .Y(_04573_));
 sky130_fd_sc_hd__o221ai_4 _07978_ (.A1(_00299_),
    .A2(_03511_),
    .B1(_00943_),
    .B2(_00921_),
    .C1(_03490_),
    .Y(_04584_));
 sky130_fd_sc_hd__nor2_2 _07979_ (.A(net60),
    .B(net61),
    .Y(_04595_));
 sky130_fd_sc_hd__and4_4 _07980_ (.A(_01216_),
    .B(_02002_),
    .C(_04595_),
    .D(_00376_),
    .X(_04606_));
 sky130_fd_sc_hd__nand4_4 _07981_ (.A(_01216_),
    .B(_02002_),
    .C(_04595_),
    .D(_00376_),
    .Y(_04616_));
 sky130_fd_sc_hd__a41oi_1 _07982_ (.A1(_01216_),
    .A2(_02002_),
    .A3(_04595_),
    .A4(_00376_),
    .B1(_00299_),
    .Y(_04627_));
 sky130_fd_sc_hd__o311a_4 _07983_ (.A1(net60),
    .A2(net61),
    .A3(_02757_),
    .B1(_00441_),
    .C1(net173),
    .X(_04638_));
 sky130_fd_sc_hd__a21oi_4 _07984_ (.A1(_04616_),
    .A2(net173),
    .B1(_00441_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_8 _07985_ (.A(net173),
    .B(net62),
    .Y(_04660_));
 sky130_fd_sc_hd__a31oi_4 _07986_ (.A1(_02013_),
    .A2(_04595_),
    .A3(_00376_),
    .B1(_04660_),
    .Y(_04671_));
 sky130_fd_sc_hd__a31o_4 _07987_ (.A1(_02013_),
    .A2(_04595_),
    .A3(_00376_),
    .B1(_04660_),
    .X(_04682_));
 sky130_fd_sc_hd__a21oi_4 _07988_ (.A1(_04616_),
    .A2(net173),
    .B1(net62),
    .Y(_04693_));
 sky130_fd_sc_hd__a21o_4 _07989_ (.A1(_04616_),
    .A2(net173),
    .B1(net62),
    .X(_04704_));
 sky130_fd_sc_hd__o21ai_4 _07990_ (.A1(_04606_),
    .A2(_04660_),
    .B1(_04704_),
    .Y(_04715_));
 sky130_fd_sc_hd__nor2_8 _07991_ (.A(_04671_),
    .B(_04693_),
    .Y(_04726_));
 sky130_fd_sc_hd__o21a_1 _07992_ (.A1(net62),
    .A2(_04627_),
    .B1(net1),
    .X(_04737_));
 sky130_fd_sc_hd__o211ai_2 _07993_ (.A1(_04606_),
    .A2(_04660_),
    .B1(net1),
    .C1(_04704_),
    .Y(_04748_));
 sky130_fd_sc_hd__a32oi_4 _07994_ (.A1(_04704_),
    .A2(net1),
    .A3(_04682_),
    .B1(_04573_),
    .B2(_03533_),
    .Y(_04759_));
 sky130_fd_sc_hd__o31ai_4 _07995_ (.A1(_00288_),
    .A2(_04671_),
    .A3(_04693_),
    .B1(_04584_),
    .Y(_04770_));
 sky130_fd_sc_hd__nor2_2 _07996_ (.A(_04584_),
    .B(_04748_),
    .Y(_04781_));
 sky130_fd_sc_hd__nand4_4 _07997_ (.A(net157),
    .B(_04737_),
    .C(_04682_),
    .D(_00998_),
    .Y(_04792_));
 sky130_fd_sc_hd__o21a_1 _07998_ (.A1(_04584_),
    .A2(_04748_),
    .B1(_04551_),
    .X(_04802_));
 sky130_fd_sc_hd__o2111ai_4 _07999_ (.A1(_01095_),
    .A2(_01117_),
    .B1(_02866_),
    .C1(_04770_),
    .D1(_04792_),
    .Y(_04813_));
 sky130_fd_sc_hd__a2bb2oi_1 _08000_ (.A1_N(net165),
    .A2_N(_02855_),
    .B1(_04770_),
    .B2(_04792_),
    .Y(_04824_));
 sky130_fd_sc_hd__o22ai_4 _08001_ (.A1(net165),
    .A2(_02855_),
    .B1(_04759_),
    .B2(_04781_),
    .Y(_04835_));
 sky130_fd_sc_hd__o21ai_1 _08002_ (.A1(_04759_),
    .A2(_04781_),
    .B1(_04551_),
    .Y(_04846_));
 sky130_fd_sc_hd__o211ai_2 _08003_ (.A1(net165),
    .A2(_02855_),
    .B1(_04770_),
    .C1(_04792_),
    .Y(_04857_));
 sky130_fd_sc_hd__a211oi_4 _08004_ (.A1(_04802_),
    .A2(_04770_),
    .B1(_04540_),
    .C1(_04824_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand3_2 _08005_ (.A(_04835_),
    .B(_04529_),
    .C(_04813_),
    .Y(_04879_));
 sky130_fd_sc_hd__a2bb2oi_2 _08006_ (.A1_N(_04485_),
    .A2_N(_04507_),
    .B1(_04813_),
    .B2(_04835_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand3_4 _08007_ (.A(_04540_),
    .B(_04846_),
    .C(_04857_),
    .Y(_04901_));
 sky130_fd_sc_hd__o2bb2ai_2 _08008_ (.A1_N(_04879_),
    .A2_N(_04901_),
    .B1(_00288_),
    .B2(_03577_),
    .Y(_04912_));
 sky130_fd_sc_hd__nand3_2 _08009_ (.A(_04901_),
    .B(_03588_),
    .C(_04879_),
    .Y(_04923_));
 sky130_fd_sc_hd__o21ai_1 _08010_ (.A1(_00288_),
    .A2(_03577_),
    .B1(_04901_),
    .Y(_04934_));
 sky130_fd_sc_hd__o211ai_1 _08011_ (.A1(_00288_),
    .A2(_03577_),
    .B1(_04879_),
    .C1(_04901_),
    .Y(_04945_));
 sky130_fd_sc_hd__o21ai_2 _08012_ (.A1(_04868_),
    .A2(_04890_),
    .B1(_03588_),
    .Y(_04956_));
 sky130_fd_sc_hd__nand3_2 _08013_ (.A(_04452_),
    .B(_04912_),
    .C(_04923_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand3_2 _08014_ (.A(_04956_),
    .B(_04441_),
    .C(_04945_),
    .Y(_04978_));
 sky130_fd_sc_hd__o211ai_4 _08015_ (.A1(_04934_),
    .A2(_04868_),
    .B1(_04452_),
    .C1(_04956_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand3_2 _08016_ (.A(_04441_),
    .B(_04912_),
    .C(_04923_),
    .Y(_04999_));
 sky130_fd_sc_hd__a2bb2oi_4 _08017_ (.A1_N(_03336_),
    .A2_N(_04343_),
    .B1(_04967_),
    .B2(_04978_),
    .Y(_05010_));
 sky130_fd_sc_hd__o211ai_4 _08018_ (.A1(_03336_),
    .A2(_04343_),
    .B1(_04988_),
    .C1(_04999_),
    .Y(_05021_));
 sky130_fd_sc_hd__a21boi_2 _08019_ (.A1(_04988_),
    .A2(_04999_),
    .B1_N(_04354_),
    .Y(_05032_));
 sky130_fd_sc_hd__nand3_2 _08020_ (.A(_04354_),
    .B(_04967_),
    .C(_04978_),
    .Y(_05043_));
 sky130_fd_sc_hd__o21a_1 _08021_ (.A1(_04321_),
    .A2(_04332_),
    .B1(_05043_),
    .X(_05054_));
 sky130_fd_sc_hd__o211a_1 _08022_ (.A1(_04321_),
    .A2(_04332_),
    .B1(_05021_),
    .C1(_05043_),
    .X(_05065_));
 sky130_fd_sc_hd__o211ai_1 _08023_ (.A1(_04321_),
    .A2(_04332_),
    .B1(_05021_),
    .C1(_05043_),
    .Y(_05076_));
 sky130_fd_sc_hd__o22ai_2 _08024_ (.A1(_04299_),
    .A2(_04310_),
    .B1(_05010_),
    .B2(_05032_),
    .Y(_05087_));
 sky130_fd_sc_hd__o211ai_4 _08025_ (.A1(_04299_),
    .A2(_04310_),
    .B1(_05021_),
    .C1(_05043_),
    .Y(_05098_));
 sky130_fd_sc_hd__o22ai_4 _08026_ (.A1(_04321_),
    .A2(_04332_),
    .B1(_05010_),
    .B2(_05032_),
    .Y(_05109_));
 sky130_fd_sc_hd__nand2_2 _08027_ (.A(_05098_),
    .B(_05109_),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(_05087_),
    .B(_04179_),
    .Y(_05131_));
 sky130_fd_sc_hd__nand3_2 _08029_ (.A(_05087_),
    .B(_04179_),
    .C(_05076_),
    .Y(_05142_));
 sky130_fd_sc_hd__o211ai_4 _08030_ (.A1(_03818_),
    .A2(_04168_),
    .B1(_05098_),
    .C1(_05109_),
    .Y(_05153_));
 sky130_fd_sc_hd__o211ai_4 _08031_ (.A1(_03292_),
    .A2(_04081_),
    .B1(_03206_),
    .C1(_03270_),
    .Y(_05164_));
 sky130_fd_sc_hd__o221ai_2 _08032_ (.A1(_03129_),
    .A2(_03173_),
    .B1(_03228_),
    .B2(_03195_),
    .C1(_04103_),
    .Y(_05174_));
 sky130_fd_sc_hd__a22oi_1 _08033_ (.A1(_05142_),
    .A2(_05153_),
    .B1(_05164_),
    .B2(_04103_),
    .Y(_05185_));
 sky130_fd_sc_hd__and4_1 _08034_ (.A(_04103_),
    .B(_05142_),
    .C(_05153_),
    .D(_05164_),
    .X(_05196_));
 sky130_fd_sc_hd__nor2_1 _08035_ (.A(_05185_),
    .B(_05196_),
    .Y(_05207_));
 sky130_fd_sc_hd__or3_1 _08036_ (.A(_00834_),
    .B(_04157_),
    .C(_05207_),
    .X(_05218_));
 sky130_fd_sc_hd__o21ai_1 _08037_ (.A1(_00834_),
    .A2(_04157_),
    .B1(_05207_),
    .Y(_05229_));
 sky130_fd_sc_hd__and2_1 _08038_ (.A(_05218_),
    .B(_05229_),
    .X(net126));
 sky130_fd_sc_hd__o2bb2a_1 _08039_ (.A1_N(_04157_),
    .A2_N(_05207_),
    .B1(_00812_),
    .B2(_00823_),
    .X(_05250_));
 sky130_fd_sc_hd__nand4_4 _08040_ (.A(net171),
    .B(_03840_),
    .C(_00430_),
    .D(_00452_),
    .Y(_05261_));
 sky130_fd_sc_hd__o211ai_4 _08041_ (.A1(net30),
    .A2(_04190_),
    .B1(net31),
    .C1(net174),
    .Y(_05272_));
 sky130_fd_sc_hd__a21o_4 _08042_ (.A1(_05261_),
    .A2(net174),
    .B1(net31),
    .X(_05283_));
 sky130_fd_sc_hd__a21bo_2 _08043_ (.A1(_05261_),
    .A2(net174),
    .B1_N(net31),
    .X(_05294_));
 sky130_fd_sc_hd__nand3b_4 _08044_ (.A_N(net31),
    .B(_05261_),
    .C(net174),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_8 _08045_ (.A(_05294_),
    .B(_05305_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_8 _08046_ (.A(_05272_),
    .B(_05283_),
    .Y(_05327_));
 sky130_fd_sc_hd__a21o_1 _08047_ (.A1(_05294_),
    .A2(_05305_),
    .B1(_00310_),
    .X(_05337_));
 sky130_fd_sc_hd__nor2_4 _08048_ (.A(net62),
    .B(_04616_),
    .Y(_05348_));
 sky130_fd_sc_hd__o311a_4 _08049_ (.A1(net61),
    .A2(net62),
    .A3(_03413_),
    .B1(_00463_),
    .C1(net173),
    .X(_05359_));
 sky130_fd_sc_hd__o21a_4 _08050_ (.A1(_00299_),
    .A2(_05348_),
    .B1(net63),
    .X(_05370_));
 sky130_fd_sc_hd__o311a_4 _08051_ (.A1(net61),
    .A2(net62),
    .A3(_03413_),
    .B1(net63),
    .C1(net173),
    .X(_05381_));
 sky130_fd_sc_hd__or3_4 _08052_ (.A(_00299_),
    .B(_00463_),
    .C(_05348_),
    .X(_05392_));
 sky130_fd_sc_hd__o21a_4 _08053_ (.A1(_00299_),
    .A2(_05348_),
    .B1(_00463_),
    .X(_05403_));
 sky130_fd_sc_hd__o21ai_4 _08054_ (.A1(_00299_),
    .A2(_05348_),
    .B1(_00463_),
    .Y(_05414_));
 sky130_fd_sc_hd__nor2_8 _08055_ (.A(_05359_),
    .B(_05370_),
    .Y(_05425_));
 sky130_fd_sc_hd__nor2_8 _08056_ (.A(_05381_),
    .B(_05403_),
    .Y(_05436_));
 sky130_fd_sc_hd__a22o_1 _08057_ (.A1(_02046_),
    .A2(_02068_),
    .B1(_02592_),
    .B2(_02603_),
    .X(_05447_));
 sky130_fd_sc_hd__nor3_2 _08058_ (.A(_02122_),
    .B(_04474_),
    .C(_02636_),
    .Y(_05458_));
 sky130_fd_sc_hd__or4_1 _08059_ (.A(_01620_),
    .B(_01958_),
    .C(_02122_),
    .D(_02636_),
    .X(_05469_));
 sky130_fd_sc_hd__a22oi_4 _08060_ (.A1(_01969_),
    .A2(_02133_),
    .B1(_02647_),
    .B2(_01631_),
    .Y(_05480_));
 sky130_fd_sc_hd__a31oi_2 _08061_ (.A1(_02133_),
    .A2(_02647_),
    .A3(_04463_),
    .B1(_05480_),
    .Y(_05491_));
 sky130_fd_sc_hd__o221ai_4 _08062_ (.A1(_00921_),
    .A2(_00943_),
    .B1(_04606_),
    .B2(_04660_),
    .C1(_04704_),
    .Y(_05501_));
 sky130_fd_sc_hd__and3_1 _08063_ (.A(_01194_),
    .B(_03490_),
    .C(_03533_),
    .X(_05512_));
 sky130_fd_sc_hd__o211ai_4 _08064_ (.A1(_00299_),
    .A2(_03511_),
    .B1(_03490_),
    .C1(_01194_),
    .Y(_05523_));
 sky130_fd_sc_hd__nand2_2 _08065_ (.A(_05501_),
    .B(_05523_),
    .Y(_05534_));
 sky130_fd_sc_hd__o211ai_4 _08066_ (.A1(_04660_),
    .A2(_04606_),
    .B1(_01194_),
    .C1(_04704_),
    .Y(_05545_));
 sky130_fd_sc_hd__nand4_2 _08067_ (.A(_04573_),
    .B(_04726_),
    .C(_01194_),
    .D(_03533_),
    .Y(_05556_));
 sky130_fd_sc_hd__o2bb2ai_1 _08068_ (.A1_N(_05501_),
    .A2_N(_05523_),
    .B1(_05545_),
    .B2(_04584_),
    .Y(_05567_));
 sky130_fd_sc_hd__and3_1 _08069_ (.A(_01499_),
    .B(_02822_),
    .C(_02844_),
    .X(_05578_));
 sky130_fd_sc_hd__a211o_1 _08070_ (.A1(_01434_),
    .A2(_01455_),
    .B1(net167),
    .C1(_02833_),
    .X(_05589_));
 sky130_fd_sc_hd__o21ai_1 _08071_ (.A1(_01488_),
    .A2(_02855_),
    .B1(_05567_),
    .Y(_05600_));
 sky130_fd_sc_hd__o2111ai_4 _08072_ (.A1(_04584_),
    .A2(_05545_),
    .B1(_05534_),
    .C1(_01499_),
    .D1(_02866_),
    .Y(_05611_));
 sky130_fd_sc_hd__o221ai_4 _08073_ (.A1(_01488_),
    .A2(_02855_),
    .B1(_04584_),
    .B2(_05545_),
    .C1(_05534_),
    .Y(_05622_));
 sky130_fd_sc_hd__nand2_1 _08074_ (.A(_05567_),
    .B(_05578_),
    .Y(_05633_));
 sky130_fd_sc_hd__o211ai_4 _08075_ (.A1(_05458_),
    .A2(_05480_),
    .B1(_05622_),
    .C1(_05633_),
    .Y(_05644_));
 sky130_fd_sc_hd__nand3_4 _08076_ (.A(_05491_),
    .B(_05600_),
    .C(_05611_),
    .Y(_05654_));
 sky130_fd_sc_hd__and3_1 _08077_ (.A(_01194_),
    .B(_02866_),
    .C(_04770_),
    .X(_05665_));
 sky130_fd_sc_hd__o31a_1 _08078_ (.A1(net165),
    .A2(_02855_),
    .A3(_04759_),
    .B1(_04792_),
    .X(_05676_));
 sky130_fd_sc_hd__o2111ai_4 _08079_ (.A1(_04562_),
    .A2(_04759_),
    .B1(_04792_),
    .C1(_05644_),
    .D1(_05654_),
    .Y(_05687_));
 sky130_fd_sc_hd__o2bb2ai_2 _08080_ (.A1_N(_05644_),
    .A2_N(_05654_),
    .B1(_05665_),
    .B2(_04781_),
    .Y(_05698_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_05687_),
    .B(_05698_),
    .Y(_05709_));
 sky130_fd_sc_hd__a31oi_2 _08082_ (.A1(_04288_),
    .A2(net33),
    .A3(_04255_),
    .B1(_04266_),
    .Y(_05720_));
 sky130_fd_sc_hd__a31o_1 _08083_ (.A1(_04288_),
    .A2(net33),
    .A3(_04255_),
    .B1(_04266_),
    .X(_05731_));
 sky130_fd_sc_hd__a31oi_1 _08084_ (.A1(_04835_),
    .A2(_04529_),
    .A3(_04813_),
    .B1(_03588_),
    .Y(_05742_));
 sky130_fd_sc_hd__a31o_1 _08085_ (.A1(_04835_),
    .A2(_04529_),
    .A3(_04813_),
    .B1(_03588_),
    .X(_05753_));
 sky130_fd_sc_hd__nor3_2 _08086_ (.A(_04890_),
    .B(_05720_),
    .C(_05742_),
    .Y(_05764_));
 sky130_fd_sc_hd__nand3_4 _08087_ (.A(_04901_),
    .B(_05731_),
    .C(_05753_),
    .Y(_05775_));
 sky130_fd_sc_hd__o211a_1 _08088_ (.A1(_03599_),
    .A2(_04890_),
    .B1(_05720_),
    .C1(_04879_),
    .X(_05786_));
 sky130_fd_sc_hd__a211o_1 _08089_ (.A1(_04901_),
    .A2(_03588_),
    .B1(_04868_),
    .C1(_05731_),
    .X(_05797_));
 sky130_fd_sc_hd__nand4_2 _08090_ (.A(_05687_),
    .B(_05698_),
    .C(_05775_),
    .D(_05797_),
    .Y(_05807_));
 sky130_fd_sc_hd__o21ai_1 _08091_ (.A1(_05764_),
    .A2(_05786_),
    .B1(_05709_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _08092_ (.A(_05709_),
    .B(_05797_),
    .Y(_05829_));
 sky130_fd_sc_hd__o211a_2 _08093_ (.A1(_05764_),
    .A2(_05786_),
    .B1(_05687_),
    .C1(_05698_),
    .X(_05840_));
 sky130_fd_sc_hd__o211ai_1 _08094_ (.A1(_05764_),
    .A2(_05786_),
    .B1(_05687_),
    .C1(_05698_),
    .Y(_05851_));
 sky130_fd_sc_hd__a31o_1 _08095_ (.A1(_04430_),
    .A2(_04912_),
    .A3(_04923_),
    .B1(_04409_),
    .X(_05862_));
 sky130_fd_sc_hd__a31oi_2 _08096_ (.A1(_04430_),
    .A2(_04912_),
    .A3(_04923_),
    .B1(_04409_),
    .Y(_05873_));
 sky130_fd_sc_hd__nand3_4 _08097_ (.A(_05807_),
    .B(_05818_),
    .C(_05873_),
    .Y(_05884_));
 sky130_fd_sc_hd__a31o_2 _08098_ (.A1(_05709_),
    .A2(_05775_),
    .A3(_05797_),
    .B1(_05873_),
    .X(_05895_));
 sky130_fd_sc_hd__o211ai_2 _08099_ (.A1(_05764_),
    .A2(_05829_),
    .B1(_05851_),
    .C1(_05862_),
    .Y(_05906_));
 sky130_fd_sc_hd__a22o_1 _08100_ (.A1(_00867_),
    .A2(_00889_),
    .B1(_04201_),
    .B2(_04212_),
    .X(_05917_));
 sky130_fd_sc_hd__nor3_1 _08101_ (.A(_01292_),
    .B(_03906_),
    .C(_04518_),
    .Y(_05928_));
 sky130_fd_sc_hd__or3_2 _08102_ (.A(_01292_),
    .B(_03906_),
    .C(_04518_),
    .X(_05939_));
 sky130_fd_sc_hd__o32a_2 _08103_ (.A1(_01488_),
    .A2(_02122_),
    .A3(_04474_),
    .B1(_03906_),
    .B2(_01292_),
    .X(_05949_));
 sky130_fd_sc_hd__o21ai_1 _08104_ (.A1(_01292_),
    .A2(_03906_),
    .B1(_04518_),
    .Y(_05960_));
 sky130_fd_sc_hd__o22a_2 _08105_ (.A1(_00900_),
    .A2(_04244_),
    .B1(_05928_),
    .B2(_05949_),
    .X(_05971_));
 sky130_fd_sc_hd__and4_2 _08106_ (.A(_00911_),
    .B(_04255_),
    .C(_05939_),
    .D(_05960_),
    .X(_05982_));
 sky130_fd_sc_hd__and3_1 _08107_ (.A(_05917_),
    .B(_05939_),
    .C(_05960_),
    .X(_05993_));
 sky130_fd_sc_hd__o211a_1 _08108_ (.A1(_05928_),
    .A2(_05949_),
    .B1(_00911_),
    .C1(_04255_),
    .X(_06004_));
 sky130_fd_sc_hd__nor2_1 _08109_ (.A(_05971_),
    .B(_05982_),
    .Y(_06015_));
 sky130_fd_sc_hd__o2bb2ai_2 _08110_ (.A1_N(_05884_),
    .A2_N(_05906_),
    .B1(_05971_),
    .B2(_05982_),
    .Y(_06026_));
 sky130_fd_sc_hd__o221ai_4 _08111_ (.A1(_05993_),
    .A2(_06004_),
    .B1(_05840_),
    .B2(_05895_),
    .C1(_05884_),
    .Y(_06037_));
 sky130_fd_sc_hd__o221ai_4 _08112_ (.A1(_05971_),
    .A2(_05982_),
    .B1(_05840_),
    .B2(_05895_),
    .C1(_05884_),
    .Y(_06048_));
 sky130_fd_sc_hd__o2bb2ai_1 _08113_ (.A1_N(_05884_),
    .A2_N(_05906_),
    .B1(_05993_),
    .B2(_06004_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_2 _08114_ (.A(_06026_),
    .B(_06037_),
    .Y(_06070_));
 sky130_fd_sc_hd__o31a_2 _08115_ (.A1(_04299_),
    .A2(_04310_),
    .A3(_05032_),
    .B1(_05021_),
    .X(_06081_));
 sky130_fd_sc_hd__nand3_4 _08116_ (.A(_06048_),
    .B(_06059_),
    .C(_06081_),
    .Y(_06091_));
 sky130_fd_sc_hd__o211ai_4 _08117_ (.A1(_05010_),
    .A2(_05054_),
    .B1(_06026_),
    .C1(_06037_),
    .Y(_06102_));
 sky130_fd_sc_hd__o211ai_4 _08118_ (.A1(_03303_),
    .A2(_04070_),
    .B1(_05142_),
    .C1(_05164_),
    .Y(_06113_));
 sky130_fd_sc_hd__o211ai_2 _08119_ (.A1(_03292_),
    .A2(_04081_),
    .B1(_05153_),
    .C1(_05174_),
    .Y(_06124_));
 sky130_fd_sc_hd__o2111ai_4 _08120_ (.A1(_04179_),
    .A2(_05120_),
    .B1(_06091_),
    .C1(_06102_),
    .D1(_06113_),
    .Y(_06135_));
 sky130_fd_sc_hd__a22o_1 _08121_ (.A1(_06091_),
    .A2(_06102_),
    .B1(_06113_),
    .B2(_05153_),
    .X(_06146_));
 sky130_fd_sc_hd__nand4_2 _08122_ (.A(_05436_),
    .B(_06135_),
    .C(_06146_),
    .D(net1),
    .Y(_06157_));
 sky130_fd_sc_hd__a22oi_1 _08123_ (.A1(_05436_),
    .A2(net1),
    .B1(_06146_),
    .B2(_06135_),
    .Y(_06168_));
 sky130_fd_sc_hd__a32o_1 _08124_ (.A1(net1),
    .A2(_05392_),
    .A3(_05414_),
    .B1(_06135_),
    .B2(_06146_),
    .X(_06179_));
 sky130_fd_sc_hd__o211ai_2 _08125_ (.A1(_00310_),
    .A2(_05327_),
    .B1(_06157_),
    .C1(_06179_),
    .Y(_06190_));
 sky130_fd_sc_hd__a221o_1 _08126_ (.A1(_05294_),
    .A2(_05305_),
    .B1(_06157_),
    .B2(_06179_),
    .C1(_00310_),
    .X(_06201_));
 sky130_fd_sc_hd__and2_1 _08127_ (.A(_06190_),
    .B(_06201_),
    .X(_06212_));
 sky130_fd_sc_hd__xnor2_1 _08128_ (.A(_05250_),
    .B(_06212_),
    .Y(net127));
 sky130_fd_sc_hd__nand4_2 _08129_ (.A(_06201_),
    .B(_05207_),
    .C(_04157_),
    .D(_06190_),
    .Y(_06232_));
 sky130_fd_sc_hd__a21oi_2 _08130_ (.A1(_05337_),
    .A2(_06157_),
    .B1(_06168_),
    .Y(_06243_));
 sky130_fd_sc_hd__nor3_4 _08131_ (.A(net62),
    .B(net63),
    .C(_04616_),
    .Y(_06254_));
 sky130_fd_sc_hd__o311a_4 _08132_ (.A1(net62),
    .A2(net63),
    .A3(_04616_),
    .B1(_00474_),
    .C1(net173),
    .X(_06265_));
 sky130_fd_sc_hd__a311o_4 _08133_ (.A1(_04606_),
    .A2(_00463_),
    .A3(_00441_),
    .B1(_00299_),
    .C1(net64),
    .X(_06276_));
 sky130_fd_sc_hd__o21a_4 _08134_ (.A1(_00299_),
    .A2(_06254_),
    .B1(net64),
    .X(_06287_));
 sky130_fd_sc_hd__o21ai_4 _08135_ (.A1(_00299_),
    .A2(_06254_),
    .B1(net64),
    .Y(_06298_));
 sky130_fd_sc_hd__a311o_4 _08136_ (.A1(_04606_),
    .A2(_00463_),
    .A3(_00441_),
    .B1(_00299_),
    .C1(_00474_),
    .X(_06309_));
 sky130_fd_sc_hd__o21ai_4 _08137_ (.A1(_00299_),
    .A2(_06254_),
    .B1(_00474_),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_8 _08138_ (.A(_06309_),
    .B(_06320_),
    .Y(_06331_));
 sky130_fd_sc_hd__nand2_8 _08139_ (.A(_06276_),
    .B(_06298_),
    .Y(_06341_));
 sky130_fd_sc_hd__o21ai_1 _08140_ (.A1(_06265_),
    .A2(_06287_),
    .B1(net1),
    .Y(_06352_));
 sky130_fd_sc_hd__and4_2 _08141_ (.A(_00998_),
    .B(_05436_),
    .C(_06341_),
    .D(net1),
    .X(_06363_));
 sky130_fd_sc_hd__or4_1 _08142_ (.A(_00987_),
    .B(_05381_),
    .C(_05403_),
    .D(_06352_),
    .X(_06374_));
 sky130_fd_sc_hd__o32a_2 _08143_ (.A1(_00987_),
    .A2(_05381_),
    .A3(_05403_),
    .B1(_00288_),
    .B2(_06331_),
    .X(_06385_));
 sky130_fd_sc_hd__nor2_1 _08144_ (.A(_06363_),
    .B(_06385_),
    .Y(_06396_));
 sky130_fd_sc_hd__o21ai_1 _08145_ (.A1(_05993_),
    .A2(_06004_),
    .B1(_05884_),
    .Y(_06407_));
 sky130_fd_sc_hd__o2bb2ai_1 _08146_ (.A1_N(_06015_),
    .A2_N(_05884_),
    .B1(_05840_),
    .B2(_05895_),
    .Y(_06418_));
 sky130_fd_sc_hd__a31oi_2 _08147_ (.A1(_05687_),
    .A2(_05698_),
    .A3(_05775_),
    .B1(_05786_),
    .Y(_06429_));
 sky130_fd_sc_hd__and3_1 _08148_ (.A(_00911_),
    .B(_04255_),
    .C(_05960_),
    .X(_06440_));
 sky130_fd_sc_hd__a31oi_1 _08149_ (.A1(_00911_),
    .A2(_04255_),
    .A3(_05960_),
    .B1(_05928_),
    .Y(_06451_));
 sky130_fd_sc_hd__nand2_1 _08150_ (.A(_05654_),
    .B(_05676_),
    .Y(_06461_));
 sky130_fd_sc_hd__o211ai_2 _08151_ (.A1(_04551_),
    .A2(_04781_),
    .B1(_05644_),
    .C1(_04770_),
    .Y(_06472_));
 sky130_fd_sc_hd__o211a_1 _08152_ (.A1(_05928_),
    .A2(_06440_),
    .B1(_06461_),
    .C1(_05644_),
    .X(_06483_));
 sky130_fd_sc_hd__nand3b_2 _08153_ (.A_N(_06451_),
    .B(_06461_),
    .C(_05644_),
    .Y(_06494_));
 sky130_fd_sc_hd__o2111ai_4 _08154_ (.A1(_05949_),
    .A2(_05917_),
    .B1(_05654_),
    .C1(_05939_),
    .D1(_06472_),
    .Y(_06505_));
 sky130_fd_sc_hd__o21ai_1 _08155_ (.A1(_04584_),
    .A2(_05545_),
    .B1(_05589_),
    .Y(_06516_));
 sky130_fd_sc_hd__nand2_1 _08156_ (.A(_05534_),
    .B(_06516_),
    .Y(_06527_));
 sky130_fd_sc_hd__a22oi_4 _08157_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_05556_),
    .B2(_05589_),
    .Y(_06538_));
 sky130_fd_sc_hd__o211a_1 _08158_ (.A1(net169),
    .A2(net163),
    .B1(_01936_),
    .C1(_01947_),
    .X(_06549_));
 sky130_fd_sc_hd__nand4_1 _08159_ (.A(_01936_),
    .B(_01947_),
    .C(_02822_),
    .D(_02844_),
    .Y(_06559_));
 sky130_fd_sc_hd__a32oi_1 _08160_ (.A1(net173),
    .A2(net61),
    .A3(_03413_),
    .B1(_01455_),
    .B2(_01434_),
    .Y(_06570_));
 sky130_fd_sc_hd__o221ai_4 _08161_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_03511_),
    .B2(_00299_),
    .C1(_03490_),
    .Y(_06581_));
 sky130_fd_sc_hd__o32a_1 _08162_ (.A1(net165),
    .A2(_04671_),
    .A3(_04693_),
    .B1(_01488_),
    .B2(_03544_),
    .X(_06592_));
 sky130_fd_sc_hd__nand2_1 _08163_ (.A(_05545_),
    .B(_06581_),
    .Y(_06603_));
 sky130_fd_sc_hd__nand4_2 _08164_ (.A(_06570_),
    .B(_04704_),
    .C(_04682_),
    .D(_03490_),
    .Y(_06614_));
 sky130_fd_sc_hd__o21ai_1 _08165_ (.A1(net165),
    .A2(_06614_),
    .B1(_06603_),
    .Y(_06625_));
 sky130_fd_sc_hd__o21ai_2 _08166_ (.A1(_01958_),
    .A2(net159),
    .B1(_06625_),
    .Y(_06636_));
 sky130_fd_sc_hd__o21ai_2 _08167_ (.A1(_05545_),
    .A2(_06581_),
    .B1(_06549_),
    .Y(_06647_));
 sky130_fd_sc_hd__nand2_1 _08168_ (.A(_06625_),
    .B(_06549_),
    .Y(_06658_));
 sky130_fd_sc_hd__o221ai_4 _08169_ (.A1(_01958_),
    .A2(net159),
    .B1(net165),
    .B2(_06614_),
    .C1(_06603_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand3_4 _08170_ (.A(_06658_),
    .B(_06668_),
    .C(_06527_),
    .Y(_06679_));
 sky130_fd_sc_hd__o211a_1 _08171_ (.A1(_06647_),
    .A2(_06592_),
    .B1(_06538_),
    .C1(_06636_),
    .X(_06690_));
 sky130_fd_sc_hd__o211ai_4 _08172_ (.A1(_06647_),
    .A2(_06592_),
    .B1(_06538_),
    .C1(_06636_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand3_2 _08173_ (.A(_06679_),
    .B(_06701_),
    .C(_05458_),
    .Y(_06712_));
 sky130_fd_sc_hd__a32o_1 _08174_ (.A1(_02133_),
    .A2(_04463_),
    .A3(_02647_),
    .B1(_06701_),
    .B2(_06679_),
    .X(_06723_));
 sky130_fd_sc_hd__a21oi_2 _08175_ (.A1(_06679_),
    .A2(_06701_),
    .B1(_05469_),
    .Y(_06734_));
 sky130_fd_sc_hd__a21o_1 _08176_ (.A1(_06679_),
    .A2(_06701_),
    .B1(_05469_),
    .X(_06745_));
 sky130_fd_sc_hd__o21ai_2 _08177_ (.A1(_04474_),
    .A2(_05447_),
    .B1(_06679_),
    .Y(_06755_));
 sky130_fd_sc_hd__o311a_1 _08178_ (.A1(_02122_),
    .A2(_02636_),
    .A3(_04474_),
    .B1(_06679_),
    .C1(_06701_),
    .X(_06766_));
 sky130_fd_sc_hd__o2111ai_4 _08179_ (.A1(_06690_),
    .A2(_06755_),
    .B1(_06745_),
    .C1(_06494_),
    .D1(_06505_),
    .Y(_06777_));
 sky130_fd_sc_hd__o2bb2ai_1 _08180_ (.A1_N(_06494_),
    .A2_N(_06505_),
    .B1(_06734_),
    .B2(_06766_),
    .Y(_06788_));
 sky130_fd_sc_hd__o2bb2ai_1 _08181_ (.A1_N(_06494_),
    .A2_N(_06505_),
    .B1(_06690_),
    .B2(_06755_),
    .Y(_06799_));
 sky130_fd_sc_hd__nand4_2 _08182_ (.A(_06494_),
    .B(_06505_),
    .C(_06712_),
    .D(_06723_),
    .Y(_06810_));
 sky130_fd_sc_hd__nand4_4 _08183_ (.A(_05775_),
    .B(_05829_),
    .C(_06777_),
    .D(_06788_),
    .Y(_06821_));
 sky130_fd_sc_hd__o211ai_4 _08184_ (.A1(_06734_),
    .A2(_06799_),
    .B1(_06810_),
    .C1(_06429_),
    .Y(_06832_));
 sky130_fd_sc_hd__a32o_2 _08185_ (.A1(_02133_),
    .A2(_02614_),
    .A3(_02625_),
    .B1(_03917_),
    .B2(_01631_),
    .X(_06842_));
 sky130_fd_sc_hd__or4_4 _08186_ (.A(_01620_),
    .B(_02122_),
    .C(_02636_),
    .D(_03906_),
    .X(_06853_));
 sky130_fd_sc_hd__a22oi_2 _08187_ (.A1(_01303_),
    .A2(_04255_),
    .B1(_06842_),
    .B2(_06853_),
    .Y(_06864_));
 sky130_fd_sc_hd__and4_1 _08188_ (.A(_01303_),
    .B(_04255_),
    .C(_06842_),
    .D(_06853_),
    .X(_06875_));
 sky130_fd_sc_hd__a211oi_1 _08189_ (.A1(_06842_),
    .A2(_06853_),
    .B1(_01292_),
    .C1(_04244_),
    .Y(_06886_));
 sky130_fd_sc_hd__o211a_1 _08190_ (.A1(_01292_),
    .A2(_04244_),
    .B1(_06842_),
    .C1(_06853_),
    .X(_06897_));
 sky130_fd_sc_hd__nor2_1 _08191_ (.A(_06886_),
    .B(_06897_),
    .Y(_06908_));
 sky130_fd_sc_hd__o211ai_2 _08192_ (.A1(_06886_),
    .A2(_06897_),
    .B1(_06821_),
    .C1(_06832_),
    .Y(_06919_));
 sky130_fd_sc_hd__o2bb2ai_1 _08193_ (.A1_N(_06821_),
    .A2_N(_06832_),
    .B1(_06864_),
    .B2(_06875_),
    .Y(_06929_));
 sky130_fd_sc_hd__a21oi_4 _08194_ (.A1(_06821_),
    .A2(_06832_),
    .B1(_06908_),
    .Y(_06940_));
 sky130_fd_sc_hd__o211ai_2 _08195_ (.A1(_06864_),
    .A2(_06875_),
    .B1(_06821_),
    .C1(_06832_),
    .Y(_06951_));
 sky130_fd_sc_hd__o211ai_4 _08196_ (.A1(_05840_),
    .A2(_05895_),
    .B1(_06407_),
    .C1(_06951_),
    .Y(_06962_));
 sky130_fd_sc_hd__nand3_4 _08197_ (.A(_06929_),
    .B(_06418_),
    .C(_06919_),
    .Y(_06973_));
 sky130_fd_sc_hd__o21a_1 _08198_ (.A1(_06940_),
    .A2(_06962_),
    .B1(_06973_),
    .X(_06984_));
 sky130_fd_sc_hd__o21ai_1 _08199_ (.A1(_06940_),
    .A2(_06962_),
    .B1(_06973_),
    .Y(_06995_));
 sky130_fd_sc_hd__o211ai_4 _08200_ (.A1(_05065_),
    .A2(_05131_),
    .B1(_06102_),
    .C1(_06124_),
    .Y(_07005_));
 sky130_fd_sc_hd__o211ai_4 _08201_ (.A1(_04179_),
    .A2(_05120_),
    .B1(_06091_),
    .C1(_06113_),
    .Y(_07016_));
 sky130_fd_sc_hd__nand3_1 _08202_ (.A(_06984_),
    .B(_07005_),
    .C(_06091_),
    .Y(_07027_));
 sky130_fd_sc_hd__o211ai_2 _08203_ (.A1(_06070_),
    .A2(_06081_),
    .B1(_06995_),
    .C1(_07016_),
    .Y(_07038_));
 sky130_fd_sc_hd__o211ai_2 _08204_ (.A1(_06070_),
    .A2(_06081_),
    .B1(_07016_),
    .C1(_06984_),
    .Y(_07049_));
 sky130_fd_sc_hd__nand3_1 _08205_ (.A(_06091_),
    .B(_06995_),
    .C(_07005_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand3_1 _08206_ (.A(_07027_),
    .B(_07038_),
    .C(_06396_),
    .Y(_07070_));
 sky130_fd_sc_hd__o211ai_4 _08207_ (.A1(_06363_),
    .A2(_06385_),
    .B1(_07049_),
    .C1(_07060_),
    .Y(_07081_));
 sky130_fd_sc_hd__nor2_2 _08208_ (.A(net30),
    .B(net31),
    .Y(_07092_));
 sky130_fd_sc_hd__nand4_4 _08209_ (.A(net171),
    .B(_03840_),
    .C(_07092_),
    .D(_00430_),
    .Y(_07103_));
 sky130_fd_sc_hd__a41o_2 _08210_ (.A1(net171),
    .A2(_03840_),
    .A3(_07092_),
    .A4(_00430_),
    .B1(_00321_),
    .X(_07114_));
 sky130_fd_sc_hd__o311a_4 _08211_ (.A1(net30),
    .A2(net31),
    .A3(_04190_),
    .B1(_00485_),
    .C1(net174),
    .X(_07125_));
 sky130_fd_sc_hd__a21oi_4 _08212_ (.A1(_07103_),
    .A2(net174),
    .B1(_00485_),
    .Y(_07135_));
 sky130_fd_sc_hd__and3_4 _08213_ (.A(_07103_),
    .B(net32),
    .C(net174),
    .X(_07146_));
 sky130_fd_sc_hd__o211ai_4 _08214_ (.A1(net31),
    .A2(_05261_),
    .B1(net32),
    .C1(net174),
    .Y(_07157_));
 sky130_fd_sc_hd__a21oi_4 _08215_ (.A1(_07103_),
    .A2(net174),
    .B1(net32),
    .Y(_07168_));
 sky130_fd_sc_hd__a21o_4 _08216_ (.A1(_07103_),
    .A2(net174),
    .B1(net32),
    .X(_07178_));
 sky130_fd_sc_hd__nand2_8 _08217_ (.A(_07157_),
    .B(_07178_),
    .Y(_07189_));
 sky130_fd_sc_hd__nor2_8 _08218_ (.A(_07146_),
    .B(_07168_),
    .Y(_07200_));
 sky130_fd_sc_hd__or3_1 _08219_ (.A(_00900_),
    .B(_07146_),
    .C(_07168_),
    .X(_07211_));
 sky130_fd_sc_hd__and4_1 _08220_ (.A(_00911_),
    .B(_07200_),
    .C(_05316_),
    .D(net33),
    .X(_07222_));
 sky130_fd_sc_hd__o32a_1 _08221_ (.A1(_00310_),
    .A2(_07146_),
    .A3(_07168_),
    .B1(_00900_),
    .B2(_05327_),
    .X(_07232_));
 sky130_fd_sc_hd__nor2_1 _08222_ (.A(_07222_),
    .B(_07232_),
    .Y(_07243_));
 sky130_fd_sc_hd__o2bb2ai_1 _08223_ (.A1_N(_07070_),
    .A2_N(_07081_),
    .B1(_07222_),
    .B2(_07232_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand3_1 _08224_ (.A(_07070_),
    .B(_07081_),
    .C(_07243_),
    .Y(_07264_));
 sky130_fd_sc_hd__nand2_1 _08225_ (.A(_07254_),
    .B(_07264_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand3_2 _08226_ (.A(_06243_),
    .B(_07254_),
    .C(_07264_),
    .Y(_07286_));
 sky130_fd_sc_hd__xnor2_2 _08227_ (.A(_06243_),
    .B(_07275_),
    .Y(_07296_));
 sky130_fd_sc_hd__a21oi_1 _08228_ (.A1(_00845_),
    .A2(_06232_),
    .B1(_07296_),
    .Y(_07307_));
 sky130_fd_sc_hd__and3_1 _08229_ (.A(_00845_),
    .B(_06232_),
    .C(_07296_),
    .X(_07318_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(_07307_),
    .B(_07318_),
    .Y(net128));
 sky130_fd_sc_hd__o21ai_1 _08231_ (.A1(_07296_),
    .A2(_06232_),
    .B1(_00845_),
    .Y(_07338_));
 sky130_fd_sc_hd__a32oi_4 _08232_ (.A1(_06396_),
    .A2(_07027_),
    .A3(_07038_),
    .B1(_07081_),
    .B2(_07243_),
    .Y(_07348_));
 sky130_fd_sc_hd__nand4b_4 _08233_ (.A_N(_04616_),
    .B(_00474_),
    .C(_00463_),
    .D(_00441_),
    .Y(_07358_));
 sky130_fd_sc_hd__o41a_1 _08234_ (.A1(net62),
    .A2(net63),
    .A3(net64),
    .A4(_04616_),
    .B1(net34),
    .X(_07365_));
 sky130_fd_sc_hd__nand2_1 _08235_ (.A(_07358_),
    .B(net34),
    .Y(_07366_));
 sky130_fd_sc_hd__a21oi_2 _08236_ (.A1(_07358_),
    .A2(net173),
    .B1(net34),
    .Y(_07367_));
 sky130_fd_sc_hd__a21o_1 _08237_ (.A1(_07358_),
    .A2(net57),
    .B1(net34),
    .X(_07368_));
 sky130_fd_sc_hd__o21ai_4 _08238_ (.A1(_00299_),
    .A2(_07366_),
    .B1(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__a21oi_4 _08239_ (.A1(net173),
    .A2(_07365_),
    .B1(_07367_),
    .Y(_07370_));
 sky130_fd_sc_hd__a221o_1 _08240_ (.A1(_00932_),
    .A2(_00954_),
    .B1(_07365_),
    .B2(net173),
    .C1(_07367_),
    .X(_07371_));
 sky130_fd_sc_hd__and4_1 _08241_ (.A(_00998_),
    .B(_06341_),
    .C(_07370_),
    .D(net1),
    .X(_07372_));
 sky130_fd_sc_hd__o22a_1 _08242_ (.A1(_00987_),
    .A2(_06331_),
    .B1(_00288_),
    .B2(net153),
    .X(_07373_));
 sky130_fd_sc_hd__o32a_1 _08243_ (.A1(net165),
    .A2(_05381_),
    .A3(_05403_),
    .B1(_07372_),
    .B2(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__a211oi_2 _08244_ (.A1(_01106_),
    .A2(_01128_),
    .B1(_07372_),
    .C1(_07373_),
    .Y(_07375_));
 sky130_fd_sc_hd__a31o_1 _08245_ (.A1(_07375_),
    .A2(_05414_),
    .A3(_05392_),
    .B1(_07374_),
    .X(_07376_));
 sky130_fd_sc_hd__o31a_1 _08246_ (.A1(_00987_),
    .A2(_05425_),
    .A3(_06352_),
    .B1(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__a211oi_2 _08247_ (.A1(_07375_),
    .A2(_05436_),
    .B1(_06374_),
    .C1(_07374_),
    .Y(_07378_));
 sky130_fd_sc_hd__nor2_1 _08248_ (.A(_07377_),
    .B(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__a31o_1 _08249_ (.A1(_06505_),
    .A2(_06712_),
    .A3(_06723_),
    .B1(_06483_),
    .X(_07380_));
 sky130_fd_sc_hd__a31oi_2 _08250_ (.A1(_06505_),
    .A2(_06712_),
    .A3(_06723_),
    .B1(_06483_),
    .Y(_07381_));
 sky130_fd_sc_hd__o211ai_2 _08251_ (.A1(_01238_),
    .A2(_01249_),
    .B1(_04255_),
    .C1(_06842_),
    .Y(_07382_));
 sky130_fd_sc_hd__nand2_1 _08252_ (.A(_06853_),
    .B(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__o21ai_1 _08253_ (.A1(_04474_),
    .A2(_05447_),
    .B1(_06701_),
    .Y(_07384_));
 sky130_fd_sc_hd__nand2_1 _08254_ (.A(_06679_),
    .B(_05458_),
    .Y(_07385_));
 sky130_fd_sc_hd__a22oi_2 _08255_ (.A1(_06853_),
    .A2(_07382_),
    .B1(_07385_),
    .B2(_06701_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand3_1 _08256_ (.A(_06679_),
    .B(_07383_),
    .C(_07384_),
    .Y(_07387_));
 sky130_fd_sc_hd__a211oi_1 _08257_ (.A1(_05458_),
    .A2(_06679_),
    .B1(_07383_),
    .C1(_06690_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand3b_2 _08258_ (.A_N(_07383_),
    .B(_07385_),
    .C(_06701_),
    .Y(_07389_));
 sky130_fd_sc_hd__a221o_1 _08259_ (.A1(_01903_),
    .A2(_01925_),
    .B1(_03501_),
    .B2(net173),
    .C1(_03479_),
    .X(_07390_));
 sky130_fd_sc_hd__o221a_1 _08260_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_04606_),
    .B2(_04660_),
    .C1(_04704_),
    .X(_07391_));
 sky130_fd_sc_hd__a211o_1 _08261_ (.A1(_01434_),
    .A2(_01455_),
    .B1(_04671_),
    .C1(_04693_),
    .X(_07392_));
 sky130_fd_sc_hd__a21oi_2 _08262_ (.A1(_05545_),
    .A2(_06581_),
    .B1(_06559_),
    .Y(_07393_));
 sky130_fd_sc_hd__o21bai_4 _08263_ (.A1(_05512_),
    .A2(_07393_),
    .B1_N(_07392_),
    .Y(_07394_));
 sky130_fd_sc_hd__a32o_1 _08264_ (.A1(_01499_),
    .A2(_04682_),
    .A3(_04704_),
    .B1(_06603_),
    .B2(_06549_),
    .X(_07395_));
 sky130_fd_sc_hd__a22oi_2 _08265_ (.A1(_01969_),
    .A2(net157),
    .B1(_07394_),
    .B2(_07395_),
    .Y(_07396_));
 sky130_fd_sc_hd__o21bai_2 _08266_ (.A1(_07391_),
    .A2(_07393_),
    .B1_N(_07390_),
    .Y(_07397_));
 sky130_fd_sc_hd__a41oi_4 _08267_ (.A1(_01969_),
    .A2(net157),
    .A3(_07394_),
    .A4(_07395_),
    .B1(_07396_),
    .Y(_07398_));
 sky130_fd_sc_hd__a41o_1 _08268_ (.A1(_01969_),
    .A2(net157),
    .A3(_07394_),
    .A4(_07395_),
    .B1(_07396_),
    .X(_07399_));
 sky130_fd_sc_hd__nand3_1 _08269_ (.A(_07387_),
    .B(_07389_),
    .C(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__o21ai_1 _08270_ (.A1(_07386_),
    .A2(_07388_),
    .B1(_07398_),
    .Y(_07401_));
 sky130_fd_sc_hd__o21ai_1 _08271_ (.A1(_07386_),
    .A2(_07388_),
    .B1(_07399_),
    .Y(_07402_));
 sky130_fd_sc_hd__nand3_1 _08272_ (.A(_07387_),
    .B(_07389_),
    .C(_07398_),
    .Y(_07403_));
 sky130_fd_sc_hd__nand3_2 _08273_ (.A(_07381_),
    .B(_07400_),
    .C(_07401_),
    .Y(_07404_));
 sky130_fd_sc_hd__nand3_2 _08274_ (.A(_07380_),
    .B(_07402_),
    .C(_07403_),
    .Y(_07405_));
 sky130_fd_sc_hd__a22o_1 _08275_ (.A1(_01543_),
    .A2(_01565_),
    .B1(_04201_),
    .B2(_04212_),
    .X(_07406_));
 sky130_fd_sc_hd__o22a_1 _08276_ (.A1(_02636_),
    .A2(net159),
    .B1(_03906_),
    .B2(_02122_),
    .X(_07407_));
 sky130_fd_sc_hd__o211a_1 _08277_ (.A1(net169),
    .A2(_02800_),
    .B1(_03884_),
    .C1(_03895_),
    .X(_07408_));
 sky130_fd_sc_hd__and3_1 _08278_ (.A(_07408_),
    .B(_02647_),
    .C(_02133_),
    .X(_07409_));
 sky130_fd_sc_hd__o32a_1 _08279_ (.A1(_01576_),
    .A2(_01598_),
    .A3(_04244_),
    .B1(_07407_),
    .B2(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__a311oi_2 _08280_ (.A1(_02133_),
    .A2(_02647_),
    .A3(_07408_),
    .B1(_07406_),
    .C1(_07407_),
    .Y(_07411_));
 sky130_fd_sc_hd__or2_1 _08281_ (.A(_07410_),
    .B(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__a21bo_1 _08282_ (.A1(_07404_),
    .A2(_07405_),
    .B1_N(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__nand3b_1 _08283_ (.A_N(_07412_),
    .B(_07405_),
    .C(_07404_),
    .Y(_07414_));
 sky130_fd_sc_hd__o211ai_2 _08284_ (.A1(_07410_),
    .A2(_07411_),
    .B1(_07404_),
    .C1(_07405_),
    .Y(_07415_));
 sky130_fd_sc_hd__a21o_1 _08285_ (.A1(_07404_),
    .A2(_07405_),
    .B1(_07412_),
    .X(_07416_));
 sky130_fd_sc_hd__nand2_2 _08286_ (.A(_07413_),
    .B(_07414_),
    .Y(_07417_));
 sky130_fd_sc_hd__a21bo_2 _08287_ (.A1(_06832_),
    .A2(_06908_),
    .B1_N(_06821_),
    .X(_07418_));
 sky130_fd_sc_hd__a21boi_1 _08288_ (.A1(_06832_),
    .A2(_06908_),
    .B1_N(_06821_),
    .Y(_07419_));
 sky130_fd_sc_hd__nand3_4 _08289_ (.A(_07418_),
    .B(_07416_),
    .C(_07415_),
    .Y(_07420_));
 sky130_fd_sc_hd__nand3_2 _08290_ (.A(_07413_),
    .B(_07414_),
    .C(_07419_),
    .Y(_07421_));
 sky130_fd_sc_hd__and2_1 _08291_ (.A(_07420_),
    .B(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__nand2_1 _08292_ (.A(_07420_),
    .B(_07421_),
    .Y(_07423_));
 sky130_fd_sc_hd__o211ai_4 _08293_ (.A1(_06070_),
    .A2(_06081_),
    .B1(_06973_),
    .C1(_07016_),
    .Y(_07424_));
 sky130_fd_sc_hd__o211ai_4 _08294_ (.A1(_06962_),
    .A2(_06940_),
    .B1(_06091_),
    .C1(_07005_),
    .Y(_07425_));
 sky130_fd_sc_hd__o211ai_2 _08295_ (.A1(_06940_),
    .A2(_06962_),
    .B1(_07423_),
    .C1(_07424_),
    .Y(_07426_));
 sky130_fd_sc_hd__nand3_1 _08296_ (.A(_06973_),
    .B(_07425_),
    .C(_07422_),
    .Y(_07427_));
 sky130_fd_sc_hd__o211ai_2 _08297_ (.A1(_06940_),
    .A2(_06962_),
    .B1(_07422_),
    .C1(_07424_),
    .Y(_07428_));
 sky130_fd_sc_hd__nand3_1 _08298_ (.A(_06973_),
    .B(_07423_),
    .C(_07425_),
    .Y(_07429_));
 sky130_fd_sc_hd__o211a_1 _08299_ (.A1(_07377_),
    .A2(_07378_),
    .B1(_07426_),
    .C1(_07427_),
    .X(_07430_));
 sky130_fd_sc_hd__o211ai_2 _08300_ (.A1(_07377_),
    .A2(_07378_),
    .B1(_07426_),
    .C1(_07427_),
    .Y(_07431_));
 sky130_fd_sc_hd__nand3_4 _08301_ (.A(_07429_),
    .B(_07379_),
    .C(_07428_),
    .Y(_07432_));
 sky130_fd_sc_hd__nor3_2 _08302_ (.A(net30),
    .B(net31),
    .C(net32),
    .Y(_07433_));
 sky130_fd_sc_hd__nand2_8 _08303_ (.A(_07092_),
    .B(_00485_),
    .Y(_07434_));
 sky130_fd_sc_hd__nor3_4 _08304_ (.A(_07434_),
    .B(net29),
    .C(_03851_),
    .Y(_07435_));
 sky130_fd_sc_hd__o211ai_4 _08305_ (.A1(_04190_),
    .A2(_07434_),
    .B1(net174),
    .C1(net2),
    .Y(_07436_));
 sky130_fd_sc_hd__o21ai_4 _08306_ (.A1(_00321_),
    .A2(_07435_),
    .B1(_00496_),
    .Y(_07437_));
 sky130_fd_sc_hd__o211ai_4 _08307_ (.A1(_04190_),
    .A2(_07434_),
    .B1(net174),
    .C1(_00496_),
    .Y(_07438_));
 sky130_fd_sc_hd__o21ai_4 _08308_ (.A1(_00321_),
    .A2(_07435_),
    .B1(net2),
    .Y(_07439_));
 sky130_fd_sc_hd__nand2_8 _08309_ (.A(_07438_),
    .B(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__nand2_8 _08310_ (.A(_07436_),
    .B(net154),
    .Y(_07441_));
 sky130_fd_sc_hd__a32o_1 _08311_ (.A1(_00911_),
    .A2(_07157_),
    .A3(_07178_),
    .B1(_05316_),
    .B2(_01303_),
    .X(_07442_));
 sky130_fd_sc_hd__a21oi_2 _08312_ (.A1(_00485_),
    .A2(_07114_),
    .B1(_01292_),
    .Y(_07443_));
 sky130_fd_sc_hd__o211ai_4 _08313_ (.A1(_01238_),
    .A2(_01249_),
    .B1(_07157_),
    .C1(_07178_),
    .Y(_07444_));
 sky130_fd_sc_hd__and4_1 _08314_ (.A(_05316_),
    .B(_07443_),
    .C(_07157_),
    .D(_00911_),
    .X(_07445_));
 sky130_fd_sc_hd__or4_1 _08315_ (.A(_00900_),
    .B(_01292_),
    .C(_05327_),
    .D(_07189_),
    .X(_07446_));
 sky130_fd_sc_hd__or4bb_4 _08316_ (.A(_07445_),
    .B(_07441_),
    .C_N(net33),
    .D_N(_07442_),
    .X(_07447_));
 sky130_fd_sc_hd__a32o_1 _08317_ (.A1(net33),
    .A2(net162),
    .A3(net154),
    .B1(_07442_),
    .B2(_07446_),
    .X(_07448_));
 sky130_fd_sc_hd__nand2_1 _08318_ (.A(_07447_),
    .B(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__o31a_1 _08319_ (.A1(_00900_),
    .A2(_05337_),
    .A3(_07189_),
    .B1(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__and3_1 _08320_ (.A(_07448_),
    .B(_07222_),
    .C(_07447_),
    .X(_07451_));
 sky130_fd_sc_hd__o211a_1 _08321_ (.A1(_05337_),
    .A2(_07211_),
    .B1(_07447_),
    .C1(_07448_),
    .X(_07452_));
 sky130_fd_sc_hd__and4b_1 _08322_ (.A_N(_05337_),
    .B(_07200_),
    .C(_07449_),
    .D(_00911_),
    .X(_07453_));
 sky130_fd_sc_hd__nor2_1 _08323_ (.A(_07452_),
    .B(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__o211ai_1 _08324_ (.A1(_07452_),
    .A2(_07453_),
    .B1(_07431_),
    .C1(_07432_),
    .Y(_07455_));
 sky130_fd_sc_hd__o2bb2ai_1 _08325_ (.A1_N(_07431_),
    .A2_N(_07432_),
    .B1(_07450_),
    .B2(_07451_),
    .Y(_07456_));
 sky130_fd_sc_hd__o2bb2ai_1 _08326_ (.A1_N(_07431_),
    .A2_N(_07432_),
    .B1(_07452_),
    .B2(_07453_),
    .Y(_07457_));
 sky130_fd_sc_hd__o211ai_2 _08327_ (.A1(_07450_),
    .A2(_07451_),
    .B1(_07431_),
    .C1(_07432_),
    .Y(_07458_));
 sky130_fd_sc_hd__nand2_1 _08328_ (.A(_07455_),
    .B(_07456_),
    .Y(_07459_));
 sky130_fd_sc_hd__a21oi_1 _08329_ (.A1(_07457_),
    .A2(_07458_),
    .B1(_07348_),
    .Y(_07460_));
 sky130_fd_sc_hd__nand2_1 _08330_ (.A(_07459_),
    .B(_07348_),
    .Y(_07461_));
 sky130_fd_sc_hd__nand2b_1 _08331_ (.A_N(_07460_),
    .B(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__xor2_2 _08332_ (.A(_07286_),
    .B(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__xnor2_1 _08333_ (.A(_07338_),
    .B(_07463_),
    .Y(net66));
 sky130_fd_sc_hd__o31ai_1 _08334_ (.A1(_06232_),
    .A2(_07296_),
    .A3(_07463_),
    .B1(_00845_),
    .Y(_07464_));
 sky130_fd_sc_hd__o21ai_1 _08335_ (.A1(_07454_),
    .A2(_07430_),
    .B1(_07432_),
    .Y(_07465_));
 sky130_fd_sc_hd__a32o_4 _08336_ (.A1(_07381_),
    .A2(_07400_),
    .A3(_07401_),
    .B1(_07405_),
    .B2(_07412_),
    .X(_07466_));
 sky130_fd_sc_hd__inv_2 _08337_ (.A(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__nor2_1 _08338_ (.A(_07406_),
    .B(_07407_),
    .Y(_07468_));
 sky130_fd_sc_hd__o32a_1 _08339_ (.A1(net159),
    .A2(_03906_),
    .A3(_05447_),
    .B1(_07406_),
    .B2(_07407_),
    .X(_07469_));
 sky130_fd_sc_hd__nand3_1 _08340_ (.A(_07469_),
    .B(_07397_),
    .C(_07394_),
    .Y(_07470_));
 sky130_fd_sc_hd__o2bb2ai_1 _08341_ (.A1_N(_07394_),
    .A2_N(_07397_),
    .B1(_07409_),
    .B2(_07468_),
    .Y(_07471_));
 sky130_fd_sc_hd__and4_1 _08342_ (.A(_01969_),
    .B(_02647_),
    .C(net157),
    .D(_04726_),
    .X(_07472_));
 sky130_fd_sc_hd__o32a_1 _08343_ (.A1(_01958_),
    .A2(_04671_),
    .A3(_04693_),
    .B1(_02636_),
    .B2(_03544_),
    .X(_07473_));
 sky130_fd_sc_hd__a32o_1 _08344_ (.A1(_01969_),
    .A2(_04682_),
    .A3(_04704_),
    .B1(_02647_),
    .B2(net157),
    .X(_07474_));
 sky130_fd_sc_hd__o32a_1 _08345_ (.A1(net167),
    .A2(_02833_),
    .A3(_03906_),
    .B1(_07472_),
    .B2(_07473_),
    .X(_07475_));
 sky130_fd_sc_hd__o22ai_1 _08346_ (.A1(net159),
    .A2(_03906_),
    .B1(_07472_),
    .B2(_07473_),
    .Y(_07476_));
 sky130_fd_sc_hd__o311a_1 _08347_ (.A1(_02636_),
    .A2(_04715_),
    .A3(_07390_),
    .B1(_07408_),
    .C1(_07474_),
    .X(_07477_));
 sky130_fd_sc_hd__o311ai_1 _08348_ (.A1(_02636_),
    .A2(_04715_),
    .A3(_07390_),
    .B1(_07408_),
    .C1(_07474_),
    .Y(_07478_));
 sky130_fd_sc_hd__nand2_1 _08349_ (.A(_07476_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__a21oi_1 _08350_ (.A1(_07470_),
    .A2(_07471_),
    .B1(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__o211a_1 _08351_ (.A1(_07475_),
    .A2(_07477_),
    .B1(_07470_),
    .C1(_07471_),
    .X(_07481_));
 sky130_fd_sc_hd__nor2_1 _08352_ (.A(_07480_),
    .B(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__nand2_1 _08353_ (.A(_07387_),
    .B(_07399_),
    .Y(_07483_));
 sky130_fd_sc_hd__a21oi_2 _08354_ (.A1(_07389_),
    .A2(_07398_),
    .B1(_07386_),
    .Y(_07484_));
 sky130_fd_sc_hd__o211a_1 _08355_ (.A1(_07480_),
    .A2(_07481_),
    .B1(_07483_),
    .C1(_07389_),
    .X(_07485_));
 sky130_fd_sc_hd__o211ai_2 _08356_ (.A1(_07480_),
    .A2(_07481_),
    .B1(_07483_),
    .C1(_07389_),
    .Y(_07486_));
 sky130_fd_sc_hd__nand2_1 _08357_ (.A(_07482_),
    .B(_07484_),
    .Y(_07487_));
 sky130_fd_sc_hd__a2bb2oi_1 _08358_ (.A1_N(_02122_),
    .A2_N(_04244_),
    .B1(_07486_),
    .B2(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__nand4_2 _08359_ (.A(_02133_),
    .B(_04255_),
    .C(_07486_),
    .D(_07487_),
    .Y(_07489_));
 sky130_fd_sc_hd__nand2b_4 _08360_ (.A_N(_07488_),
    .B(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__inv_2 _08361_ (.A(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__and2_1 _08362_ (.A(_07490_),
    .B(_07466_),
    .X(_07492_));
 sky130_fd_sc_hd__nor2_1 _08363_ (.A(_07466_),
    .B(_07490_),
    .Y(_07493_));
 sky130_fd_sc_hd__xor2_1 _08364_ (.A(_07466_),
    .B(_07490_),
    .X(_07494_));
 sky130_fd_sc_hd__o211ai_4 _08365_ (.A1(_07418_),
    .A2(_07417_),
    .B1(_06973_),
    .C1(_07425_),
    .Y(_07495_));
 sky130_fd_sc_hd__o211ai_4 _08366_ (.A1(_06940_),
    .A2(_06962_),
    .B1(_07420_),
    .C1(_07424_),
    .Y(_07496_));
 sky130_fd_sc_hd__o211ai_1 _08367_ (.A1(_07492_),
    .A2(_07493_),
    .B1(_07495_),
    .C1(_07420_),
    .Y(_07497_));
 sky130_fd_sc_hd__o211ai_1 _08368_ (.A1(_07417_),
    .A2(_07418_),
    .B1(_07494_),
    .C1(_07496_),
    .Y(_07498_));
 sky130_fd_sc_hd__o221ai_4 _08369_ (.A1(_07417_),
    .A2(_07418_),
    .B1(_07492_),
    .B2(_07493_),
    .C1(_07496_),
    .Y(_07499_));
 sky130_fd_sc_hd__nand3_1 _08370_ (.A(_07420_),
    .B(_07495_),
    .C(_07494_),
    .Y(_07500_));
 sky130_fd_sc_hd__and3_1 _08371_ (.A(_01499_),
    .B(_05392_),
    .C(_05414_),
    .X(_07501_));
 sky130_fd_sc_hd__nor2_8 _08372_ (.A(net64),
    .B(net34),
    .Y(_07502_));
 sky130_fd_sc_hd__or2_1 _08373_ (.A(net64),
    .B(net34),
    .X(_07503_));
 sky130_fd_sc_hd__nor4_2 _08374_ (.A(net62),
    .B(_07503_),
    .C(net63),
    .D(_04616_),
    .Y(_07504_));
 sky130_fd_sc_hd__nand4b_4 _08375_ (.A_N(_04616_),
    .B(_07502_),
    .C(_00441_),
    .D(_00463_),
    .Y(_07505_));
 sky130_fd_sc_hd__and3_1 _08376_ (.A(_07505_),
    .B(net57),
    .C(_00507_),
    .X(_07506_));
 sky130_fd_sc_hd__a21oi_1 _08377_ (.A1(_07505_),
    .A2(net57),
    .B1(_00507_),
    .Y(_07507_));
 sky130_fd_sc_hd__a21oi_4 _08378_ (.A1(_07505_),
    .A2(net57),
    .B1(net35),
    .Y(_07508_));
 sky130_fd_sc_hd__o21ai_4 _08379_ (.A1(_00299_),
    .A2(net161),
    .B1(_00507_),
    .Y(_07509_));
 sky130_fd_sc_hd__and3_4 _08380_ (.A(_07505_),
    .B(net35),
    .C(net173),
    .X(_07510_));
 sky130_fd_sc_hd__o211ai_4 _08381_ (.A1(net34),
    .A2(_07358_),
    .B1(net35),
    .C1(net57),
    .Y(_07511_));
 sky130_fd_sc_hd__nand2_8 _08382_ (.A(_07509_),
    .B(_07511_),
    .Y(_07512_));
 sky130_fd_sc_hd__nor2_8 _08383_ (.A(_07508_),
    .B(_07510_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand3_4 _08384_ (.A(_07509_),
    .B(_07511_),
    .C(net1),
    .Y(_07514_));
 sky130_fd_sc_hd__o21ai_1 _08385_ (.A1(_00987_),
    .A2(net153),
    .B1(_07514_),
    .Y(_07515_));
 sky130_fd_sc_hd__nand4_2 _08386_ (.A(_00998_),
    .B(_07370_),
    .C(_07513_),
    .D(net1),
    .Y(_07516_));
 sky130_fd_sc_hd__and4_1 _08387_ (.A(net164),
    .B(_06341_),
    .C(_07515_),
    .D(_07516_),
    .X(_07517_));
 sky130_fd_sc_hd__nand4_2 _08388_ (.A(net164),
    .B(_06341_),
    .C(_07515_),
    .D(_07516_),
    .Y(_07518_));
 sky130_fd_sc_hd__a32o_1 _08389_ (.A1(net164),
    .A2(_06309_),
    .A3(_06320_),
    .B1(_07515_),
    .B2(_07516_),
    .X(_07519_));
 sky130_fd_sc_hd__o2111ai_4 _08390_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_05436_),
    .C1(_07518_),
    .D1(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__a32o_1 _08391_ (.A1(_01499_),
    .A2(_05392_),
    .A3(_05414_),
    .B1(_07518_),
    .B2(_07519_),
    .X(_07521_));
 sky130_fd_sc_hd__or4bb_2 _08392_ (.A(_06352_),
    .B(_07371_),
    .C_N(_07520_),
    .D_N(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__a21oi_2 _08393_ (.A1(_07520_),
    .A2(_07521_),
    .B1(_07372_),
    .Y(_07523_));
 sky130_fd_sc_hd__inv_2 _08394_ (.A(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__o2bb2ai_1 _08395_ (.A1_N(_05436_),
    .A2_N(_07375_),
    .B1(_07374_),
    .B2(_06374_),
    .Y(_07525_));
 sky130_fd_sc_hd__o2bb2a_1 _08396_ (.A1_N(_05436_),
    .A2_N(_07375_),
    .B1(_07374_),
    .B2(_06374_),
    .X(_07526_));
 sky130_fd_sc_hd__a21oi_2 _08397_ (.A1(_07522_),
    .A2(_07524_),
    .B1(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__and3_1 _08398_ (.A(_07522_),
    .B(_07524_),
    .C(_07526_),
    .X(_07528_));
 sky130_fd_sc_hd__nor2_1 _08399_ (.A(_07527_),
    .B(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__nand3_2 _08400_ (.A(_07497_),
    .B(_07498_),
    .C(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__o211ai_4 _08401_ (.A1(_07527_),
    .A2(_07528_),
    .B1(_07499_),
    .C1(_07500_),
    .Y(_07531_));
 sky130_fd_sc_hd__inv_2 _08402_ (.A(_07531_),
    .Y(_07532_));
 sky130_fd_sc_hd__o31ai_4 _08403_ (.A1(_07434_),
    .A2(net2),
    .A3(_04190_),
    .B1(net174),
    .Y(_07533_));
 sky130_fd_sc_hd__o311ai_4 _08404_ (.A1(_07434_),
    .A2(net2),
    .A3(_04190_),
    .B1(_00518_),
    .C1(net174),
    .Y(_07534_));
 sky130_fd_sc_hd__nand2_8 _08405_ (.A(_07533_),
    .B(net3),
    .Y(_07535_));
 sky130_fd_sc_hd__nand2_8 _08406_ (.A(_00518_),
    .B(_07533_),
    .Y(_07536_));
 sky130_fd_sc_hd__o31ai_4 _08407_ (.A1(_07434_),
    .A2(net2),
    .A3(_04190_),
    .B1(net3),
    .Y(_07537_));
 sky130_fd_sc_hd__o311ai_4 _08408_ (.A1(_07434_),
    .A2(net2),
    .A3(_04190_),
    .B1(net3),
    .C1(net174),
    .Y(_07538_));
 sky130_fd_sc_hd__o21ai_4 _08409_ (.A1(_00321_),
    .A2(_07537_),
    .B1(_07536_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_8 _08410_ (.A(_07534_),
    .B(_07535_),
    .Y(_07540_));
 sky130_fd_sc_hd__a21o_1 _08411_ (.A1(_07534_),
    .A2(_07535_),
    .B1(_00310_),
    .X(_07541_));
 sky130_fd_sc_hd__a31o_1 _08412_ (.A1(net174),
    .A2(net32),
    .A3(_07103_),
    .B1(_01620_),
    .X(_07542_));
 sky130_fd_sc_hd__o211ai_4 _08413_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_05272_),
    .C1(_05283_),
    .Y(_07543_));
 sky130_fd_sc_hd__and4_1 _08414_ (.A(_05316_),
    .B(_07443_),
    .C(_07157_),
    .D(_01631_),
    .X(_07544_));
 sky130_fd_sc_hd__nand4_1 _08415_ (.A(_05316_),
    .B(_07443_),
    .C(_07157_),
    .D(_01631_),
    .Y(_07545_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(_07444_),
    .B(_07543_),
    .Y(_07546_));
 sky130_fd_sc_hd__nand4_2 _08417_ (.A(_05316_),
    .B(_07444_),
    .C(_01587_),
    .D(_01609_),
    .Y(_07547_));
 sky130_fd_sc_hd__o211ai_2 _08418_ (.A1(_00485_),
    .A2(_07114_),
    .B1(_07443_),
    .C1(_07543_),
    .Y(_07548_));
 sky130_fd_sc_hd__nand4_4 _08419_ (.A(_00911_),
    .B(_07545_),
    .C(_07546_),
    .D(_07440_),
    .Y(_07549_));
 sky130_fd_sc_hd__o211ai_4 _08420_ (.A1(_07441_),
    .A2(_00900_),
    .B1(_07548_),
    .C1(_07547_),
    .Y(_07550_));
 sky130_fd_sc_hd__a32o_1 _08421_ (.A1(net33),
    .A2(_07536_),
    .A3(_07538_),
    .B1(_07549_),
    .B2(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__nand4_1 _08422_ (.A(_07540_),
    .B(_07549_),
    .C(_07550_),
    .D(net33),
    .Y(_07552_));
 sky130_fd_sc_hd__a211o_1 _08423_ (.A1(_07549_),
    .A2(_07550_),
    .B1(_00310_),
    .C1(net150),
    .X(_07553_));
 sky130_fd_sc_hd__nand3_2 _08424_ (.A(_07551_),
    .B(_07552_),
    .C(_07445_),
    .Y(_07554_));
 sky130_fd_sc_hd__a31oi_1 _08425_ (.A1(_07541_),
    .A2(_07549_),
    .A3(_07550_),
    .B1(_07445_),
    .Y(_07555_));
 sky130_fd_sc_hd__nand2_2 _08426_ (.A(_07555_),
    .B(_07553_),
    .Y(_07556_));
 sky130_fd_sc_hd__a2111o_1 _08427_ (.A1(_01303_),
    .A2(_07441_),
    .B1(_05327_),
    .C1(_00310_),
    .D1(_07211_),
    .X(_07557_));
 sky130_fd_sc_hd__nand2_1 _08428_ (.A(_07447_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__a22oi_2 _08429_ (.A1(_07554_),
    .A2(_07556_),
    .B1(_07557_),
    .B2(_07447_),
    .Y(_07559_));
 sky130_fd_sc_hd__and4_1 _08430_ (.A(_07447_),
    .B(_07554_),
    .C(_07556_),
    .D(_07557_),
    .X(_07560_));
 sky130_fd_sc_hd__and3_1 _08431_ (.A(_07558_),
    .B(_07556_),
    .C(_07554_),
    .X(_07561_));
 sky130_fd_sc_hd__a21oi_1 _08432_ (.A1(_07554_),
    .A2(_07556_),
    .B1(_07558_),
    .Y(_07562_));
 sky130_fd_sc_hd__o21a_1 _08433_ (.A1(_07559_),
    .A2(_07560_),
    .B1(_07530_),
    .X(_07563_));
 sky130_fd_sc_hd__o211ai_1 _08434_ (.A1(_07559_),
    .A2(_07560_),
    .B1(_07530_),
    .C1(_07531_),
    .Y(_07564_));
 sky130_fd_sc_hd__o2bb2ai_1 _08435_ (.A1_N(_07530_),
    .A2_N(_07531_),
    .B1(_07561_),
    .B2(_07562_),
    .Y(_07565_));
 sky130_fd_sc_hd__o211ai_2 _08436_ (.A1(_07561_),
    .A2(_07562_),
    .B1(_07530_),
    .C1(_07531_),
    .Y(_07566_));
 sky130_fd_sc_hd__o2bb2ai_1 _08437_ (.A1_N(_07530_),
    .A2_N(_07531_),
    .B1(_07559_),
    .B2(_07560_),
    .Y(_07567_));
 sky130_fd_sc_hd__o2111ai_4 _08438_ (.A1(_07454_),
    .A2(_07430_),
    .B1(_07432_),
    .C1(_07566_),
    .D1(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__nand3_2 _08439_ (.A(_07565_),
    .B(_07465_),
    .C(_07564_),
    .Y(_07569_));
 sky130_fd_sc_hd__a31oi_1 _08440_ (.A1(_07457_),
    .A2(_07458_),
    .A3(_07348_),
    .B1(_07286_),
    .Y(_07570_));
 sky130_fd_sc_hd__a31o_1 _08441_ (.A1(_07457_),
    .A2(_07458_),
    .A3(_07348_),
    .B1(_07286_),
    .X(_07571_));
 sky130_fd_sc_hd__o2111a_1 _08442_ (.A1(_07459_),
    .A2(_07348_),
    .B1(_07569_),
    .C1(_07568_),
    .D1(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__o2bb2ai_1 _08443_ (.A1_N(_07568_),
    .A2_N(_07569_),
    .B1(_07570_),
    .B2(_07460_),
    .Y(_07573_));
 sky130_fd_sc_hd__nand2b_1 _08444_ (.A_N(_07572_),
    .B(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__xnor2_1 _08445_ (.A(_07464_),
    .B(_07574_),
    .Y(net67));
 sky130_fd_sc_hd__o211ai_2 _08446_ (.A1(_07459_),
    .A2(_07348_),
    .B1(_07571_),
    .C1(_07569_),
    .Y(_07575_));
 sky130_fd_sc_hd__o21ai_1 _08447_ (.A1(_07460_),
    .A2(_07570_),
    .B1(_07568_),
    .Y(_07576_));
 sky130_fd_sc_hd__o21ai_1 _08448_ (.A1(_07561_),
    .A2(_07562_),
    .B1(_07531_),
    .Y(_07577_));
 sky130_fd_sc_hd__nand2_1 _08449_ (.A(_07530_),
    .B(_07577_),
    .Y(_07578_));
 sky130_fd_sc_hd__o31a_1 _08450_ (.A1(_07532_),
    .A2(_07559_),
    .A3(_07560_),
    .B1(_07530_),
    .X(_07579_));
 sky130_fd_sc_hd__a31oi_1 _08451_ (.A1(_07520_),
    .A2(_07521_),
    .A3(_07372_),
    .B1(_07525_),
    .Y(_07580_));
 sky130_fd_sc_hd__o21ai_2 _08452_ (.A1(_07526_),
    .A2(_07523_),
    .B1(_07522_),
    .Y(_07581_));
 sky130_fd_sc_hd__a21oi_1 _08453_ (.A1(_07519_),
    .A2(_07501_),
    .B1(_07517_),
    .Y(_07582_));
 sky130_fd_sc_hd__o21ai_1 _08454_ (.A1(_01892_),
    .A2(_01914_),
    .B1(_05414_),
    .Y(_07583_));
 sky130_fd_sc_hd__and3_1 _08455_ (.A(_01969_),
    .B(_05392_),
    .C(_05414_),
    .X(_07584_));
 sky130_fd_sc_hd__and3_1 _08456_ (.A(_01499_),
    .B(_06309_),
    .C(_06320_),
    .X(_00000_));
 sky130_fd_sc_hd__o211a_1 _08457_ (.A1(_00299_),
    .A2(_07366_),
    .B1(_07368_),
    .C1(net164),
    .X(_00001_));
 sky130_fd_sc_hd__nand4_4 _08458_ (.A(_05348_),
    .B(_07502_),
    .C(_00463_),
    .D(_00507_),
    .Y(_00002_));
 sky130_fd_sc_hd__o211a_4 _08459_ (.A1(net35),
    .A2(_07505_),
    .B1(_00529_),
    .C1(net57),
    .X(_00003_));
 sky130_fd_sc_hd__a21oi_4 _08460_ (.A1(_00002_),
    .A2(net57),
    .B1(_00529_),
    .Y(_00004_));
 sky130_fd_sc_hd__a21oi_4 _08461_ (.A1(_00002_),
    .A2(net57),
    .B1(net36),
    .Y(_00005_));
 sky130_fd_sc_hd__a21o_4 _08462_ (.A1(_00002_),
    .A2(net57),
    .B1(net36),
    .X(_00006_));
 sky130_fd_sc_hd__o211a_4 _08463_ (.A1(net35),
    .A2(_07505_),
    .B1(net36),
    .C1(net57),
    .X(_00007_));
 sky130_fd_sc_hd__a311o_4 _08464_ (.A1(_06254_),
    .A2(_07502_),
    .A3(_00507_),
    .B1(_00529_),
    .C1(_00299_),
    .X(_00008_));
 sky130_fd_sc_hd__nand2_8 _08465_ (.A(_00006_),
    .B(_00008_),
    .Y(_00009_));
 sky130_fd_sc_hd__nor2_8 _08466_ (.A(_00005_),
    .B(_00007_),
    .Y(_00010_));
 sky130_fd_sc_hd__o21ai_4 _08467_ (.A1(_00003_),
    .A2(_00004_),
    .B1(_00998_),
    .Y(_00011_));
 sky130_fd_sc_hd__a31oi_1 _08468_ (.A1(_00002_),
    .A2(net36),
    .A3(net57),
    .B1(_00288_),
    .Y(_00012_));
 sky130_fd_sc_hd__a31o_1 _08469_ (.A1(_00002_),
    .A2(net36),
    .A3(net57),
    .B1(_00288_),
    .X(_00013_));
 sky130_fd_sc_hd__nand4_2 _08470_ (.A(_07513_),
    .B(_00012_),
    .C(_00006_),
    .D(_00998_),
    .Y(_00014_));
 sky130_fd_sc_hd__o32ai_4 _08471_ (.A1(_00987_),
    .A2(_07508_),
    .A3(_07510_),
    .B1(_00005_),
    .B2(_00013_),
    .Y(_00015_));
 sky130_fd_sc_hd__o311a_1 _08472_ (.A1(_00987_),
    .A2(_07514_),
    .A3(_00009_),
    .B1(_00015_),
    .C1(_00001_),
    .X(_00016_));
 sky130_fd_sc_hd__o2111ai_2 _08473_ (.A1(_07514_),
    .A2(_00011_),
    .B1(_00015_),
    .C1(_07370_),
    .D1(net164),
    .Y(_00017_));
 sky130_fd_sc_hd__a21oi_2 _08474_ (.A1(_00014_),
    .A2(_00015_),
    .B1(_00001_),
    .Y(_00018_));
 sky130_fd_sc_hd__nand3b_1 _08475_ (.A_N(_00018_),
    .B(_00000_),
    .C(_00017_),
    .Y(_00019_));
 sky130_fd_sc_hd__o22ai_2 _08476_ (.A1(_01488_),
    .A2(_06331_),
    .B1(_00016_),
    .B2(_00018_),
    .Y(_00020_));
 sky130_fd_sc_hd__nand3b_2 _08477_ (.A_N(_07516_),
    .B(_00019_),
    .C(_00020_),
    .Y(_00021_));
 sky130_fd_sc_hd__o2bb2ai_2 _08478_ (.A1_N(_00019_),
    .A2_N(_00020_),
    .B1(_07371_),
    .B2(_07514_),
    .Y(_00022_));
 sky130_fd_sc_hd__o2bb2ai_2 _08479_ (.A1_N(_00021_),
    .A2_N(_00022_),
    .B1(_05381_),
    .B2(_07583_),
    .Y(_00023_));
 sky130_fd_sc_hd__nand4_1 _08480_ (.A(_01969_),
    .B(_05436_),
    .C(_00021_),
    .D(_00022_),
    .Y(_00024_));
 sky130_fd_sc_hd__a31oi_2 _08481_ (.A1(_00022_),
    .A2(_07584_),
    .A3(_00021_),
    .B1(_07582_),
    .Y(_00025_));
 sky130_fd_sc_hd__a21boi_2 _08482_ (.A1(_00023_),
    .A2(_00024_),
    .B1_N(_07582_),
    .Y(_00026_));
 sky130_fd_sc_hd__a21oi_2 _08483_ (.A1(_00023_),
    .A2(_00025_),
    .B1(_00026_),
    .Y(_00027_));
 sky130_fd_sc_hd__xor2_4 _08484_ (.A(_07581_),
    .B(_00027_),
    .X(_00028_));
 sky130_fd_sc_hd__inv_2 _08485_ (.A(_00028_),
    .Y(_00029_));
 sky130_fd_sc_hd__a31o_2 _08486_ (.A1(_02866_),
    .A2(_03917_),
    .A3(_07474_),
    .B1(_07472_),
    .X(_00030_));
 sky130_fd_sc_hd__a32oi_2 _08487_ (.A1(_07394_),
    .A2(_07469_),
    .A3(_07397_),
    .B1(_07479_),
    .B2(_07471_),
    .Y(_00031_));
 sky130_fd_sc_hd__or3_1 _08488_ (.A(net167),
    .B(_02833_),
    .C(_04244_),
    .X(_00032_));
 sky130_fd_sc_hd__o32a_1 _08489_ (.A1(_03479_),
    .A2(_03522_),
    .A3(_03906_),
    .B1(_04715_),
    .B2(_02636_),
    .X(_00033_));
 sky130_fd_sc_hd__and3_1 _08490_ (.A(_02647_),
    .B(_03917_),
    .C(_04726_),
    .X(_00034_));
 sky130_fd_sc_hd__a21oi_1 _08491_ (.A1(_00034_),
    .A2(net157),
    .B1(_00033_),
    .Y(_00035_));
 sky130_fd_sc_hd__xnor2_1 _08492_ (.A(_00032_),
    .B(_00035_),
    .Y(_00036_));
 sky130_fd_sc_hd__and2_1 _08493_ (.A(_00031_),
    .B(_00036_),
    .X(_00037_));
 sky130_fd_sc_hd__nor2_1 _08494_ (.A(_00031_),
    .B(_00036_),
    .Y(_00038_));
 sky130_fd_sc_hd__nor2_1 _08495_ (.A(_00037_),
    .B(_00038_),
    .Y(_00039_));
 sky130_fd_sc_hd__o21bai_4 _08496_ (.A1(_00030_),
    .A2(_00037_),
    .B1_N(_00038_),
    .Y(_00040_));
 sky130_fd_sc_hd__o21ba_2 _08497_ (.A1(_00030_),
    .A2(_00037_),
    .B1_N(_00038_),
    .X(_00041_));
 sky130_fd_sc_hd__xnor2_4 _08498_ (.A(_00030_),
    .B(_00039_),
    .Y(_00042_));
 sky130_fd_sc_hd__and3_2 _08499_ (.A(_02133_),
    .B(_04255_),
    .C(_07487_),
    .X(_00043_));
 sky130_fd_sc_hd__nor2_1 _08500_ (.A(_07485_),
    .B(_00043_),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_1 _08501_ (.A(_00044_),
    .B(_00042_),
    .Y(_00045_));
 sky130_fd_sc_hd__inv_2 _08502_ (.A(_00045_),
    .Y(_00046_));
 sky130_fd_sc_hd__o21ai_4 _08503_ (.A1(_07482_),
    .A2(_07484_),
    .B1(_00042_),
    .Y(_00047_));
 sky130_fd_sc_hd__nand2_1 _08504_ (.A(_00042_),
    .B(_00044_),
    .Y(_00048_));
 sky130_fd_sc_hd__and2b_1 _08505_ (.A_N(_00045_),
    .B(_00048_),
    .X(_00049_));
 sky130_fd_sc_hd__o21bai_2 _08506_ (.A1(_00043_),
    .A2(_00047_),
    .B1_N(_00045_),
    .Y(_00050_));
 sky130_fd_sc_hd__o211ai_4 _08507_ (.A1(_07490_),
    .A2(_07466_),
    .B1(_07421_),
    .C1(_07496_),
    .Y(_00051_));
 sky130_fd_sc_hd__o211ai_4 _08508_ (.A1(_07491_),
    .A2(_07467_),
    .B1(_07420_),
    .C1(_07495_),
    .Y(_00052_));
 sky130_fd_sc_hd__o211ai_1 _08509_ (.A1(_07467_),
    .A2(_07491_),
    .B1(_00050_),
    .C1(_00051_),
    .Y(_00053_));
 sky130_fd_sc_hd__o211ai_1 _08510_ (.A1(_07466_),
    .A2(_07490_),
    .B1(_00049_),
    .C1(_00052_),
    .Y(_00054_));
 sky130_fd_sc_hd__o211ai_4 _08511_ (.A1(_07466_),
    .A2(_07490_),
    .B1(_00050_),
    .C1(_00052_),
    .Y(_00055_));
 sky130_fd_sc_hd__o211ai_4 _08512_ (.A1(_07467_),
    .A2(_07491_),
    .B1(_00049_),
    .C1(_00051_),
    .Y(_00056_));
 sky130_fd_sc_hd__nand3_2 _08513_ (.A(_00055_),
    .B(_00056_),
    .C(_00028_),
    .Y(_00057_));
 sky130_fd_sc_hd__a21oi_4 _08514_ (.A1(_00055_),
    .A2(_00056_),
    .B1(_00028_),
    .Y(_00058_));
 sky130_fd_sc_hd__nand3_1 _08515_ (.A(_00029_),
    .B(_00053_),
    .C(_00054_),
    .Y(_00059_));
 sky130_fd_sc_hd__a21bo_1 _08516_ (.A1(_07556_),
    .A2(_07558_),
    .B1_N(_07554_),
    .X(_00060_));
 sky130_fd_sc_hd__a21boi_1 _08517_ (.A1(_07558_),
    .A2(_07556_),
    .B1_N(_07554_),
    .Y(_00061_));
 sky130_fd_sc_hd__nor2_4 _08518_ (.A(net2),
    .B(net3),
    .Y(_00062_));
 sky130_fd_sc_hd__nor4_4 _08519_ (.A(net2),
    .B(_07434_),
    .C(net3),
    .D(_04190_),
    .Y(_00063_));
 sky130_fd_sc_hd__nand3b_2 _08520_ (.A_N(_04190_),
    .B(_07433_),
    .C(_00062_),
    .Y(_00064_));
 sky130_fd_sc_hd__o41ai_1 _08521_ (.A1(net2),
    .A2(_07434_),
    .A3(net3),
    .A4(_04190_),
    .B1(net174),
    .Y(_00065_));
 sky130_fd_sc_hd__nand2_8 _08522_ (.A(net174),
    .B(net4),
    .Y(_00066_));
 sky130_fd_sc_hd__a21oi_4 _08523_ (.A1(_07435_),
    .A2(_00062_),
    .B1(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__a31o_1 _08524_ (.A1(_07435_),
    .A2(_00518_),
    .A3(_00496_),
    .B1(_00066_),
    .X(_00068_));
 sky130_fd_sc_hd__a21oi_4 _08525_ (.A1(_00064_),
    .A2(net174),
    .B1(net4),
    .Y(_00069_));
 sky130_fd_sc_hd__o21ai_4 _08526_ (.A1(_00321_),
    .A2(net160),
    .B1(_00540_),
    .Y(_00070_));
 sky130_fd_sc_hd__o21ai_4 _08527_ (.A1(net160),
    .A2(_00066_),
    .B1(_00070_),
    .Y(_00071_));
 sky130_fd_sc_hd__o21a_4 _08528_ (.A1(net160),
    .A2(_00066_),
    .B1(_00070_),
    .X(_00072_));
 sky130_fd_sc_hd__or3_1 _08529_ (.A(_00310_),
    .B(_00067_),
    .C(_00069_),
    .X(_00073_));
 sky130_fd_sc_hd__o221ai_4 _08530_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_07537_),
    .B2(_00321_),
    .C1(_07536_),
    .Y(_00074_));
 sky130_fd_sc_hd__o211ai_2 _08531_ (.A1(net170),
    .A2(_02057_),
    .B1(_05272_),
    .C1(_05283_),
    .Y(_00075_));
 sky130_fd_sc_hd__o21ai_4 _08532_ (.A1(_07168_),
    .A2(_07542_),
    .B1(_00075_),
    .Y(_00076_));
 sky130_fd_sc_hd__a22oi_4 _08533_ (.A1(_02046_),
    .A2(_02068_),
    .B1(_07114_),
    .B2(_00485_),
    .Y(_00077_));
 sky130_fd_sc_hd__o211ai_4 _08534_ (.A1(net170),
    .A2(_02057_),
    .B1(_07157_),
    .C1(_07178_),
    .Y(_00078_));
 sky130_fd_sc_hd__o2111ai_4 _08535_ (.A1(_00485_),
    .A2(_07114_),
    .B1(_00077_),
    .C1(_01631_),
    .D1(_05316_),
    .Y(_00079_));
 sky130_fd_sc_hd__a22oi_4 _08536_ (.A1(_07440_),
    .A2(_01303_),
    .B1(_00079_),
    .B2(_00076_),
    .Y(_00080_));
 sky130_fd_sc_hd__a32o_1 _08537_ (.A1(_01270_),
    .A2(_07440_),
    .A3(_01281_),
    .B1(_00079_),
    .B2(_00076_),
    .X(_00081_));
 sky130_fd_sc_hd__o2111a_1 _08538_ (.A1(_07543_),
    .A2(_00078_),
    .B1(_07440_),
    .C1(_00076_),
    .D1(_01303_),
    .X(_00082_));
 sky130_fd_sc_hd__o2111ai_2 _08539_ (.A1(_07543_),
    .A2(_00078_),
    .B1(_07440_),
    .C1(_00076_),
    .D1(_01303_),
    .Y(_00083_));
 sky130_fd_sc_hd__o22ai_4 _08540_ (.A1(_00900_),
    .A2(net150),
    .B1(_00080_),
    .B2(_00082_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand3b_2 _08541_ (.A_N(_00074_),
    .B(_00081_),
    .C(_00083_),
    .Y(_00085_));
 sky130_fd_sc_hd__nand3_2 _08542_ (.A(_00085_),
    .B(_07544_),
    .C(_00084_),
    .Y(_00086_));
 sky130_fd_sc_hd__a21oi_1 _08543_ (.A1(_00084_),
    .A2(_00085_),
    .B1(_07544_),
    .Y(_00087_));
 sky130_fd_sc_hd__o2bb2ai_2 _08544_ (.A1_N(_00084_),
    .A2_N(_00085_),
    .B1(_07444_),
    .B2(_07543_),
    .Y(_00088_));
 sky130_fd_sc_hd__a22o_1 _08545_ (.A1(_00072_),
    .A2(net33),
    .B1(_00088_),
    .B2(_00086_),
    .X(_00089_));
 sky130_fd_sc_hd__nand4_4 _08546_ (.A(_00072_),
    .B(_00086_),
    .C(_00088_),
    .D(net33),
    .Y(_00090_));
 sky130_fd_sc_hd__and2_1 _08547_ (.A(_00089_),
    .B(_00090_),
    .X(_00091_));
 sky130_fd_sc_hd__a21boi_4 _08548_ (.A1(_07541_),
    .A2(_07549_),
    .B1_N(_07550_),
    .Y(_00092_));
 sky130_fd_sc_hd__a21oi_2 _08549_ (.A1(_00089_),
    .A2(_00090_),
    .B1(_00092_),
    .Y(_00093_));
 sky130_fd_sc_hd__and3_1 _08550_ (.A(_00089_),
    .B(_00090_),
    .C(_00092_),
    .X(_00094_));
 sky130_fd_sc_hd__or2_1 _08551_ (.A(_00093_),
    .B(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__and2_1 _08552_ (.A(_00061_),
    .B(_00095_),
    .X(_00096_));
 sky130_fd_sc_hd__nor2_1 _08553_ (.A(_00061_),
    .B(_00095_),
    .Y(_00097_));
 sky130_fd_sc_hd__a31oi_4 _08554_ (.A1(_00089_),
    .A2(_00090_),
    .A3(_00092_),
    .B1(_00060_),
    .Y(_00098_));
 sky130_fd_sc_hd__o21a_1 _08555_ (.A1(_00091_),
    .A2(_00092_),
    .B1(_00098_),
    .X(_00099_));
 sky130_fd_sc_hd__and2_1 _08556_ (.A(_00095_),
    .B(_00060_),
    .X(_00100_));
 sky130_fd_sc_hd__nor2_1 _08557_ (.A(_00099_),
    .B(_00100_),
    .Y(_00101_));
 sky130_fd_sc_hd__o211ai_1 _08558_ (.A1(_00096_),
    .A2(_00097_),
    .B1(_00057_),
    .C1(_00059_),
    .Y(_00102_));
 sky130_fd_sc_hd__o2bb2ai_1 _08559_ (.A1_N(_00057_),
    .A2_N(_00059_),
    .B1(_00099_),
    .B2(_00100_),
    .Y(_00103_));
 sky130_fd_sc_hd__o2bb2ai_2 _08560_ (.A1_N(_00057_),
    .A2_N(_00059_),
    .B1(_00096_),
    .B2(_00097_),
    .Y(_00104_));
 sky130_fd_sc_hd__a31o_1 _08561_ (.A1(_00055_),
    .A2(_00056_),
    .A3(_00028_),
    .B1(_00101_),
    .X(_00105_));
 sky130_fd_sc_hd__o21ai_1 _08562_ (.A1(_00058_),
    .A2(_00105_),
    .B1(_00104_),
    .Y(_00106_));
 sky130_fd_sc_hd__o21a_1 _08563_ (.A1(_00058_),
    .A2(_00105_),
    .B1(_00104_),
    .X(_00107_));
 sky130_fd_sc_hd__nand3_1 _08564_ (.A(_00103_),
    .B(_07578_),
    .C(_00102_),
    .Y(_00108_));
 sky130_fd_sc_hd__o221ai_4 _08565_ (.A1(_07532_),
    .A2(_07563_),
    .B1(_00058_),
    .B2(_00105_),
    .C1(_00104_),
    .Y(_00109_));
 sky130_fd_sc_hd__a22oi_1 _08566_ (.A1(_07568_),
    .A2(_07575_),
    .B1(_00108_),
    .B2(_00109_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand3_1 _08567_ (.A(_07569_),
    .B(_07576_),
    .C(_00109_),
    .Y(_00111_));
 sky130_fd_sc_hd__nand3_1 _08568_ (.A(_07568_),
    .B(_07575_),
    .C(_00108_),
    .Y(_00112_));
 sky130_fd_sc_hd__a41o_1 _08569_ (.A1(_07568_),
    .A2(_07575_),
    .A3(_00108_),
    .A4(_00109_),
    .B1(_00110_),
    .X(_00113_));
 sky130_fd_sc_hd__nor4_2 _08570_ (.A(_06232_),
    .B(_07296_),
    .C(_07574_),
    .D(_07463_),
    .Y(_00114_));
 sky130_fd_sc_hd__or3_1 _08571_ (.A(_00834_),
    .B(_00113_),
    .C(_00114_),
    .X(_00115_));
 sky130_fd_sc_hd__o21ai_1 _08572_ (.A1(_00834_),
    .A2(_00114_),
    .B1(_00113_),
    .Y(_00116_));
 sky130_fd_sc_hd__and2_1 _08573_ (.A(_00115_),
    .B(_00116_),
    .X(net68));
 sky130_fd_sc_hd__o2bb2a_1 _08574_ (.A1_N(_00113_),
    .A2_N(_00114_),
    .B1(_00812_),
    .B2(_00823_),
    .X(_00117_));
 sky130_fd_sc_hd__a221o_4 _08575_ (.A1(net173),
    .A2(_03501_),
    .B1(_04201_),
    .B2(_04212_),
    .C1(_03479_),
    .X(_00118_));
 sky130_fd_sc_hd__a2bb2o_1 _08576_ (.A1_N(_00033_),
    .A2_N(_00032_),
    .B1(net157),
    .B2(_02647_),
    .X(_00119_));
 sky130_fd_sc_hd__or4b_1 _08577_ (.A(_03906_),
    .B(_04671_),
    .C(_04693_),
    .D_N(_00119_),
    .X(_00120_));
 sky130_fd_sc_hd__o32a_1 _08578_ (.A1(net159),
    .A2(_04244_),
    .A3(_00033_),
    .B1(_04715_),
    .B2(_03906_),
    .X(_00121_));
 sky130_fd_sc_hd__a31o_2 _08579_ (.A1(_03917_),
    .A2(_04726_),
    .A3(_00119_),
    .B1(_00121_),
    .X(_00122_));
 sky130_fd_sc_hd__xor2_4 _08580_ (.A(_00118_),
    .B(_00122_),
    .X(_00123_));
 sky130_fd_sc_hd__xnor2_2 _08581_ (.A(_00118_),
    .B(_00122_),
    .Y(_00124_));
 sky130_fd_sc_hd__xor2_2 _08582_ (.A(_00040_),
    .B(_00123_),
    .X(_00125_));
 sky130_fd_sc_hd__inv_2 _08583_ (.A(_00125_),
    .Y(_00126_));
 sky130_fd_sc_hd__o211ai_4 _08584_ (.A1(_07466_),
    .A2(_07490_),
    .B1(_00046_),
    .C1(_00052_),
    .Y(_00127_));
 sky130_fd_sc_hd__o211ai_2 _08585_ (.A1(_07467_),
    .A2(_07491_),
    .B1(_00048_),
    .C1(_00051_),
    .Y(_00128_));
 sky130_fd_sc_hd__o211ai_2 _08586_ (.A1(_00043_),
    .A2(_00047_),
    .B1(_00126_),
    .C1(_00127_),
    .Y(_00129_));
 sky130_fd_sc_hd__o211ai_2 _08587_ (.A1(_00042_),
    .A2(_00044_),
    .B1(_00125_),
    .C1(_00128_),
    .Y(_00130_));
 sky130_fd_sc_hd__o211ai_1 _08588_ (.A1(_00043_),
    .A2(_00047_),
    .B1(_00125_),
    .C1(_00127_),
    .Y(_00131_));
 sky130_fd_sc_hd__o211ai_1 _08589_ (.A1(_00042_),
    .A2(_00044_),
    .B1(_00126_),
    .C1(_00128_),
    .Y(_00132_));
 sky130_fd_sc_hd__and3_2 _08590_ (.A(_02647_),
    .B(_05392_),
    .C(_05414_),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _08591_ (.A1(_01903_),
    .A2(_01925_),
    .B1(_06276_),
    .B2(_06298_),
    .X(_00134_));
 sky130_fd_sc_hd__and3_1 _08592_ (.A(_00000_),
    .B(_07370_),
    .C(_01969_),
    .X(_00135_));
 sky130_fd_sc_hd__o22a_1 _08593_ (.A1(_01958_),
    .A2(_06331_),
    .B1(net153),
    .B2(_01488_),
    .X(_00136_));
 sky130_fd_sc_hd__a31oi_1 _08594_ (.A1(_01969_),
    .A2(_07370_),
    .A3(_00000_),
    .B1(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__a31o_1 _08595_ (.A1(_01969_),
    .A2(_07370_),
    .A3(_00000_),
    .B1(_00136_),
    .X(_00138_));
 sky130_fd_sc_hd__o221a_1 _08596_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_07506_),
    .B2(_07507_),
    .C1(_01172_),
    .X(_00139_));
 sky130_fd_sc_hd__nor2_8 _08597_ (.A(net35),
    .B(net36),
    .Y(_00140_));
 sky130_fd_sc_hd__or2_1 _08598_ (.A(net35),
    .B(net36),
    .X(_00141_));
 sky130_fd_sc_hd__and3_4 _08599_ (.A(_06254_),
    .B(_07502_),
    .C(_00140_),
    .X(_00142_));
 sky130_fd_sc_hd__nand4_4 _08600_ (.A(_05348_),
    .B(_07502_),
    .C(_00140_),
    .D(_00463_),
    .Y(_00143_));
 sky130_fd_sc_hd__nand2_8 _08601_ (.A(net57),
    .B(net37),
    .Y(_00144_));
 sky130_fd_sc_hd__a21oi_4 _08602_ (.A1(net161),
    .A2(_00140_),
    .B1(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__a31o_4 _08603_ (.A1(net161),
    .A2(_00529_),
    .A3(_00507_),
    .B1(_00144_),
    .X(_00146_));
 sky130_fd_sc_hd__a21oi_4 _08604_ (.A1(_00143_),
    .A2(net57),
    .B1(net37),
    .Y(_00147_));
 sky130_fd_sc_hd__a21o_4 _08605_ (.A1(_00143_),
    .A2(net57),
    .B1(net37),
    .X(_00148_));
 sky130_fd_sc_hd__o21ai_4 _08606_ (.A1(_00142_),
    .A2(_00144_),
    .B1(_00148_),
    .Y(_00149_));
 sky130_fd_sc_hd__nor2_8 _08607_ (.A(_00145_),
    .B(_00147_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand3_1 _08608_ (.A(_00148_),
    .B(net1),
    .C(_00146_),
    .Y(_00151_));
 sky130_fd_sc_hd__o31ai_4 _08609_ (.A1(_00987_),
    .A2(_00005_),
    .A3(_00007_),
    .B1(_00151_),
    .Y(_00152_));
 sky130_fd_sc_hd__a31oi_2 _08610_ (.A1(_00143_),
    .A2(net37),
    .A3(net57),
    .B1(_00987_),
    .Y(_00153_));
 sky130_fd_sc_hd__o2111ai_4 _08611_ (.A1(net172),
    .A2(_00943_),
    .B1(net1),
    .C1(_00146_),
    .D1(_00148_),
    .Y(_00154_));
 sky130_fd_sc_hd__o21ai_1 _08612_ (.A1(_00009_),
    .A2(_00154_),
    .B1(_00152_),
    .Y(_00155_));
 sky130_fd_sc_hd__nand2_1 _08613_ (.A(_00155_),
    .B(_00139_),
    .Y(_00156_));
 sky130_fd_sc_hd__o221ai_4 _08614_ (.A1(net165),
    .A2(_07512_),
    .B1(_00009_),
    .B2(_00154_),
    .C1(_00152_),
    .Y(_00157_));
 sky130_fd_sc_hd__o21ai_1 _08615_ (.A1(net165),
    .A2(_07512_),
    .B1(_00155_),
    .Y(_00158_));
 sky130_fd_sc_hd__o2111ai_2 _08616_ (.A1(_00154_),
    .A2(_00009_),
    .B1(_07513_),
    .C1(net164),
    .D1(_00152_),
    .Y(_00159_));
 sky130_fd_sc_hd__o211a_1 _08617_ (.A1(_00135_),
    .A2(_00136_),
    .B1(_00156_),
    .C1(_00157_),
    .X(_00160_));
 sky130_fd_sc_hd__nand3_2 _08618_ (.A(_00138_),
    .B(_00156_),
    .C(_00157_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand3_2 _08619_ (.A(_00158_),
    .B(_00159_),
    .C(_00137_),
    .Y(_00162_));
 sky130_fd_sc_hd__o2bb2ai_1 _08620_ (.A1_N(_00161_),
    .A2_N(_00162_),
    .B1(_07514_),
    .B2(_00011_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand3b_1 _08621_ (.A_N(_00014_),
    .B(_00161_),
    .C(_00162_),
    .Y(_00164_));
 sky130_fd_sc_hd__o21ai_4 _08622_ (.A1(_07514_),
    .A2(_00011_),
    .B1(_00162_),
    .Y(_00165_));
 sky130_fd_sc_hd__a21o_1 _08623_ (.A1(_00161_),
    .A2(_00162_),
    .B1(_00014_),
    .X(_00166_));
 sky130_fd_sc_hd__o31ai_2 _08624_ (.A1(_01488_),
    .A2(_06331_),
    .A3(_00018_),
    .B1(_00017_),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _08625_ (.A(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__o211ai_4 _08626_ (.A1(_00165_),
    .A2(_00160_),
    .B1(_00168_),
    .C1(_00166_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand3_2 _08627_ (.A(_00163_),
    .B(_00164_),
    .C(_00167_),
    .Y(_00170_));
 sky130_fd_sc_hd__a21oi_1 _08628_ (.A1(_00169_),
    .A2(_00170_),
    .B1(_00133_),
    .Y(_00171_));
 sky130_fd_sc_hd__a32o_1 _08629_ (.A1(_02647_),
    .A2(_05392_),
    .A3(_05414_),
    .B1(_00169_),
    .B2(_00170_),
    .X(_00172_));
 sky130_fd_sc_hd__and3_1 _08630_ (.A(_00169_),
    .B(_00170_),
    .C(_00133_),
    .X(_00173_));
 sky130_fd_sc_hd__a21boi_1 _08631_ (.A1(_00022_),
    .A2(_07584_),
    .B1_N(_00021_),
    .Y(_00174_));
 sky130_fd_sc_hd__o21ai_2 _08632_ (.A1(_00171_),
    .A2(_00173_),
    .B1(_00174_),
    .Y(_00175_));
 sky130_fd_sc_hd__a31oi_1 _08633_ (.A1(_00169_),
    .A2(_00170_),
    .A3(_00133_),
    .B1(_00174_),
    .Y(_00176_));
 sky130_fd_sc_hd__a31o_1 _08634_ (.A1(_00169_),
    .A2(_00170_),
    .A3(_00133_),
    .B1(_00174_),
    .X(_00177_));
 sky130_fd_sc_hd__o21ai_1 _08635_ (.A1(_00171_),
    .A2(_00177_),
    .B1(_00175_),
    .Y(_00178_));
 sky130_fd_sc_hd__a2bb2oi_1 _08636_ (.A1_N(_07523_),
    .A2_N(_07580_),
    .B1(_00023_),
    .B2(_00025_),
    .Y(_00179_));
 sky130_fd_sc_hd__nor2_1 _08637_ (.A(_00026_),
    .B(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__xor2_2 _08638_ (.A(_00178_),
    .B(_00180_),
    .X(_00181_));
 sky130_fd_sc_hd__inv_2 _08639_ (.A(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand3_2 _08640_ (.A(_00129_),
    .B(_00130_),
    .C(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand3_2 _08641_ (.A(_00131_),
    .B(_00132_),
    .C(_00181_),
    .Y(_00184_));
 sky130_fd_sc_hd__nand4b_4 _08642_ (.A_N(_04190_),
    .B(_07433_),
    .C(_00062_),
    .D(_00540_),
    .Y(_00185_));
 sky130_fd_sc_hd__and3_1 _08643_ (.A(_00185_),
    .B(net25),
    .C(_00561_),
    .X(_00186_));
 sky130_fd_sc_hd__a21oi_1 _08644_ (.A1(_00185_),
    .A2(net25),
    .B1(_00561_),
    .Y(_00187_));
 sky130_fd_sc_hd__and3_4 _08645_ (.A(_00185_),
    .B(net5),
    .C(net174),
    .X(_00188_));
 sky130_fd_sc_hd__o211ai_4 _08646_ (.A1(net4),
    .A2(_00064_),
    .B1(net5),
    .C1(net174),
    .Y(_00189_));
 sky130_fd_sc_hd__a21oi_4 _08647_ (.A1(_00185_),
    .A2(net174),
    .B1(net5),
    .Y(_00190_));
 sky130_fd_sc_hd__a21o_4 _08648_ (.A1(_00185_),
    .A2(net174),
    .B1(net5),
    .X(_00191_));
 sky130_fd_sc_hd__nand2_8 _08649_ (.A(_00189_),
    .B(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__nor2_8 _08650_ (.A(_00188_),
    .B(_00190_),
    .Y(_00193_));
 sky130_fd_sc_hd__o21a_1 _08651_ (.A1(_00900_),
    .A2(net150),
    .B1(_00083_),
    .X(_00194_));
 sky130_fd_sc_hd__a31o_1 _08652_ (.A1(_00911_),
    .A2(_07540_),
    .A3(_00081_),
    .B1(_00082_),
    .X(_00195_));
 sky130_fd_sc_hd__o221ai_4 _08653_ (.A1(_01238_),
    .A2(_01249_),
    .B1(_00063_),
    .B2(_00066_),
    .C1(_00070_),
    .Y(_00196_));
 sky130_fd_sc_hd__nor2_2 _08654_ (.A(_00074_),
    .B(_00196_),
    .Y(_00197_));
 sky130_fd_sc_hd__or3_1 _08655_ (.A(_00900_),
    .B(_00067_),
    .C(_00069_),
    .X(_00198_));
 sky130_fd_sc_hd__o32a_1 _08656_ (.A1(_00900_),
    .A2(_00067_),
    .A3(_00069_),
    .B1(_01292_),
    .B2(net150),
    .X(_00199_));
 sky130_fd_sc_hd__a32o_1 _08657_ (.A1(_00911_),
    .A2(_00068_),
    .A3(_00070_),
    .B1(_01303_),
    .B2(_07540_),
    .X(_00200_));
 sky130_fd_sc_hd__o211ai_4 _08658_ (.A1(net169),
    .A2(net163),
    .B1(_05272_),
    .C1(_05283_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_2 _08659_ (.A(_00078_),
    .B(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__and4_1 _08660_ (.A(_05316_),
    .B(_07157_),
    .C(_00077_),
    .D(_02866_),
    .X(_00203_));
 sky130_fd_sc_hd__nand4_2 _08661_ (.A(_05316_),
    .B(_07157_),
    .C(_00077_),
    .D(_02866_),
    .Y(_00204_));
 sky130_fd_sc_hd__and3_1 _08662_ (.A(_01631_),
    .B(net162),
    .C(net154),
    .X(_00205_));
 sky130_fd_sc_hd__a22o_1 _08663_ (.A1(_01543_),
    .A2(_01565_),
    .B1(_07438_),
    .B2(_07439_),
    .X(_00206_));
 sky130_fd_sc_hd__nand4_1 _08664_ (.A(_01631_),
    .B(_00202_),
    .C(_00204_),
    .D(_07440_),
    .Y(_00207_));
 sky130_fd_sc_hd__o2bb2ai_1 _08665_ (.A1_N(_00202_),
    .A2_N(_00204_),
    .B1(_01620_),
    .B2(_07441_),
    .Y(_00208_));
 sky130_fd_sc_hd__o211ai_2 _08666_ (.A1(_01620_),
    .A2(_07441_),
    .B1(_00202_),
    .C1(_00204_),
    .Y(_00209_));
 sky130_fd_sc_hd__a21o_1 _08667_ (.A1(_00202_),
    .A2(_00204_),
    .B1(_00206_),
    .X(_00210_));
 sky130_fd_sc_hd__nand4b_2 _08668_ (.A_N(_00197_),
    .B(_00200_),
    .C(_00207_),
    .D(_00208_),
    .Y(_00211_));
 sky130_fd_sc_hd__a2bb2oi_1 _08669_ (.A1_N(_00197_),
    .A2_N(_00199_),
    .B1(_00207_),
    .B2(_00208_),
    .Y(_00212_));
 sky130_fd_sc_hd__o211ai_4 _08670_ (.A1(_00197_),
    .A2(_00199_),
    .B1(_00209_),
    .C1(_00210_),
    .Y(_00213_));
 sky130_fd_sc_hd__o2bb2ai_1 _08671_ (.A1_N(_00211_),
    .A2_N(_00213_),
    .B1(_07543_),
    .B2(_00078_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand3b_1 _08672_ (.A_N(_00079_),
    .B(_00211_),
    .C(_00213_),
    .Y(_00215_));
 sky130_fd_sc_hd__o211ai_2 _08673_ (.A1(_07543_),
    .A2(_00078_),
    .B1(_00211_),
    .C1(_00213_),
    .Y(_00216_));
 sky130_fd_sc_hd__a21o_1 _08674_ (.A1(_00211_),
    .A2(_00213_),
    .B1(_00079_),
    .X(_00217_));
 sky130_fd_sc_hd__o211ai_4 _08675_ (.A1(_00080_),
    .A2(_00194_),
    .B1(_00216_),
    .C1(_00217_),
    .Y(_00218_));
 sky130_fd_sc_hd__and3_1 _08676_ (.A(_00214_),
    .B(_00215_),
    .C(_00195_),
    .X(_00219_));
 sky130_fd_sc_hd__nand3_2 _08677_ (.A(_00214_),
    .B(_00215_),
    .C(_00195_),
    .Y(_00220_));
 sky130_fd_sc_hd__a22oi_2 _08678_ (.A1(net33),
    .A2(_00193_),
    .B1(_00218_),
    .B2(_00220_),
    .Y(_00221_));
 sky130_fd_sc_hd__a32o_1 _08679_ (.A1(net33),
    .A2(_00189_),
    .A3(_00191_),
    .B1(_00218_),
    .B2(_00220_),
    .X(_00222_));
 sky130_fd_sc_hd__and4_1 _08680_ (.A(_00218_),
    .B(net33),
    .C(_00193_),
    .D(_00220_),
    .X(_00223_));
 sky130_fd_sc_hd__o21a_1 _08681_ (.A1(_00073_),
    .A2(_00087_),
    .B1(_00086_),
    .X(_00224_));
 sky130_fd_sc_hd__o221a_1 _08682_ (.A1(_00073_),
    .A2(_00087_),
    .B1(_00221_),
    .B2(_00223_),
    .C1(_00086_),
    .X(_00225_));
 sky130_fd_sc_hd__o21ai_2 _08683_ (.A1(_00221_),
    .A2(_00223_),
    .B1(_00224_),
    .Y(_00226_));
 sky130_fd_sc_hd__a41oi_4 _08684_ (.A1(_00193_),
    .A2(_00218_),
    .A3(_00220_),
    .A4(net33),
    .B1(_00224_),
    .Y(_00227_));
 sky130_fd_sc_hd__or3_1 _08685_ (.A(_00221_),
    .B(_00224_),
    .C(_00223_),
    .X(_00228_));
 sky130_fd_sc_hd__a2bb2oi_1 _08686_ (.A1_N(_00093_),
    .A2_N(_00098_),
    .B1(_00226_),
    .B2(_00228_),
    .Y(_00229_));
 sky130_fd_sc_hd__a2111oi_2 _08687_ (.A1(_00227_),
    .A2(_00222_),
    .B1(_00098_),
    .C1(_00093_),
    .D1(_00225_),
    .Y(_00230_));
 sky130_fd_sc_hd__nor2_1 _08688_ (.A(_00229_),
    .B(_00230_),
    .Y(_00231_));
 sky130_fd_sc_hd__or2_1 _08689_ (.A(_00229_),
    .B(_00230_),
    .X(_00232_));
 sky130_fd_sc_hd__nand3_1 _08690_ (.A(_00183_),
    .B(_00184_),
    .C(_00231_),
    .Y(_00233_));
 sky130_fd_sc_hd__o2bb2ai_1 _08691_ (.A1_N(_00183_),
    .A2_N(_00184_),
    .B1(_00229_),
    .B2(_00230_),
    .Y(_00234_));
 sky130_fd_sc_hd__a21o_1 _08692_ (.A1(_00183_),
    .A2(_00184_),
    .B1(_00232_),
    .X(_00235_));
 sky130_fd_sc_hd__o211ai_1 _08693_ (.A1(_00229_),
    .A2(_00230_),
    .B1(_00183_),
    .C1(_00184_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _08694_ (.A(_00235_),
    .B(_00236_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(_00233_),
    .B(_00234_),
    .Y(_00238_));
 sky130_fd_sc_hd__a21o_1 _08696_ (.A1(_00057_),
    .A2(_00101_),
    .B1(_00058_),
    .X(_00239_));
 sky130_fd_sc_hd__a21oi_2 _08697_ (.A1(_00057_),
    .A2(_00101_),
    .B1(_00058_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand3_1 _08698_ (.A(_00233_),
    .B(_00234_),
    .C(_00240_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand3_1 _08699_ (.A(_00235_),
    .B(_00236_),
    .C(_00239_),
    .Y(_00242_));
 sky130_fd_sc_hd__a22oi_1 _08700_ (.A1(_00109_),
    .A2(_00112_),
    .B1(_00241_),
    .B2(_00242_),
    .Y(_00243_));
 sky130_fd_sc_hd__and4_1 _08701_ (.A(_00109_),
    .B(_00112_),
    .C(_00241_),
    .D(_00242_),
    .X(_00244_));
 sky130_fd_sc_hd__nor2_1 _08702_ (.A(_00243_),
    .B(_00244_),
    .Y(_00245_));
 sky130_fd_sc_hd__xnor2_1 _08703_ (.A(_00117_),
    .B(_00245_),
    .Y(net69));
 sky130_fd_sc_hd__and3_1 _08704_ (.A(_00114_),
    .B(_00245_),
    .C(_00113_),
    .X(_00246_));
 sky130_fd_sc_hd__a21bo_1 _08705_ (.A1(_00183_),
    .A2(_00232_),
    .B1_N(_00184_),
    .X(_00247_));
 sky130_fd_sc_hd__a32o_1 _08706_ (.A1(_00129_),
    .A2(_00130_),
    .A3(_00182_),
    .B1(_00184_),
    .B2(_00231_),
    .X(_00248_));
 sky130_fd_sc_hd__o22a_1 _08707_ (.A1(_02636_),
    .A2(_06331_),
    .B1(net153),
    .B2(_01958_),
    .X(_00249_));
 sky130_fd_sc_hd__a32o_1 _08708_ (.A1(_02647_),
    .A2(_06309_),
    .A3(_06320_),
    .B1(_07370_),
    .B2(_01969_),
    .X(_00250_));
 sky130_fd_sc_hd__o31a_2 _08709_ (.A1(_02636_),
    .A2(net153),
    .A3(_00134_),
    .B1(_00250_),
    .X(_00251_));
 sky130_fd_sc_hd__or3_4 _08710_ (.A(_03906_),
    .B(_05381_),
    .C(_05403_),
    .X(_00252_));
 sky130_fd_sc_hd__xor2_4 _08711_ (.A(_00251_),
    .B(_00252_),
    .X(_00253_));
 sky130_fd_sc_hd__a21o_1 _08712_ (.A1(_00014_),
    .A2(_00162_),
    .B1(_00160_),
    .X(_00254_));
 sky130_fd_sc_hd__o22ai_4 _08713_ (.A1(net165),
    .A2(_07512_),
    .B1(_00009_),
    .B2(_00154_),
    .Y(_00255_));
 sky130_fd_sc_hd__a21oi_2 _08714_ (.A1(_00152_),
    .A2(_00255_),
    .B1(_00135_),
    .Y(_00256_));
 sky130_fd_sc_hd__a21o_1 _08715_ (.A1(_00152_),
    .A2(_00255_),
    .B1(_00135_),
    .X(_00257_));
 sky130_fd_sc_hd__nand3_2 _08716_ (.A(_00135_),
    .B(_00152_),
    .C(_00255_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _08717_ (.A(_00257_),
    .B(_00258_),
    .Y(_00259_));
 sky130_fd_sc_hd__and3_1 _08718_ (.A(_01499_),
    .B(_07509_),
    .C(_07511_),
    .X(_00260_));
 sky130_fd_sc_hd__a211o_1 _08719_ (.A1(_01434_),
    .A2(_01455_),
    .B1(_07508_),
    .C1(_07510_),
    .X(_00261_));
 sky130_fd_sc_hd__o221a_2 _08720_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_00003_),
    .B2(_00004_),
    .C1(_01172_),
    .X(_00262_));
 sky130_fd_sc_hd__nand4_4 _08721_ (.A(_06254_),
    .B(_07502_),
    .C(_00140_),
    .D(_00551_),
    .Y(_00263_));
 sky130_fd_sc_hd__a41oi_4 _08722_ (.A1(_06254_),
    .A2(_07502_),
    .A3(_00140_),
    .A4(_00551_),
    .B1(_00299_),
    .Y(_00264_));
 sky130_fd_sc_hd__a41o_2 _08723_ (.A1(_06254_),
    .A2(_07502_),
    .A3(_00140_),
    .A4(_00551_),
    .B1(_00299_),
    .X(_00265_));
 sky130_fd_sc_hd__o311a_1 _08724_ (.A1(_00141_),
    .A2(net37),
    .A3(_07505_),
    .B1(_00572_),
    .C1(net57),
    .X(_00266_));
 sky130_fd_sc_hd__a311o_4 _08725_ (.A1(net161),
    .A2(_00140_),
    .A3(_00551_),
    .B1(net38),
    .C1(_00299_),
    .X(_00267_));
 sky130_fd_sc_hd__a21oi_2 _08726_ (.A1(_00263_),
    .A2(net57),
    .B1(_00572_),
    .Y(_00268_));
 sky130_fd_sc_hd__a21o_2 _08727_ (.A1(_00263_),
    .A2(net57),
    .B1(_00572_),
    .X(_00269_));
 sky130_fd_sc_hd__a21oi_4 _08728_ (.A1(_00263_),
    .A2(net57),
    .B1(net38),
    .Y(_00270_));
 sky130_fd_sc_hd__a21o_4 _08729_ (.A1(_00263_),
    .A2(net57),
    .B1(net38),
    .X(_00271_));
 sky130_fd_sc_hd__o311a_4 _08730_ (.A1(_00141_),
    .A2(net37),
    .A3(_07505_),
    .B1(net38),
    .C1(net57),
    .X(_00272_));
 sky130_fd_sc_hd__a311o_4 _08731_ (.A1(net161),
    .A2(_00140_),
    .A3(_00551_),
    .B1(_00572_),
    .C1(_00299_),
    .X(_00273_));
 sky130_fd_sc_hd__nand2_8 _08732_ (.A(_00271_),
    .B(_00273_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_8 _08733_ (.A(_00267_),
    .B(_00269_),
    .Y(_00275_));
 sky130_fd_sc_hd__a31oi_1 _08734_ (.A1(_00263_),
    .A2(net38),
    .A3(net57),
    .B1(_00288_),
    .Y(_00276_));
 sky130_fd_sc_hd__a31o_1 _08735_ (.A1(_00263_),
    .A2(net38),
    .A3(net57),
    .B1(_00288_),
    .X(_00277_));
 sky130_fd_sc_hd__o21ai_1 _08736_ (.A1(net38),
    .A2(_00264_),
    .B1(_00276_),
    .Y(_00278_));
 sky130_fd_sc_hd__o32ai_4 _08737_ (.A1(_00987_),
    .A2(_00145_),
    .A3(_00147_),
    .B1(_00270_),
    .B2(_00277_),
    .Y(_00279_));
 sky130_fd_sc_hd__o2111ai_4 _08738_ (.A1(_00572_),
    .A2(_00265_),
    .B1(_00153_),
    .C1(net1),
    .D1(_00148_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand4_4 _08739_ (.A(_00150_),
    .B(_00271_),
    .C(_00273_),
    .D(_02177_),
    .Y(_00281_));
 sky130_fd_sc_hd__o311a_1 _08740_ (.A1(_00270_),
    .A2(_00272_),
    .A3(_00154_),
    .B1(_00279_),
    .C1(_00262_),
    .X(_00282_));
 sky130_fd_sc_hd__o2111ai_4 _08741_ (.A1(_00270_),
    .A2(_00280_),
    .B1(_00279_),
    .C1(net164),
    .D1(_00010_),
    .Y(_00283_));
 sky130_fd_sc_hd__a21oi_2 _08742_ (.A1(_00279_),
    .A2(_00281_),
    .B1(_00262_),
    .Y(_00284_));
 sky130_fd_sc_hd__a22o_2 _08743_ (.A1(net164),
    .A2(_00010_),
    .B1(_00279_),
    .B2(_00281_),
    .X(_00285_));
 sky130_fd_sc_hd__o21ai_1 _08744_ (.A1(_00282_),
    .A2(_00284_),
    .B1(_00260_),
    .Y(_00286_));
 sky130_fd_sc_hd__o211ai_1 _08745_ (.A1(_01488_),
    .A2(_07512_),
    .B1(_00283_),
    .C1(_00285_),
    .Y(_00287_));
 sky130_fd_sc_hd__o22ai_4 _08746_ (.A1(_01488_),
    .A2(_07512_),
    .B1(_00282_),
    .B2(_00284_),
    .Y(_00289_));
 sky130_fd_sc_hd__o2111ai_4 _08747_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_07513_),
    .C1(_00283_),
    .D1(_00285_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(_00289_),
    .B(_00290_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand3_1 _08749_ (.A(_00259_),
    .B(_00286_),
    .C(_00287_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand4_2 _08750_ (.A(_00257_),
    .B(_00258_),
    .C(_00289_),
    .D(_00290_),
    .Y(_00293_));
 sky130_fd_sc_hd__a21o_1 _08751_ (.A1(_00289_),
    .A2(_00290_),
    .B1(_00259_),
    .X(_00294_));
 sky130_fd_sc_hd__nand3_1 _08752_ (.A(_00259_),
    .B(_00289_),
    .C(_00290_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand4_4 _08753_ (.A(_00161_),
    .B(_00165_),
    .C(_00292_),
    .D(_00293_),
    .Y(_00296_));
 sky130_fd_sc_hd__and4_1 _08754_ (.A(_00254_),
    .B(_00294_),
    .C(_00295_),
    .D(_00253_),
    .X(_00297_));
 sky130_fd_sc_hd__a32oi_4 _08755_ (.A1(_00254_),
    .A2(_00294_),
    .A3(_00295_),
    .B1(_00296_),
    .B2(_00253_),
    .Y(_00298_));
 sky130_fd_sc_hd__o22ai_4 _08756_ (.A1(_00253_),
    .A2(_00296_),
    .B1(_00297_),
    .B2(_00298_),
    .Y(_00300_));
 sky130_fd_sc_hd__o22a_1 _08757_ (.A1(_00253_),
    .A2(_00296_),
    .B1(_00297_),
    .B2(_00298_),
    .X(_00301_));
 sky130_fd_sc_hd__a21bo_1 _08758_ (.A1(_00133_),
    .A2(_00169_),
    .B1_N(_00170_),
    .X(_00302_));
 sky130_fd_sc_hd__a21boi_4 _08759_ (.A1(_00169_),
    .A2(_00133_),
    .B1_N(_00170_),
    .Y(_00303_));
 sky130_fd_sc_hd__xnor2_1 _08760_ (.A(_00300_),
    .B(_00303_),
    .Y(_00304_));
 sky130_fd_sc_hd__o2bb2ai_1 _08761_ (.A1_N(_00176_),
    .A2_N(_00172_),
    .B1(_00026_),
    .B2(_00179_),
    .Y(_00305_));
 sky130_fd_sc_hd__o2bb2a_1 _08762_ (.A1_N(_00175_),
    .A2_N(_00180_),
    .B1(_00177_),
    .B2(_00171_),
    .X(_00306_));
 sky130_fd_sc_hd__xnor2_2 _08763_ (.A(_00304_),
    .B(_00306_),
    .Y(_00307_));
 sky130_fd_sc_hd__and3_1 _08764_ (.A(_04222_),
    .B(_04233_),
    .C(_04726_),
    .X(_00308_));
 sky130_fd_sc_hd__o21ai_4 _08765_ (.A1(_00118_),
    .A2(_00121_),
    .B1(_00120_),
    .Y(_00309_));
 sky130_fd_sc_hd__or4b_2 _08766_ (.A(_04244_),
    .B(_04671_),
    .C(_04693_),
    .D_N(_00309_),
    .X(_00311_));
 sky130_fd_sc_hd__a31o_1 _08767_ (.A1(_04222_),
    .A2(_04233_),
    .A3(_04726_),
    .B1(_00309_),
    .X(_00312_));
 sky130_fd_sc_hd__and2_1 _08768_ (.A(_00311_),
    .B(_00312_),
    .X(_00313_));
 sky130_fd_sc_hd__nand2_1 _08769_ (.A(_00311_),
    .B(_00312_),
    .Y(_00314_));
 sky130_fd_sc_hd__o211ai_2 _08770_ (.A1(_00124_),
    .A2(_00040_),
    .B1(_00046_),
    .C1(_00128_),
    .Y(_00315_));
 sky130_fd_sc_hd__o221ai_4 _08771_ (.A1(_00043_),
    .A2(_00047_),
    .B1(_00123_),
    .B2(_00041_),
    .C1(_00127_),
    .Y(_00316_));
 sky130_fd_sc_hd__o211ai_1 _08772_ (.A1(_00041_),
    .A2(_00123_),
    .B1(_00314_),
    .C1(_00315_),
    .Y(_00317_));
 sky130_fd_sc_hd__o211ai_1 _08773_ (.A1(_00040_),
    .A2(_00124_),
    .B1(_00313_),
    .C1(_00316_),
    .Y(_00318_));
 sky130_fd_sc_hd__o211ai_2 _08774_ (.A1(_00040_),
    .A2(_00124_),
    .B1(_00314_),
    .C1(_00316_),
    .Y(_00319_));
 sky130_fd_sc_hd__o211ai_2 _08775_ (.A1(_00041_),
    .A2(_00123_),
    .B1(_00313_),
    .C1(_00315_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand3_4 _08776_ (.A(_00319_),
    .B(_00320_),
    .C(_00307_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand3b_2 _08777_ (.A_N(_00307_),
    .B(_00317_),
    .C(_00318_),
    .Y(_00323_));
 sky130_fd_sc_hd__o2bb2ai_2 _08778_ (.A1_N(_00222_),
    .A2_N(_00227_),
    .B1(_00093_),
    .B2(_00098_),
    .Y(_00324_));
 sky130_fd_sc_hd__a31o_1 _08779_ (.A1(net33),
    .A2(_00193_),
    .A3(_00218_),
    .B1(_00219_),
    .X(_00325_));
 sky130_fd_sc_hd__inv_2 _08780_ (.A(_00325_),
    .Y(_00326_));
 sky130_fd_sc_hd__o21ai_1 _08781_ (.A1(_00079_),
    .A2(_00212_),
    .B1(_00211_),
    .Y(_00327_));
 sky130_fd_sc_hd__o211a_1 _08782_ (.A1(_00203_),
    .A2(_00205_),
    .B1(_00197_),
    .C1(_00202_),
    .X(_00328_));
 sky130_fd_sc_hd__o211ai_1 _08783_ (.A1(_00203_),
    .A2(_00205_),
    .B1(_00197_),
    .C1(_00202_),
    .Y(_00329_));
 sky130_fd_sc_hd__a311oi_2 _08784_ (.A1(_01631_),
    .A2(_07440_),
    .A3(_00202_),
    .B1(_00203_),
    .C1(_00197_),
    .Y(_00330_));
 sky130_fd_sc_hd__a311o_1 _08785_ (.A1(_01631_),
    .A2(_07440_),
    .A3(_00202_),
    .B1(_00203_),
    .C1(_00197_),
    .X(_00331_));
 sky130_fd_sc_hd__a22o_2 _08786_ (.A1(_01543_),
    .A2(_01565_),
    .B1(_07534_),
    .B2(_07535_),
    .X(_00333_));
 sky130_fd_sc_hd__o2111ai_4 _08787_ (.A1(_00299_),
    .A2(_03511_),
    .B1(_05272_),
    .C1(_05283_),
    .D1(_03490_),
    .Y(_00334_));
 sky130_fd_sc_hd__o21ai_4 _08788_ (.A1(net159),
    .A2(_07189_),
    .B1(_00334_),
    .Y(_00335_));
 sky130_fd_sc_hd__o21ai_4 _08789_ (.A1(_07125_),
    .A2(_07135_),
    .B1(_03555_),
    .Y(_00336_));
 sky130_fd_sc_hd__and4_1 _08790_ (.A(_05316_),
    .B(_07200_),
    .C(_02866_),
    .D(net157),
    .X(_00337_));
 sky130_fd_sc_hd__nand4_2 _08791_ (.A(_05316_),
    .B(_07200_),
    .C(_02866_),
    .D(net157),
    .Y(_00338_));
 sky130_fd_sc_hd__a22oi_2 _08792_ (.A1(_07440_),
    .A2(_02133_),
    .B1(_00338_),
    .B2(_00335_),
    .Y(_00339_));
 sky130_fd_sc_hd__o2bb2ai_2 _08793_ (.A1_N(_00335_),
    .A2_N(_00338_),
    .B1(_02122_),
    .B2(_07441_),
    .Y(_00340_));
 sky130_fd_sc_hd__o2111a_1 _08794_ (.A1(_00201_),
    .A2(_00336_),
    .B1(_07440_),
    .C1(_00335_),
    .D1(_02133_),
    .X(_00341_));
 sky130_fd_sc_hd__o2111ai_4 _08795_ (.A1(_00201_),
    .A2(_00336_),
    .B1(_07440_),
    .C1(_00335_),
    .D1(_02133_),
    .Y(_00342_));
 sky130_fd_sc_hd__o2111ai_2 _08796_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_07540_),
    .C1(_00340_),
    .D1(_00342_),
    .Y(_00344_));
 sky130_fd_sc_hd__a22o_1 _08797_ (.A1(_01631_),
    .A2(_07540_),
    .B1(_00340_),
    .B2(_00342_),
    .X(_00345_));
 sky130_fd_sc_hd__o21bai_1 _08798_ (.A1(_00339_),
    .A2(_00341_),
    .B1_N(_00333_),
    .Y(_00346_));
 sky130_fd_sc_hd__o211ai_1 _08799_ (.A1(_01620_),
    .A2(net150),
    .B1(_00340_),
    .C1(_00342_),
    .Y(_00347_));
 sky130_fd_sc_hd__o211ai_1 _08800_ (.A1(_00328_),
    .A2(_00330_),
    .B1(_00346_),
    .C1(_00347_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand4_1 _08801_ (.A(_00329_),
    .B(_00331_),
    .C(_00344_),
    .D(_00345_),
    .Y(_00349_));
 sky130_fd_sc_hd__o211ai_1 _08802_ (.A1(_00328_),
    .A2(_00330_),
    .B1(_00344_),
    .C1(_00345_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand4_1 _08803_ (.A(_00329_),
    .B(_00331_),
    .C(_00346_),
    .D(_00347_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand3_1 _08804_ (.A(_00349_),
    .B(_00327_),
    .C(_00348_),
    .Y(_00352_));
 sky130_fd_sc_hd__nand3b_1 _08805_ (.A_N(_00327_),
    .B(_00350_),
    .C(_00351_),
    .Y(_00353_));
 sky130_fd_sc_hd__o211ai_4 _08806_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_00189_),
    .C1(_00191_),
    .Y(_00355_));
 sky130_fd_sc_hd__a32o_1 _08807_ (.A1(_00911_),
    .A2(_00189_),
    .A3(_00191_),
    .B1(_01303_),
    .B2(_00072_),
    .X(_00356_));
 sky130_fd_sc_hd__nor2_1 _08808_ (.A(_00196_),
    .B(_00355_),
    .Y(_00357_));
 sky130_fd_sc_hd__o31ai_1 _08809_ (.A1(_01292_),
    .A2(_00192_),
    .A3(_00198_),
    .B1(_00356_),
    .Y(_00358_));
 sky130_fd_sc_hd__nor2_1 _08810_ (.A(net5),
    .B(_00185_),
    .Y(_00359_));
 sky130_fd_sc_hd__nand4_2 _08811_ (.A(_07435_),
    .B(_00062_),
    .C(_00540_),
    .D(_00561_),
    .Y(_00360_));
 sky130_fd_sc_hd__o211a_4 _08812_ (.A1(net5),
    .A2(_00185_),
    .B1(net6),
    .C1(net174),
    .X(_00361_));
 sky130_fd_sc_hd__o211ai_4 _08813_ (.A1(net5),
    .A2(_00185_),
    .B1(net6),
    .C1(net174),
    .Y(_00362_));
 sky130_fd_sc_hd__a21oi_4 _08814_ (.A1(_00360_),
    .A2(net174),
    .B1(net6),
    .Y(_00363_));
 sky130_fd_sc_hd__a21o_4 _08815_ (.A1(_00360_),
    .A2(net174),
    .B1(net6),
    .X(_00364_));
 sky130_fd_sc_hd__nand2_8 _08816_ (.A(_00362_),
    .B(_00364_),
    .Y(_00366_));
 sky130_fd_sc_hd__nor2_8 _08817_ (.A(_00361_),
    .B(_00363_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand3_1 _08818_ (.A(_00364_),
    .B(net33),
    .C(_00362_),
    .Y(_00368_));
 sky130_fd_sc_hd__and4b_1 _08819_ (.A_N(_00357_),
    .B(net33),
    .C(_00356_),
    .D(_00367_),
    .X(_00369_));
 sky130_fd_sc_hd__o31a_1 _08820_ (.A1(_00310_),
    .A2(_00361_),
    .A3(_00363_),
    .B1(_00358_),
    .X(_00370_));
 sky130_fd_sc_hd__and3_1 _08821_ (.A(_00358_),
    .B(_00367_),
    .C(net33),
    .X(_00371_));
 sky130_fd_sc_hd__o311a_1 _08822_ (.A1(_01292_),
    .A2(_00192_),
    .A3(_00198_),
    .B1(_00356_),
    .C1(_00368_),
    .X(_00372_));
 sky130_fd_sc_hd__nor2_1 _08823_ (.A(_00369_),
    .B(_00370_),
    .Y(_00373_));
 sky130_fd_sc_hd__o2bb2ai_1 _08824_ (.A1_N(_00352_),
    .A2_N(_00353_),
    .B1(_00371_),
    .B2(_00372_),
    .Y(_00374_));
 sky130_fd_sc_hd__o211ai_2 _08825_ (.A1(_00369_),
    .A2(_00370_),
    .B1(_00352_),
    .C1(_00353_),
    .Y(_00375_));
 sky130_fd_sc_hd__and2_1 _08826_ (.A(_00374_),
    .B(_00375_),
    .X(_00377_));
 sky130_fd_sc_hd__nand2_1 _08827_ (.A(_00374_),
    .B(_00375_),
    .Y(_00378_));
 sky130_fd_sc_hd__xnor2_1 _08828_ (.A(_00325_),
    .B(_00378_),
    .Y(_00379_));
 sky130_fd_sc_hd__o311a_1 _08829_ (.A1(_00093_),
    .A2(_00098_),
    .A3(_00225_),
    .B1(_00228_),
    .C1(_00379_),
    .X(_00380_));
 sky130_fd_sc_hd__and3b_1 _08830_ (.A_N(_00379_),
    .B(_00324_),
    .C(_00226_),
    .X(_00381_));
 sky130_fd_sc_hd__and3_1 _08831_ (.A(_00226_),
    .B(_00324_),
    .C(_00379_),
    .X(_00382_));
 sky130_fd_sc_hd__a21oi_1 _08832_ (.A1(_00226_),
    .A2(_00324_),
    .B1(_00379_),
    .Y(_00383_));
 sky130_fd_sc_hd__o211ai_2 _08833_ (.A1(_00380_),
    .A2(_00381_),
    .B1(_00322_),
    .C1(_00323_),
    .Y(_00384_));
 sky130_fd_sc_hd__o2bb2ai_1 _08834_ (.A1_N(_00322_),
    .A2_N(_00323_),
    .B1(_00382_),
    .B2(_00383_),
    .Y(_00385_));
 sky130_fd_sc_hd__o2bb2ai_1 _08835_ (.A1_N(_00322_),
    .A2_N(_00323_),
    .B1(_00380_),
    .B2(_00381_),
    .Y(_00386_));
 sky130_fd_sc_hd__o211ai_1 _08836_ (.A1(_00382_),
    .A2(_00383_),
    .B1(_00322_),
    .C1(_00323_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _08837_ (.A(_00384_),
    .B(_00385_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand3_1 _08838_ (.A(_00385_),
    .B(_00247_),
    .C(_00384_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand3_2 _08839_ (.A(_00248_),
    .B(_00386_),
    .C(_00388_),
    .Y(_00391_));
 sky130_fd_sc_hd__o211ai_2 _08840_ (.A1(_07578_),
    .A2(_00106_),
    .B1(_00112_),
    .C1(_00241_),
    .Y(_00392_));
 sky130_fd_sc_hd__o211ai_1 _08841_ (.A1(_07579_),
    .A2(_00107_),
    .B1(_00111_),
    .C1(_00242_),
    .Y(_00393_));
 sky130_fd_sc_hd__o21ai_1 _08842_ (.A1(_00237_),
    .A2(_00240_),
    .B1(_00392_),
    .Y(_00394_));
 sky130_fd_sc_hd__a21oi_1 _08843_ (.A1(_00390_),
    .A2(_00391_),
    .B1(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__and3_1 _08844_ (.A(_00390_),
    .B(_00391_),
    .C(_00394_),
    .X(_00396_));
 sky130_fd_sc_hd__nor2_1 _08845_ (.A(_00395_),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__a311o_1 _08846_ (.A1(_00114_),
    .A2(_00245_),
    .A3(_00113_),
    .B1(_00834_),
    .C1(_00397_),
    .X(_00399_));
 sky130_fd_sc_hd__o21ai_1 _08847_ (.A1(_00834_),
    .A2(_00246_),
    .B1(_00397_),
    .Y(_00400_));
 sky130_fd_sc_hd__and2_1 _08848_ (.A(_00399_),
    .B(_00400_),
    .X(net70));
 sky130_fd_sc_hd__or3b_1 _08849_ (.A(_00395_),
    .B(_00396_),
    .C_N(_00246_),
    .X(_00401_));
 sky130_fd_sc_hd__o21ai_2 _08850_ (.A1(_00382_),
    .A2(_00383_),
    .B1(_00323_),
    .Y(_00402_));
 sky130_fd_sc_hd__o31ai_2 _08851_ (.A1(_02636_),
    .A2(net153),
    .A3(_00134_),
    .B1(_00252_),
    .Y(_00403_));
 sky130_fd_sc_hd__o32a_1 _08852_ (.A1(_02636_),
    .A2(net153),
    .A3(_00134_),
    .B1(_00252_),
    .B2(_00249_),
    .X(_00404_));
 sky130_fd_sc_hd__a31oi_1 _08853_ (.A1(_00281_),
    .A2(_00262_),
    .A3(_00279_),
    .B1(_00260_),
    .Y(_00405_));
 sky130_fd_sc_hd__a31o_1 _08854_ (.A1(_00281_),
    .A2(_00262_),
    .A3(_00279_),
    .B1(_00260_),
    .X(_00406_));
 sky130_fd_sc_hd__a22oi_4 _08855_ (.A1(_00250_),
    .A2(_00403_),
    .B1(_00406_),
    .B2(_00285_),
    .Y(_00407_));
 sky130_fd_sc_hd__nor3_1 _08856_ (.A(_00284_),
    .B(_00404_),
    .C(_00405_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2_1 _08857_ (.A(_00407_),
    .B(_00409_),
    .Y(_00410_));
 sky130_fd_sc_hd__o211ai_4 _08858_ (.A1(_01892_),
    .A2(_01914_),
    .B1(_07509_),
    .C1(_07511_),
    .Y(_00411_));
 sky130_fd_sc_hd__or4_2 _08859_ (.A(_01488_),
    .B(_00005_),
    .C(_00007_),
    .D(_00411_),
    .X(_00412_));
 sky130_fd_sc_hd__a32o_1 _08860_ (.A1(_01499_),
    .A2(_00006_),
    .A3(_00008_),
    .B1(_01969_),
    .B2(_07513_),
    .X(_00413_));
 sky130_fd_sc_hd__o311a_1 _08861_ (.A1(_01488_),
    .A2(_00005_),
    .A3(_00007_),
    .B1(_01969_),
    .C1(_07513_),
    .X(_00414_));
 sky130_fd_sc_hd__o311a_1 _08862_ (.A1(_01958_),
    .A2(_07508_),
    .A3(_07510_),
    .B1(_00010_),
    .C1(_01499_),
    .X(_00415_));
 sky130_fd_sc_hd__o31a_1 _08863_ (.A1(_01958_),
    .A2(_00009_),
    .A3(_00261_),
    .B1(_00413_),
    .X(_00416_));
 sky130_fd_sc_hd__o221a_1 _08864_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_00144_),
    .B2(_00142_),
    .C1(_01172_),
    .X(_00417_));
 sky130_fd_sc_hd__and3_1 _08865_ (.A(net164),
    .B(_00146_),
    .C(_00148_),
    .X(_00418_));
 sky130_fd_sc_hd__nand4_2 _08866_ (.A(net161),
    .B(_00140_),
    .C(_00551_),
    .D(_00572_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _08867_ (.A(net57),
    .B(net38),
    .Y(_00421_));
 sky130_fd_sc_hd__o211ai_4 _08868_ (.A1(net38),
    .A2(_00263_),
    .B1(_00583_),
    .C1(net57),
    .Y(_00422_));
 sky130_fd_sc_hd__nand3_4 _08869_ (.A(_00265_),
    .B(_00421_),
    .C(net39),
    .Y(_00423_));
 sky130_fd_sc_hd__a41o_4 _08870_ (.A1(net161),
    .A2(_00140_),
    .A3(_00551_),
    .A4(_00572_),
    .B1(_00583_),
    .X(_00424_));
 sky130_fd_sc_hd__o211ai_4 _08871_ (.A1(net38),
    .A2(_00263_),
    .B1(net39),
    .C1(net57),
    .Y(_00425_));
 sky130_fd_sc_hd__a21oi_2 _08872_ (.A1(_00420_),
    .A2(net57),
    .B1(net39),
    .Y(_00426_));
 sky130_fd_sc_hd__o211ai_4 _08873_ (.A1(_00299_),
    .A2(_00572_),
    .B1(_00583_),
    .C1(_00265_),
    .Y(_00427_));
 sky130_fd_sc_hd__o21ai_4 _08874_ (.A1(_00299_),
    .A2(_00424_),
    .B1(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_8 _08875_ (.A(_00422_),
    .B(_00423_),
    .Y(_00429_));
 sky130_fd_sc_hd__a31o_1 _08876_ (.A1(_00420_),
    .A2(net39),
    .A3(net57),
    .B1(_00987_),
    .X(_00431_));
 sky130_fd_sc_hd__o22a_2 _08877_ (.A1(net172),
    .A2(_00943_),
    .B1(_00264_),
    .B2(net38),
    .X(_00432_));
 sky130_fd_sc_hd__o211ai_4 _08878_ (.A1(net172),
    .A2(_00943_),
    .B1(_00271_),
    .C1(_00273_),
    .Y(_00433_));
 sky130_fd_sc_hd__nor3_2 _08879_ (.A(_00426_),
    .B(_00431_),
    .C(_00278_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand4_4 _08880_ (.A(_00273_),
    .B(_00429_),
    .C(_00432_),
    .D(net1),
    .Y(_00435_));
 sky130_fd_sc_hd__a32oi_4 _08881_ (.A1(_00427_),
    .A2(net1),
    .A3(_00425_),
    .B1(_00432_),
    .B2(_00273_),
    .Y(_00436_));
 sky130_fd_sc_hd__o32ai_4 _08882_ (.A1(_00987_),
    .A2(_00270_),
    .A3(_00272_),
    .B1(_00288_),
    .B2(_00428_),
    .Y(_00437_));
 sky130_fd_sc_hd__o2bb2ai_4 _08883_ (.A1_N(_00417_),
    .A2_N(_00148_),
    .B1(_00436_),
    .B2(_00434_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand3_4 _08884_ (.A(_00435_),
    .B(_00437_),
    .C(_00418_),
    .Y(_00439_));
 sky130_fd_sc_hd__a22oi_4 _08885_ (.A1(_00412_),
    .A2(_00413_),
    .B1(_00438_),
    .B2(_00439_),
    .Y(_00440_));
 sky130_fd_sc_hd__a22o_1 _08886_ (.A1(_00412_),
    .A2(_00413_),
    .B1(_00438_),
    .B2(_00439_),
    .X(_00442_));
 sky130_fd_sc_hd__o211a_1 _08887_ (.A1(_00414_),
    .A2(_00415_),
    .B1(_00438_),
    .C1(_00439_),
    .X(_00443_));
 sky130_fd_sc_hd__nand3_2 _08888_ (.A(_00438_),
    .B(_00439_),
    .C(_00416_),
    .Y(_00444_));
 sky130_fd_sc_hd__o32ai_4 _08889_ (.A1(_02188_),
    .A2(net143),
    .A3(_00274_),
    .B1(_00440_),
    .B2(_00443_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand3b_1 _08890_ (.A_N(_00281_),
    .B(_00442_),
    .C(_00444_),
    .Y(_00446_));
 sky130_fd_sc_hd__o21bai_1 _08891_ (.A1(_00440_),
    .A2(_00443_),
    .B1_N(_00281_),
    .Y(_00447_));
 sky130_fd_sc_hd__o211ai_2 _08892_ (.A1(_00280_),
    .A2(_00270_),
    .B1(_00444_),
    .C1(_00442_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _08893_ (.A(_00445_),
    .B(_00446_),
    .Y(_00449_));
 sky130_fd_sc_hd__o211ai_1 _08894_ (.A1(_00407_),
    .A2(_00409_),
    .B1(_00447_),
    .C1(_00448_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand3_1 _08895_ (.A(_00445_),
    .B(_00446_),
    .C(_00410_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand3_1 _08896_ (.A(_00447_),
    .B(_00448_),
    .C(_00410_),
    .Y(_00453_));
 sky130_fd_sc_hd__o211ai_2 _08897_ (.A1(_00407_),
    .A2(_00409_),
    .B1(_00445_),
    .C1(_00446_),
    .Y(_00454_));
 sky130_fd_sc_hd__o21ai_1 _08898_ (.A1(_00256_),
    .A2(_00291_),
    .B1(_00258_),
    .Y(_00455_));
 sky130_fd_sc_hd__o2111ai_4 _08899_ (.A1(_00256_),
    .A2(_00291_),
    .B1(_00453_),
    .C1(_00454_),
    .D1(_00258_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand3_2 _08900_ (.A(_00450_),
    .B(_00451_),
    .C(_00455_),
    .Y(_00457_));
 sky130_fd_sc_hd__or3_1 _08901_ (.A(_04244_),
    .B(_05381_),
    .C(_05403_),
    .X(_00458_));
 sky130_fd_sc_hd__nor4_1 _08902_ (.A(_02636_),
    .B(_03906_),
    .C(_06331_),
    .D(net153),
    .Y(_00459_));
 sky130_fd_sc_hd__o22ai_1 _08903_ (.A1(_03906_),
    .A2(_06331_),
    .B1(net153),
    .B2(_02636_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2b_1 _08904_ (.A_N(_00459_),
    .B(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__xor2_1 _08905_ (.A(_00458_),
    .B(_00461_),
    .X(_00462_));
 sky130_fd_sc_hd__xnor2_1 _08906_ (.A(_00458_),
    .B(_00461_),
    .Y(_00464_));
 sky130_fd_sc_hd__a21o_1 _08907_ (.A1(_00456_),
    .A2(_00457_),
    .B1(_00464_),
    .X(_00465_));
 sky130_fd_sc_hd__nand3_1 _08908_ (.A(_00456_),
    .B(_00457_),
    .C(_00464_),
    .Y(_00466_));
 sky130_fd_sc_hd__a21o_1 _08909_ (.A1(_00456_),
    .A2(_00457_),
    .B1(_00462_),
    .X(_00467_));
 sky130_fd_sc_hd__nand3_1 _08910_ (.A(_00456_),
    .B(_00457_),
    .C(_00462_),
    .Y(_00468_));
 sky130_fd_sc_hd__nand3_2 _08911_ (.A(_00467_),
    .B(_00468_),
    .C(_00298_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand3b_4 _08912_ (.A_N(_00298_),
    .B(_00465_),
    .C(_00466_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _08913_ (.A(_00469_),
    .B(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__o211ai_2 _08914_ (.A1(_00300_),
    .A2(_00302_),
    .B1(_00305_),
    .C1(_00175_),
    .Y(_00472_));
 sky130_fd_sc_hd__o2bb2ai_1 _08915_ (.A1_N(_00175_),
    .A2_N(_00305_),
    .B1(_00303_),
    .B2(_00301_),
    .Y(_00473_));
 sky130_fd_sc_hd__o211ai_2 _08916_ (.A1(_00300_),
    .A2(_00302_),
    .B1(_00470_),
    .C1(_00473_),
    .Y(_00475_));
 sky130_fd_sc_hd__o2111a_1 _08917_ (.A1(_00301_),
    .A2(_00303_),
    .B1(_00469_),
    .C1(_00470_),
    .D1(_00472_),
    .X(_00476_));
 sky130_fd_sc_hd__o211a_1 _08918_ (.A1(_00300_),
    .A2(_00302_),
    .B1(_00471_),
    .C1(_00473_),
    .X(_00477_));
 sky130_fd_sc_hd__o211ai_2 _08919_ (.A1(_00040_),
    .A2(_00124_),
    .B1(_00311_),
    .C1(_00316_),
    .Y(_00478_));
 sky130_fd_sc_hd__o211ai_1 _08920_ (.A1(_00041_),
    .A2(_00123_),
    .B1(_00312_),
    .C1(_00315_),
    .Y(_00479_));
 sky130_fd_sc_hd__o221ai_4 _08921_ (.A1(_00308_),
    .A2(_00309_),
    .B1(_00476_),
    .B2(_00477_),
    .C1(_00478_),
    .Y(_00480_));
 sky130_fd_sc_hd__a311oi_1 _08922_ (.A1(_04255_),
    .A2(_04726_),
    .A3(_00309_),
    .B1(_00476_),
    .C1(_00477_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _08923_ (.A(_00479_),
    .B(_00481_),
    .Y(_00482_));
 sky130_fd_sc_hd__a32o_1 _08924_ (.A1(_00327_),
    .A2(_00348_),
    .A3(_00349_),
    .B1(_00373_),
    .B2(_00353_),
    .X(_00483_));
 sky130_fd_sc_hd__a31o_1 _08925_ (.A1(_00331_),
    .A2(_00344_),
    .A3(_00345_),
    .B1(_00328_),
    .X(_00484_));
 sky130_fd_sc_hd__a21oi_1 _08926_ (.A1(_00196_),
    .A2(_00355_),
    .B1(_00368_),
    .Y(_00486_));
 sky130_fd_sc_hd__nor2_1 _08927_ (.A(_00357_),
    .B(_00486_),
    .Y(_00487_));
 sky130_fd_sc_hd__o21ai_1 _08928_ (.A1(_01620_),
    .A2(net150),
    .B1(_00342_),
    .Y(_00488_));
 sky130_fd_sc_hd__o311a_1 _08929_ (.A1(_01620_),
    .A2(net150),
    .A3(_00339_),
    .B1(_00342_),
    .C1(_00487_),
    .X(_00489_));
 sky130_fd_sc_hd__o211ai_2 _08930_ (.A1(_00333_),
    .A2(_00339_),
    .B1(_00342_),
    .C1(_00487_),
    .Y(_00490_));
 sky130_fd_sc_hd__o211a_1 _08931_ (.A1(_00357_),
    .A2(_00486_),
    .B1(_00488_),
    .C1(_00340_),
    .X(_00491_));
 sky130_fd_sc_hd__o211ai_1 _08932_ (.A1(_00357_),
    .A2(_00486_),
    .B1(_00488_),
    .C1(_00340_),
    .Y(_00492_));
 sky130_fd_sc_hd__o221ai_4 _08933_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_00063_),
    .B2(_00066_),
    .C1(_00070_),
    .Y(_00493_));
 sky130_fd_sc_hd__o21ai_1 _08934_ (.A1(_02122_),
    .A2(net150),
    .B1(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__a22oi_2 _08935_ (.A1(_02046_),
    .A2(_02068_),
    .B1(_00065_),
    .B2(_00540_),
    .Y(_00495_));
 sky130_fd_sc_hd__o21ai_4 _08936_ (.A1(_00063_),
    .A2(_00066_),
    .B1(_00495_),
    .Y(_00497_));
 sky130_fd_sc_hd__o31a_1 _08937_ (.A1(_01620_),
    .A2(net150),
    .A3(_00497_),
    .B1(_00494_),
    .X(_00498_));
 sky130_fd_sc_hd__o21ai_1 _08938_ (.A1(_00333_),
    .A2(_00497_),
    .B1(_00494_),
    .Y(_00499_));
 sky130_fd_sc_hd__and3_1 _08939_ (.A(_02866_),
    .B(net162),
    .C(net154),
    .X(_00500_));
 sky130_fd_sc_hd__a32oi_4 _08940_ (.A1(_03555_),
    .A2(_07157_),
    .A3(_07178_),
    .B1(_05316_),
    .B2(_04726_),
    .Y(_00501_));
 sky130_fd_sc_hd__a32o_1 _08941_ (.A1(_03555_),
    .A2(_07157_),
    .A3(_07178_),
    .B1(_05316_),
    .B2(_04726_),
    .X(_00502_));
 sky130_fd_sc_hd__o2111ai_4 _08942_ (.A1(_04606_),
    .A2(_04660_),
    .B1(_04704_),
    .C1(_07157_),
    .D1(_07178_),
    .Y(_00503_));
 sky130_fd_sc_hd__nor2_1 _08943_ (.A(_00334_),
    .B(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__o22ai_1 _08944_ (.A1(net159),
    .A2(_07441_),
    .B1(_00501_),
    .B2(_00504_),
    .Y(_00505_));
 sky130_fd_sc_hd__o2111ai_1 _08945_ (.A1(_00334_),
    .A2(_00503_),
    .B1(_07440_),
    .C1(_00502_),
    .D1(_02866_),
    .Y(_00506_));
 sky130_fd_sc_hd__o21ai_1 _08946_ (.A1(_00501_),
    .A2(_00504_),
    .B1(_00500_),
    .Y(_00508_));
 sky130_fd_sc_hd__o221ai_2 _08947_ (.A1(net159),
    .A2(_07441_),
    .B1(_00334_),
    .B2(_00503_),
    .C1(_00502_),
    .Y(_00509_));
 sky130_fd_sc_hd__and3_1 _08948_ (.A(_00499_),
    .B(_00508_),
    .C(_00509_),
    .X(_00510_));
 sky130_fd_sc_hd__nand3_2 _08949_ (.A(_00499_),
    .B(_00508_),
    .C(_00509_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand3_2 _08950_ (.A(_00498_),
    .B(_00505_),
    .C(_00506_),
    .Y(_00512_));
 sky130_fd_sc_hd__o21ai_2 _08951_ (.A1(_00201_),
    .A2(_00336_),
    .B1(_00512_),
    .Y(_00513_));
 sky130_fd_sc_hd__a21o_1 _08952_ (.A1(_00511_),
    .A2(_00512_),
    .B1(_00338_),
    .X(_00514_));
 sky130_fd_sc_hd__a21o_1 _08953_ (.A1(_00511_),
    .A2(_00512_),
    .B1(_00337_),
    .X(_00515_));
 sky130_fd_sc_hd__nand3_1 _08954_ (.A(_00511_),
    .B(_00512_),
    .C(_00337_),
    .Y(_00516_));
 sky130_fd_sc_hd__nand4_1 _08955_ (.A(_00490_),
    .B(_00492_),
    .C(_00515_),
    .D(_00516_),
    .Y(_00517_));
 sky130_fd_sc_hd__o221ai_1 _08956_ (.A1(_00513_),
    .A2(_00510_),
    .B1(_00491_),
    .B2(_00489_),
    .C1(_00514_),
    .Y(_00519_));
 sky130_fd_sc_hd__o2111ai_1 _08957_ (.A1(_00513_),
    .A2(_00510_),
    .B1(_00492_),
    .C1(_00490_),
    .D1(_00514_),
    .Y(_00520_));
 sky130_fd_sc_hd__o211ai_1 _08958_ (.A1(_00489_),
    .A2(_00491_),
    .B1(_00515_),
    .C1(_00516_),
    .Y(_00521_));
 sky130_fd_sc_hd__nand3_1 _08959_ (.A(_00517_),
    .B(_00519_),
    .C(_00484_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand3b_2 _08960_ (.A_N(_00484_),
    .B(_00520_),
    .C(_00521_),
    .Y(_00523_));
 sky130_fd_sc_hd__nor2_4 _08961_ (.A(net5),
    .B(net6),
    .Y(_00524_));
 sky130_fd_sc_hd__or2_2 _08962_ (.A(net5),
    .B(net6),
    .X(_00525_));
 sky130_fd_sc_hd__nand4_4 _08963_ (.A(_07435_),
    .B(_00062_),
    .C(_00524_),
    .D(_00540_),
    .Y(_00526_));
 sky130_fd_sc_hd__a21oi_4 _08964_ (.A1(_00526_),
    .A2(net174),
    .B1(net7),
    .Y(_00527_));
 sky130_fd_sc_hd__a21o_2 _08965_ (.A1(_00526_),
    .A2(net174),
    .B1(net7),
    .X(_00528_));
 sky130_fd_sc_hd__o31a_4 _08966_ (.A1(net5),
    .A2(net6),
    .A3(_00185_),
    .B1(net7),
    .X(_00530_));
 sky130_fd_sc_hd__nand2_4 _08967_ (.A(net25),
    .B(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__a21o_4 _08968_ (.A1(net174),
    .A2(_00530_),
    .B1(_00527_),
    .X(_00532_));
 sky130_fd_sc_hd__a21oi_4 _08969_ (.A1(net25),
    .A2(_00530_),
    .B1(_00527_),
    .Y(_00533_));
 sky130_fd_sc_hd__o32ai_2 _08970_ (.A1(_00900_),
    .A2(_00361_),
    .A3(_00363_),
    .B1(_01292_),
    .B2(_00192_),
    .Y(_00534_));
 sky130_fd_sc_hd__o31a_1 _08971_ (.A1(_01292_),
    .A2(_00355_),
    .A3(_00366_),
    .B1(_00534_),
    .X(_00535_));
 sky130_fd_sc_hd__a21oi_1 _08972_ (.A1(net33),
    .A2(_00533_),
    .B1(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__and3_1 _08973_ (.A(net33),
    .B(_00535_),
    .C(_00533_),
    .X(_00537_));
 sky130_fd_sc_hd__nor2_1 _08974_ (.A(_00536_),
    .B(_00537_),
    .Y(_00538_));
 sky130_fd_sc_hd__o2bb2ai_1 _08975_ (.A1_N(_00522_),
    .A2_N(_00523_),
    .B1(_00536_),
    .B2(_00537_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand3_1 _08976_ (.A(_00522_),
    .B(_00523_),
    .C(_00538_),
    .Y(_00541_));
 sky130_fd_sc_hd__and2_1 _08977_ (.A(_00539_),
    .B(_00541_),
    .X(_00542_));
 sky130_fd_sc_hd__a21o_1 _08978_ (.A1(_00539_),
    .A2(_00541_),
    .B1(_00483_),
    .X(_00543_));
 sky130_fd_sc_hd__nand3_1 _08979_ (.A(_00483_),
    .B(_00539_),
    .C(_00541_),
    .Y(_00544_));
 sky130_fd_sc_hd__and2_1 _08980_ (.A(_00543_),
    .B(_00544_),
    .X(_00545_));
 sky130_fd_sc_hd__o211ai_1 _08981_ (.A1(_00325_),
    .A2(_00378_),
    .B1(_00226_),
    .C1(_00324_),
    .Y(_00546_));
 sky130_fd_sc_hd__o21ai_1 _08982_ (.A1(_00326_),
    .A2(_00377_),
    .B1(_00546_),
    .Y(_00547_));
 sky130_fd_sc_hd__xor2_2 _08983_ (.A(_00545_),
    .B(_00547_),
    .X(_00548_));
 sky130_fd_sc_hd__a21oi_2 _08984_ (.A1(_00480_),
    .A2(_00482_),
    .B1(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__and3_2 _08985_ (.A(_00480_),
    .B(_00482_),
    .C(_00548_),
    .X(_00550_));
 sky130_fd_sc_hd__o211ai_4 _08986_ (.A1(_00549_),
    .A2(_00550_),
    .B1(_00322_),
    .C1(_00402_),
    .Y(_00552_));
 sky130_fd_sc_hd__a21o_2 _08987_ (.A1(_00322_),
    .A2(_00402_),
    .B1(_00549_),
    .X(_00553_));
 sky130_fd_sc_hd__o21ai_1 _08988_ (.A1(_00550_),
    .A2(_00553_),
    .B1(_00552_),
    .Y(_00554_));
 sky130_fd_sc_hd__o211ai_1 _08989_ (.A1(_00238_),
    .A2(_00239_),
    .B1(_00391_),
    .C1(_00393_),
    .Y(_00555_));
 sky130_fd_sc_hd__o211ai_2 _08990_ (.A1(_00237_),
    .A2(_00240_),
    .B1(_00390_),
    .C1(_00392_),
    .Y(_00556_));
 sky130_fd_sc_hd__a32o_1 _08991_ (.A1(_00247_),
    .A2(_00384_),
    .A3(_00385_),
    .B1(_00391_),
    .B2(_00394_),
    .X(_00557_));
 sky130_fd_sc_hd__xor2_1 _08992_ (.A(_00554_),
    .B(_00557_),
    .X(_00558_));
 sky130_fd_sc_hd__and3_1 _08993_ (.A(_00845_),
    .B(_00401_),
    .C(_00558_),
    .X(_00559_));
 sky130_fd_sc_hd__a21oi_1 _08994_ (.A1(_00845_),
    .A2(_00401_),
    .B1(_00558_),
    .Y(_00560_));
 sky130_fd_sc_hd__nor2_1 _08995_ (.A(_00559_),
    .B(_00560_),
    .Y(net71));
 sky130_fd_sc_hd__or4b_2 _08996_ (.A(_00395_),
    .B(_00396_),
    .C(_00558_),
    .D_N(_00246_),
    .X(_00562_));
 sky130_fd_sc_hd__nor2_1 _08997_ (.A(net6),
    .B(net7),
    .Y(_00563_));
 sky130_fd_sc_hd__nor3_4 _08998_ (.A(_00525_),
    .B(net7),
    .C(_00185_),
    .Y(_00564_));
 sky130_fd_sc_hd__o211ai_4 _08999_ (.A1(net7),
    .A2(_00526_),
    .B1(net8),
    .C1(net174),
    .Y(_00565_));
 sky130_fd_sc_hd__o21ai_4 _09000_ (.A1(_00321_),
    .A2(_00564_),
    .B1(_00594_),
    .Y(_00566_));
 sky130_fd_sc_hd__o21ai_4 _09001_ (.A1(_00321_),
    .A2(_00564_),
    .B1(net8),
    .Y(_00567_));
 sky130_fd_sc_hd__o211ai_4 _09002_ (.A1(net7),
    .A2(_00526_),
    .B1(_00594_),
    .C1(net174),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_8 _09003_ (.A(_00567_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_8 _09004_ (.A(net147),
    .B(net146),
    .Y(_00570_));
 sky130_fd_sc_hd__a21o_4 _09005_ (.A1(_00567_),
    .A2(_00568_),
    .B1(_00310_),
    .X(_00571_));
 sky130_fd_sc_hd__nor2_4 _09006_ (.A(net38),
    .B(net39),
    .Y(_00573_));
 sky130_fd_sc_hd__or2_2 _09007_ (.A(net38),
    .B(net39),
    .X(_00574_));
 sky130_fd_sc_hd__nand4_4 _09008_ (.A(_07504_),
    .B(_00140_),
    .C(_00573_),
    .D(_00551_),
    .Y(_00575_));
 sky130_fd_sc_hd__a21oi_4 _09009_ (.A1(_00575_),
    .A2(net57),
    .B1(net40),
    .Y(_00576_));
 sky130_fd_sc_hd__a21o_4 _09010_ (.A1(_00575_),
    .A2(net57),
    .B1(net40),
    .X(_00577_));
 sky130_fd_sc_hd__o311a_4 _09011_ (.A1(_00574_),
    .A2(net37),
    .A3(_00143_),
    .B1(net40),
    .C1(net57),
    .X(_00578_));
 sky130_fd_sc_hd__o211ai_4 _09012_ (.A1(_00263_),
    .A2(_00574_),
    .B1(net57),
    .C1(net40),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_8 _09013_ (.A(_00577_),
    .B(_00579_),
    .Y(_00580_));
 sky130_fd_sc_hd__nor2_8 _09014_ (.A(_00576_),
    .B(_00578_),
    .Y(_00581_));
 sky130_fd_sc_hd__or3_4 _09015_ (.A(_00288_),
    .B(_00576_),
    .C(_00578_),
    .X(_00582_));
 sky130_fd_sc_hd__a21bo_4 _09016_ (.A1(_00482_),
    .A2(_00548_),
    .B1_N(_00480_),
    .X(_00584_));
 sky130_fd_sc_hd__inv_2 _09017_ (.A(_00584_),
    .Y(_00585_));
 sky130_fd_sc_hd__a21boi_2 _09018_ (.A1(_00523_),
    .A2(_00538_),
    .B1_N(_00522_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand4_1 _09019_ (.A(_00528_),
    .B(_00531_),
    .C(_00534_),
    .D(net33),
    .Y(_00587_));
 sky130_fd_sc_hd__o31ai_2 _09020_ (.A1(_01292_),
    .A2(_00355_),
    .A3(_00366_),
    .B1(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _09021_ (.A(_00511_),
    .B(_00337_),
    .Y(_00589_));
 sky130_fd_sc_hd__a21oi_1 _09022_ (.A1(_00511_),
    .A2(_00513_),
    .B1(_00588_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand3b_1 _09023_ (.A_N(_00588_),
    .B(_00589_),
    .C(_00512_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand3_2 _09024_ (.A(_00511_),
    .B(_00513_),
    .C(_00588_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _09025_ (.A(_00591_),
    .B(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__o221a_1 _09026_ (.A1(_02790_),
    .A2(net163),
    .B1(_07537_),
    .B2(_00321_),
    .C1(_07536_),
    .X(_00595_));
 sky130_fd_sc_hd__a2bb2oi_1 _09027_ (.A1_N(_04638_),
    .A2_N(_04649_),
    .B1(_07438_),
    .B2(_07439_),
    .Y(_00596_));
 sky130_fd_sc_hd__o2111ai_4 _09028_ (.A1(_04606_),
    .A2(_04660_),
    .B1(_04704_),
    .C1(net162),
    .D1(_07437_),
    .Y(_00597_));
 sky130_fd_sc_hd__and3_1 _09029_ (.A(net156),
    .B(_07436_),
    .C(net154),
    .X(_00598_));
 sky130_fd_sc_hd__o211ai_4 _09030_ (.A1(_03435_),
    .A2(_03457_),
    .B1(net162),
    .C1(_07437_),
    .Y(_00599_));
 sky130_fd_sc_hd__nor2_2 _09031_ (.A(_00503_),
    .B(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__o31a_1 _09032_ (.A1(_04715_),
    .A2(_07146_),
    .A3(_07168_),
    .B1(_00599_),
    .X(_00601_));
 sky130_fd_sc_hd__o21ai_4 _09033_ (.A1(_04715_),
    .A2(_07189_),
    .B1(_00599_),
    .Y(_00602_));
 sky130_fd_sc_hd__o22ai_2 _09034_ (.A1(net159),
    .A2(net150),
    .B1(_00600_),
    .B2(_00601_),
    .Y(_00603_));
 sky130_fd_sc_hd__o2111ai_4 _09035_ (.A1(_00336_),
    .A2(_00597_),
    .B1(_00602_),
    .C1(_07540_),
    .D1(_02866_),
    .Y(_00604_));
 sky130_fd_sc_hd__o21ai_1 _09036_ (.A1(_00600_),
    .A2(_00601_),
    .B1(_00595_),
    .Y(_00606_));
 sky130_fd_sc_hd__o221ai_4 _09037_ (.A1(net159),
    .A2(net150),
    .B1(_00336_),
    .B2(_00597_),
    .C1(_00602_),
    .Y(_00607_));
 sky130_fd_sc_hd__o211ai_1 _09038_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_00189_),
    .C1(_00191_),
    .Y(_00608_));
 sky130_fd_sc_hd__or4_2 _09039_ (.A(_02079_),
    .B(_02100_),
    .C(_00188_),
    .D(_00190_),
    .X(_00609_));
 sky130_fd_sc_hd__o2111ai_1 _09040_ (.A1(_00066_),
    .A2(net160),
    .B1(_01631_),
    .C1(_00189_),
    .D1(_00495_),
    .Y(_00610_));
 sky130_fd_sc_hd__or4_1 _09041_ (.A(_01620_),
    .B(_00188_),
    .C(_00190_),
    .D(_00497_),
    .X(_00611_));
 sky130_fd_sc_hd__o2bb2ai_2 _09042_ (.A1_N(_00497_),
    .A2_N(_00608_),
    .B1(_00190_),
    .B2(_00610_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand3b_4 _09043_ (.A_N(_00612_),
    .B(_00604_),
    .C(_00603_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand3_4 _09044_ (.A(_00606_),
    .B(_00607_),
    .C(_00612_),
    .Y(_00614_));
 sky130_fd_sc_hd__o32a_1 _09045_ (.A1(_04715_),
    .A2(_05327_),
    .A3(_00336_),
    .B1(_07441_),
    .B2(net159),
    .X(_00615_));
 sky130_fd_sc_hd__a31o_1 _09046_ (.A1(_02866_),
    .A2(_00502_),
    .A3(_07440_),
    .B1(_00504_),
    .X(_00617_));
 sky130_fd_sc_hd__o211ai_2 _09047_ (.A1(_00501_),
    .A2(_00615_),
    .B1(_00614_),
    .C1(_00613_),
    .Y(_00618_));
 sky130_fd_sc_hd__a21bo_1 _09048_ (.A1(_00613_),
    .A2(_00614_),
    .B1_N(_00617_),
    .X(_00619_));
 sky130_fd_sc_hd__o2111ai_2 _09049_ (.A1(_00500_),
    .A2(_00504_),
    .B1(_00613_),
    .C1(_00614_),
    .D1(_00502_),
    .Y(_00620_));
 sky130_fd_sc_hd__a21o_1 _09050_ (.A1(_00613_),
    .A2(_00614_),
    .B1(_00617_),
    .X(_00621_));
 sky130_fd_sc_hd__nand2_1 _09051_ (.A(_00620_),
    .B(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _09052_ (.A(_00618_),
    .B(_00619_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _09053_ (.A(_00593_),
    .B(_00622_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand4_1 _09054_ (.A(_00591_),
    .B(_00592_),
    .C(_00620_),
    .D(_00621_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand4_1 _09055_ (.A(_00591_),
    .B(_00592_),
    .C(_00618_),
    .D(_00619_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _09056_ (.A(_00593_),
    .B(_00623_),
    .Y(_00628_));
 sky130_fd_sc_hd__a31oi_1 _09057_ (.A1(_00490_),
    .A2(_00515_),
    .A3(_00516_),
    .B1(_00491_),
    .Y(_00629_));
 sky130_fd_sc_hd__a31o_1 _09058_ (.A1(_00490_),
    .A2(_00515_),
    .A3(_00516_),
    .B1(_00491_),
    .X(_00630_));
 sky130_fd_sc_hd__nand3_2 _09059_ (.A(_00624_),
    .B(_00625_),
    .C(_00630_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand3_2 _09060_ (.A(_00626_),
    .B(_00628_),
    .C(_00629_),
    .Y(_00632_));
 sky130_fd_sc_hd__and3_1 _09061_ (.A(_00911_),
    .B(_00528_),
    .C(_00531_),
    .X(_00633_));
 sky130_fd_sc_hd__o22ai_4 _09062_ (.A1(_00333_),
    .A2(_00497_),
    .B1(_00366_),
    .B2(_01292_),
    .Y(_00634_));
 sky130_fd_sc_hd__or4_2 _09063_ (.A(_01292_),
    .B(_00333_),
    .C(_00497_),
    .D(_00366_),
    .X(_00635_));
 sky130_fd_sc_hd__a21oi_1 _09064_ (.A1(_00634_),
    .A2(_00635_),
    .B1(_00633_),
    .Y(_00636_));
 sky130_fd_sc_hd__and3_1 _09065_ (.A(_00635_),
    .B(_00633_),
    .C(_00634_),
    .X(_00637_));
 sky130_fd_sc_hd__a221oi_2 _09066_ (.A1(_00867_),
    .A2(_00889_),
    .B1(_00634_),
    .B2(_00635_),
    .C1(_00532_),
    .Y(_00639_));
 sky130_fd_sc_hd__o211a_1 _09067_ (.A1(_00900_),
    .A2(_00532_),
    .B1(_00634_),
    .C1(_00635_),
    .X(_00640_));
 sky130_fd_sc_hd__nor2_1 _09068_ (.A(_00636_),
    .B(_00637_),
    .Y(_00641_));
 sky130_fd_sc_hd__o211ai_1 _09069_ (.A1(_00636_),
    .A2(_00637_),
    .B1(_00631_),
    .C1(_00632_),
    .Y(_00642_));
 sky130_fd_sc_hd__o2bb2ai_1 _09070_ (.A1_N(_00631_),
    .A2_N(_00632_),
    .B1(_00639_),
    .B2(_00640_),
    .Y(_00643_));
 sky130_fd_sc_hd__a211o_1 _09071_ (.A1(_00631_),
    .A2(_00632_),
    .B1(_00639_),
    .C1(_00640_),
    .X(_00644_));
 sky130_fd_sc_hd__and2_1 _09072_ (.A(_00642_),
    .B(_00643_),
    .X(_00645_));
 sky130_fd_sc_hd__a31oi_2 _09073_ (.A1(_00631_),
    .A2(_00632_),
    .A3(_00641_),
    .B1(_00586_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand3_1 _09074_ (.A(_00586_),
    .B(_00642_),
    .C(_00643_),
    .Y(_00647_));
 sky130_fd_sc_hd__a21boi_2 _09075_ (.A1(_00646_),
    .A2(_00644_),
    .B1_N(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__o211ai_1 _09076_ (.A1(_00326_),
    .A2(_00377_),
    .B1(_00544_),
    .C1(_00546_),
    .Y(_00650_));
 sky130_fd_sc_hd__o21a_2 _09077_ (.A1(_00483_),
    .A2(_00542_),
    .B1(_00650_),
    .X(_00651_));
 sky130_fd_sc_hd__xnor2_4 _09078_ (.A(_00648_),
    .B(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__a21bo_1 _09079_ (.A1(_00456_),
    .A2(_00462_),
    .B1_N(_00457_),
    .X(_00653_));
 sky130_fd_sc_hd__o311a_1 _09080_ (.A1(_00284_),
    .A2(_00404_),
    .A3(_00405_),
    .B1(_00447_),
    .C1(_00448_),
    .X(_00654_));
 sky130_fd_sc_hd__o21bai_1 _09081_ (.A1(_00407_),
    .A2(_00449_),
    .B1_N(_00409_),
    .Y(_00655_));
 sky130_fd_sc_hd__a31o_1 _09082_ (.A1(_04255_),
    .A2(_05436_),
    .A3(_00460_),
    .B1(_00459_),
    .X(_00656_));
 sky130_fd_sc_hd__inv_2 _09083_ (.A(_00656_),
    .Y(_00657_));
 sky130_fd_sc_hd__o21ai_1 _09084_ (.A1(_00270_),
    .A2(_00280_),
    .B1(_00444_),
    .Y(_00658_));
 sky130_fd_sc_hd__a211oi_1 _09085_ (.A1(_00281_),
    .A2(_00444_),
    .B1(_00657_),
    .C1(_00440_),
    .Y(_00659_));
 sky130_fd_sc_hd__a211o_1 _09086_ (.A1(_00281_),
    .A2(_00444_),
    .B1(_00657_),
    .C1(_00440_),
    .X(_00661_));
 sky130_fd_sc_hd__a21oi_1 _09087_ (.A1(_00442_),
    .A2(_00658_),
    .B1(_00656_),
    .Y(_00662_));
 sky130_fd_sc_hd__a21o_1 _09088_ (.A1(_00442_),
    .A2(_00658_),
    .B1(_00656_),
    .X(_00663_));
 sky130_fd_sc_hd__or3_1 _09089_ (.A(_02636_),
    .B(_00005_),
    .C(_00007_),
    .X(_00664_));
 sky130_fd_sc_hd__or3_1 _09090_ (.A(_02636_),
    .B(_07508_),
    .C(_07510_),
    .X(_00665_));
 sky130_fd_sc_hd__and4_1 _09091_ (.A(_01969_),
    .B(_02647_),
    .C(_07513_),
    .D(_00010_),
    .X(_00666_));
 sky130_fd_sc_hd__or4_2 _09092_ (.A(_02636_),
    .B(_00005_),
    .C(_00007_),
    .D(_00411_),
    .X(_00667_));
 sky130_fd_sc_hd__o22ai_1 _09093_ (.A1(_02636_),
    .A2(_07512_),
    .B1(_00009_),
    .B2(_01958_),
    .Y(_00668_));
 sky130_fd_sc_hd__o31a_1 _09094_ (.A1(_02636_),
    .A2(_00009_),
    .A3(_00411_),
    .B1(_00668_),
    .X(_00669_));
 sky130_fd_sc_hd__o21a_1 _09095_ (.A1(net38),
    .A2(_00264_),
    .B1(net164),
    .X(_00670_));
 sky130_fd_sc_hd__o2bb2ai_4 _09096_ (.A1_N(_00273_),
    .A2_N(_00670_),
    .B1(_00426_),
    .B2(_00431_),
    .Y(_00672_));
 sky130_fd_sc_hd__o2111ai_4 _09097_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01172_),
    .C1(_00425_),
    .D1(_00427_),
    .Y(_00673_));
 sky130_fd_sc_hd__o21ai_1 _09098_ (.A1(_00433_),
    .A2(_00673_),
    .B1(_00672_),
    .Y(_00674_));
 sky130_fd_sc_hd__o221a_1 _09099_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_00142_),
    .B2(_00144_),
    .C1(_00148_),
    .X(_00675_));
 sky130_fd_sc_hd__o21ai_1 _09100_ (.A1(_01488_),
    .A2(net143),
    .B1(_00674_),
    .Y(_00676_));
 sky130_fd_sc_hd__o2111ai_4 _09101_ (.A1(_00433_),
    .A2(_00673_),
    .B1(_00672_),
    .C1(_01499_),
    .D1(_00150_),
    .Y(_00677_));
 sky130_fd_sc_hd__o221ai_4 _09102_ (.A1(_01488_),
    .A2(net143),
    .B1(_00433_),
    .B2(_00673_),
    .C1(_00672_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand2_1 _09103_ (.A(_00674_),
    .B(_00675_),
    .Y(_00679_));
 sky130_fd_sc_hd__nand3b_4 _09104_ (.A_N(_00669_),
    .B(_00678_),
    .C(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand3_4 _09105_ (.A(_00676_),
    .B(_00677_),
    .C(_00669_),
    .Y(_00681_));
 sky130_fd_sc_hd__a31o_1 _09106_ (.A1(_00148_),
    .A2(_00437_),
    .A3(_00417_),
    .B1(_00434_),
    .X(_00683_));
 sky130_fd_sc_hd__a21oi_1 _09107_ (.A1(_00680_),
    .A2(_00681_),
    .B1(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__and3_1 _09108_ (.A(_00680_),
    .B(_00681_),
    .C(_00683_),
    .X(_00685_));
 sky130_fd_sc_hd__nand3b_1 _09109_ (.A_N(_00683_),
    .B(_00681_),
    .C(_00680_),
    .Y(_00686_));
 sky130_fd_sc_hd__a21bo_1 _09110_ (.A1(_00680_),
    .A2(_00681_),
    .B1_N(_00683_),
    .X(_00687_));
 sky130_fd_sc_hd__nand2_1 _09111_ (.A(_00686_),
    .B(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__o211ai_2 _09112_ (.A1(_00684_),
    .A2(_00685_),
    .B1(_00661_),
    .C1(_00663_),
    .Y(_00689_));
 sky130_fd_sc_hd__o21ai_1 _09113_ (.A1(_00659_),
    .A2(_00662_),
    .B1(_00688_),
    .Y(_00690_));
 sky130_fd_sc_hd__nand3_1 _09114_ (.A(_00688_),
    .B(_00663_),
    .C(_00661_),
    .Y(_00691_));
 sky130_fd_sc_hd__o22ai_1 _09115_ (.A1(_00659_),
    .A2(_00662_),
    .B1(_00684_),
    .B2(_00685_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand3_1 _09116_ (.A(_00655_),
    .B(_00691_),
    .C(_00692_),
    .Y(_00694_));
 sky130_fd_sc_hd__o211ai_4 _09117_ (.A1(_00407_),
    .A2(_00654_),
    .B1(_00689_),
    .C1(_00690_),
    .Y(_00695_));
 sky130_fd_sc_hd__o21ai_2 _09118_ (.A1(_06265_),
    .A2(_06287_),
    .B1(_04255_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand3b_2 _09119_ (.A_N(_00412_),
    .B(_07370_),
    .C(_03917_),
    .Y(_00697_));
 sky130_fd_sc_hd__o32a_1 _09120_ (.A1(_01488_),
    .A2(_00411_),
    .A3(_00009_),
    .B1(net153),
    .B2(_03906_),
    .X(_00698_));
 sky130_fd_sc_hd__a32o_1 _09121_ (.A1(_00260_),
    .A2(_00010_),
    .A3(_01969_),
    .B1(_07370_),
    .B2(_03917_),
    .X(_00699_));
 sky130_fd_sc_hd__and3_1 _09122_ (.A(_00696_),
    .B(_00697_),
    .C(_00699_),
    .X(_00700_));
 sky130_fd_sc_hd__a21oi_1 _09123_ (.A1(_00697_),
    .A2(_00699_),
    .B1(_00696_),
    .Y(_00701_));
 sky130_fd_sc_hd__nor2_1 _09124_ (.A(_00700_),
    .B(_00701_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand3_1 _09125_ (.A(_00694_),
    .B(_00695_),
    .C(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__a21o_1 _09126_ (.A1(_00694_),
    .A2(_00695_),
    .B1(_00702_),
    .X(_00705_));
 sky130_fd_sc_hd__a21bo_1 _09127_ (.A1(_00694_),
    .A2(_00695_),
    .B1_N(_00702_),
    .X(_00706_));
 sky130_fd_sc_hd__o211ai_1 _09128_ (.A1(_00700_),
    .A2(_00701_),
    .B1(_00694_),
    .C1(_00695_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand3b_4 _09129_ (.A_N(_00653_),
    .B(_00703_),
    .C(_00705_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand3_2 _09130_ (.A(_00706_),
    .B(_00707_),
    .C(_00653_),
    .Y(_00709_));
 sky130_fd_sc_hd__o211ai_4 _09131_ (.A1(_00301_),
    .A2(_00303_),
    .B1(_00469_),
    .C1(_00472_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand4_2 _09132_ (.A(_00470_),
    .B(_00708_),
    .C(_00709_),
    .D(_00710_),
    .Y(_00711_));
 sky130_fd_sc_hd__a22o_1 _09133_ (.A1(_00708_),
    .A2(_00709_),
    .B1(_00710_),
    .B2(_00470_),
    .X(_00712_));
 sky130_fd_sc_hd__o2111ai_2 _09134_ (.A1(_05359_),
    .A2(_05370_),
    .B1(_05316_),
    .C1(_00711_),
    .D1(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__o2bb2a_1 _09135_ (.A1_N(_00711_),
    .A2_N(_00712_),
    .B1(_05327_),
    .B2(_05425_),
    .X(_00714_));
 sky130_fd_sc_hd__a32o_1 _09136_ (.A1(_05316_),
    .A2(_05392_),
    .A3(_05414_),
    .B1(_00711_),
    .B2(_00712_),
    .X(_00716_));
 sky130_fd_sc_hd__nand2_2 _09137_ (.A(_00713_),
    .B(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__xnor2_2 _09138_ (.A(_00652_),
    .B(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__xor2_4 _09139_ (.A(_00652_),
    .B(_00717_),
    .X(_00719_));
 sky130_fd_sc_hd__nand2_1 _09140_ (.A(_00585_),
    .B(_00718_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand2_2 _09141_ (.A(_00719_),
    .B(_00584_),
    .Y(_00721_));
 sky130_fd_sc_hd__nand2_1 _09142_ (.A(_00720_),
    .B(_00721_),
    .Y(_00722_));
 sky130_fd_sc_hd__o211ai_2 _09143_ (.A1(_00248_),
    .A2(_00389_),
    .B1(_00552_),
    .C1(_00555_),
    .Y(_00723_));
 sky130_fd_sc_hd__o211ai_4 _09144_ (.A1(_00553_),
    .A2(_00550_),
    .B1(_00391_),
    .C1(_00556_),
    .Y(_00724_));
 sky130_fd_sc_hd__a21o_1 _09145_ (.A1(_00552_),
    .A2(_00724_),
    .B1(_00722_),
    .X(_00725_));
 sky130_fd_sc_hd__nand3_1 _09146_ (.A(_00552_),
    .B(_00722_),
    .C(_00724_),
    .Y(_00727_));
 sky130_fd_sc_hd__and2_1 _09147_ (.A(_00725_),
    .B(_00727_),
    .X(_00728_));
 sky130_fd_sc_hd__xnor2_2 _09148_ (.A(_00582_),
    .B(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__xor2_4 _09149_ (.A(_00571_),
    .B(_00729_),
    .X(_00730_));
 sky130_fd_sc_hd__o221a_1 _09150_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_00401_),
    .B2(_00558_),
    .C1(_00730_),
    .X(_00731_));
 sky130_fd_sc_hd__a21oi_1 _09151_ (.A1(_00845_),
    .A2(_00562_),
    .B1(_00730_),
    .Y(_00732_));
 sky130_fd_sc_hd__nor2_1 _09152_ (.A(_00731_),
    .B(_00732_),
    .Y(net72));
 sky130_fd_sc_hd__o21ai_1 _09153_ (.A1(_00562_),
    .A2(_00730_),
    .B1(_00845_),
    .Y(_00733_));
 sky130_fd_sc_hd__a31o_1 _09154_ (.A1(_00582_),
    .A2(_00725_),
    .A3(_00727_),
    .B1(_00571_),
    .X(_00734_));
 sky130_fd_sc_hd__o21ai_2 _09155_ (.A1(_00582_),
    .A2(_00728_),
    .B1(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__nor4_1 _09156_ (.A(net37),
    .B(_00141_),
    .C(net40),
    .D(_07505_),
    .Y(_00737_));
 sky130_fd_sc_hd__nor3_4 _09157_ (.A(_00574_),
    .B(net40),
    .C(_00263_),
    .Y(_00738_));
 sky130_fd_sc_hd__o211ai_4 _09158_ (.A1(net40),
    .A2(_00575_),
    .B1(net41),
    .C1(net173),
    .Y(_00739_));
 sky130_fd_sc_hd__o21bai_4 _09159_ (.A1(_00299_),
    .A2(_00738_),
    .B1_N(net41),
    .Y(_00740_));
 sky130_fd_sc_hd__o21ai_4 _09160_ (.A1(_00299_),
    .A2(_00738_),
    .B1(net41),
    .Y(_00741_));
 sky130_fd_sc_hd__a311o_4 _09161_ (.A1(_00737_),
    .A2(_00583_),
    .A3(_00572_),
    .B1(_00299_),
    .C1(net41),
    .X(_00742_));
 sky130_fd_sc_hd__nand2_8 _09162_ (.A(_00741_),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_8 _09163_ (.A(_00739_),
    .B(_00740_),
    .Y(_00744_));
 sky130_fd_sc_hd__and3_1 _09164_ (.A(_00998_),
    .B(_00739_),
    .C(_00740_),
    .X(_00745_));
 sky130_fd_sc_hd__a22o_2 _09165_ (.A1(_00932_),
    .A2(_00954_),
    .B1(_00741_),
    .B2(_00742_),
    .X(_00746_));
 sky130_fd_sc_hd__and3_1 _09166_ (.A(net1),
    .B(_00745_),
    .C(_00581_),
    .X(_00748_));
 sky130_fd_sc_hd__or4_4 _09167_ (.A(_00288_),
    .B(_00987_),
    .C(_00580_),
    .D(_00744_),
    .X(_00749_));
 sky130_fd_sc_hd__a32o_4 _09168_ (.A1(net1),
    .A2(_00739_),
    .A3(_00740_),
    .B1(_00998_),
    .B2(_00581_),
    .X(_00750_));
 sky130_fd_sc_hd__o21a_2 _09169_ (.A1(_00652_),
    .A2(_00714_),
    .B1(_00713_),
    .X(_00751_));
 sky130_fd_sc_hd__inv_2 _09170_ (.A(_00751_),
    .Y(_00752_));
 sky130_fd_sc_hd__o32a_1 _09171_ (.A1(_05381_),
    .A2(_05403_),
    .A3(_07189_),
    .B1(_06331_),
    .B2(_05327_),
    .X(_00753_));
 sky130_fd_sc_hd__or3_1 _09172_ (.A(_06331_),
    .B(_07146_),
    .C(_07168_),
    .X(_00754_));
 sky130_fd_sc_hd__and4_1 _09173_ (.A(_05436_),
    .B(_06341_),
    .C(_07200_),
    .D(_05316_),
    .X(_00755_));
 sky130_fd_sc_hd__nor2_1 _09174_ (.A(_00753_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__a311o_1 _09175_ (.A1(_00655_),
    .A2(_00691_),
    .A3(_00692_),
    .B1(_00700_),
    .C1(_00701_),
    .X(_00757_));
 sky130_fd_sc_hd__nand2_1 _09176_ (.A(_00695_),
    .B(_00757_),
    .Y(_00759_));
 sky130_fd_sc_hd__and2_1 _09177_ (.A(_00695_),
    .B(_00757_),
    .X(_00760_));
 sky130_fd_sc_hd__a31oi_1 _09178_ (.A1(_00661_),
    .A2(_00686_),
    .A3(_00687_),
    .B1(_00662_),
    .Y(_00761_));
 sky130_fd_sc_hd__a31o_1 _09179_ (.A1(_00661_),
    .A2(_00686_),
    .A3(_00687_),
    .B1(_00662_),
    .X(_00762_));
 sky130_fd_sc_hd__o21ai_1 _09180_ (.A1(_04244_),
    .A2(_06331_),
    .B1(_00697_),
    .Y(_00763_));
 sky130_fd_sc_hd__o311ai_4 _09181_ (.A1(net165),
    .A2(net143),
    .A3(_00436_),
    .B1(_00681_),
    .C1(_00435_),
    .Y(_00764_));
 sky130_fd_sc_hd__nand2_1 _09182_ (.A(_00680_),
    .B(_00683_),
    .Y(_00765_));
 sky130_fd_sc_hd__o2111a_1 _09183_ (.A1(_00698_),
    .A2(_00696_),
    .B1(_00681_),
    .C1(_00697_),
    .D1(_00765_),
    .X(_00766_));
 sky130_fd_sc_hd__o2111ai_4 _09184_ (.A1(_00698_),
    .A2(_00696_),
    .B1(_00681_),
    .C1(_00697_),
    .D1(_00765_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand4_4 _09185_ (.A(_00680_),
    .B(_00699_),
    .C(_00763_),
    .D(_00764_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2_1 _09186_ (.A(_00672_),
    .B(_00675_),
    .Y(_00770_));
 sky130_fd_sc_hd__a41o_1 _09187_ (.A1(_00998_),
    .A2(net164),
    .A3(_00275_),
    .A4(_00429_),
    .B1(_00675_),
    .X(_00771_));
 sky130_fd_sc_hd__o21ai_1 _09188_ (.A1(_00433_),
    .A2(_00673_),
    .B1(_00770_),
    .Y(_00772_));
 sky130_fd_sc_hd__a31o_1 _09189_ (.A1(_00143_),
    .A2(net37),
    .A3(net57),
    .B1(_01958_),
    .X(_00773_));
 sky130_fd_sc_hd__o221a_1 _09190_ (.A1(_01892_),
    .A2(_01914_),
    .B1(_00142_),
    .B2(_00144_),
    .C1(_00148_),
    .X(_00774_));
 sky130_fd_sc_hd__o31ai_4 _09191_ (.A1(_01488_),
    .A2(_00270_),
    .A3(_00272_),
    .B1(_00673_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand4_4 _09192_ (.A(net164),
    .B(_01499_),
    .C(_00275_),
    .D(_00429_),
    .Y(_00776_));
 sky130_fd_sc_hd__o2bb2ai_4 _09193_ (.A1_N(_00775_),
    .A2_N(_00776_),
    .B1(_00147_),
    .B2(_00773_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand4_4 _09194_ (.A(_01969_),
    .B(_00150_),
    .C(_00775_),
    .D(_00776_),
    .Y(_00778_));
 sky130_fd_sc_hd__a21oi_2 _09195_ (.A1(_00777_),
    .A2(_00778_),
    .B1(_00772_),
    .Y(_00779_));
 sky130_fd_sc_hd__a22o_1 _09196_ (.A1(_00672_),
    .A2(_00771_),
    .B1(_00777_),
    .B2(_00778_),
    .X(_00781_));
 sky130_fd_sc_hd__and3_1 _09197_ (.A(_00772_),
    .B(_00777_),
    .C(_00778_),
    .X(_00782_));
 sky130_fd_sc_hd__nand4_4 _09198_ (.A(_00672_),
    .B(_00771_),
    .C(_00777_),
    .D(_00778_),
    .Y(_00783_));
 sky130_fd_sc_hd__nand3_1 _09199_ (.A(_00781_),
    .B(_00783_),
    .C(_00666_),
    .Y(_00784_));
 sky130_fd_sc_hd__o21ai_1 _09200_ (.A1(_00779_),
    .A2(_00782_),
    .B1(_00667_),
    .Y(_00785_));
 sky130_fd_sc_hd__o21ai_1 _09201_ (.A1(_00411_),
    .A2(_00664_),
    .B1(_00783_),
    .Y(_00786_));
 sky130_fd_sc_hd__o311a_1 _09202_ (.A1(_02636_),
    .A2(_00411_),
    .A3(_00009_),
    .B1(_00783_),
    .C1(_00781_),
    .X(_00787_));
 sky130_fd_sc_hd__a21oi_1 _09203_ (.A1(_00781_),
    .A2(_00783_),
    .B1(_00667_),
    .Y(_00788_));
 sky130_fd_sc_hd__o21ai_1 _09204_ (.A1(_00779_),
    .A2(_00782_),
    .B1(_00666_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand2_1 _09205_ (.A(_00784_),
    .B(_00785_),
    .Y(_00790_));
 sky130_fd_sc_hd__o2111ai_1 _09206_ (.A1(_00786_),
    .A2(_00779_),
    .B1(_00768_),
    .C1(_00767_),
    .D1(_00789_),
    .Y(_00792_));
 sky130_fd_sc_hd__o2bb2ai_1 _09207_ (.A1_N(_00767_),
    .A2_N(_00768_),
    .B1(_00787_),
    .B2(_00788_),
    .Y(_00793_));
 sky130_fd_sc_hd__a22o_1 _09208_ (.A1(_00767_),
    .A2(_00768_),
    .B1(_00784_),
    .B2(_00785_),
    .X(_00794_));
 sky130_fd_sc_hd__nand4_1 _09209_ (.A(_00767_),
    .B(_00768_),
    .C(_00784_),
    .D(_00785_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand3_1 _09210_ (.A(_00762_),
    .B(_00792_),
    .C(_00793_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand3_1 _09211_ (.A(_00794_),
    .B(_00795_),
    .C(_00761_),
    .Y(_00797_));
 sky130_fd_sc_hd__a32o_1 _09212_ (.A1(_02647_),
    .A2(_00006_),
    .A3(_00008_),
    .B1(_03917_),
    .B2(_07513_),
    .X(_00798_));
 sky130_fd_sc_hd__and4_1 _09213_ (.A(_02647_),
    .B(_03917_),
    .C(_07513_),
    .D(_00010_),
    .X(_00799_));
 sky130_fd_sc_hd__o31a_1 _09214_ (.A1(_03906_),
    .A2(_00009_),
    .A3(_00665_),
    .B1(_00798_),
    .X(_00800_));
 sky130_fd_sc_hd__a21oi_1 _09215_ (.A1(_04255_),
    .A2(_07370_),
    .B1(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__and3_1 _09216_ (.A(_00800_),
    .B(_07370_),
    .C(_04255_),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _09217_ (.A(_00801_),
    .B(_00802_),
    .X(_00803_));
 sky130_fd_sc_hd__a21o_1 _09218_ (.A1(_00796_),
    .A2(_00797_),
    .B1(_00803_),
    .X(_00804_));
 sky130_fd_sc_hd__nand3_1 _09219_ (.A(_00796_),
    .B(_00797_),
    .C(_00803_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand2_1 _09220_ (.A(_00804_),
    .B(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__and2_1 _09221_ (.A(_00804_),
    .B(_00805_),
    .X(_00807_));
 sky130_fd_sc_hd__a21o_1 _09222_ (.A1(_00695_),
    .A2(_00757_),
    .B1(_00806_),
    .X(_00808_));
 sky130_fd_sc_hd__a21o_1 _09223_ (.A1(_00804_),
    .A2(_00805_),
    .B1(_00759_),
    .X(_00809_));
 sky130_fd_sc_hd__nand3_2 _09224_ (.A(_00469_),
    .B(_00475_),
    .C(_00709_),
    .Y(_00810_));
 sky130_fd_sc_hd__nand3_1 _09225_ (.A(_00470_),
    .B(_00708_),
    .C(_00710_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand4_1 _09226_ (.A(_00708_),
    .B(_00808_),
    .C(_00809_),
    .D(_00810_),
    .Y(_00813_));
 sky130_fd_sc_hd__a22o_1 _09227_ (.A1(_00808_),
    .A2(_00809_),
    .B1(_00810_),
    .B2(_00708_),
    .X(_00814_));
 sky130_fd_sc_hd__and2_1 _09228_ (.A(_00813_),
    .B(_00814_),
    .X(_00815_));
 sky130_fd_sc_hd__a2bb2o_1 _09229_ (.A1_N(_00753_),
    .A2_N(_00755_),
    .B1(_00813_),
    .B2(_00814_),
    .X(_00816_));
 sky130_fd_sc_hd__nand3_1 _09230_ (.A(_00814_),
    .B(_00756_),
    .C(_00813_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_2 _09231_ (.A(_00816_),
    .B(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__a32o_1 _09232_ (.A1(_01631_),
    .A2(_00362_),
    .A3(_00364_),
    .B1(_02133_),
    .B2(_00193_),
    .X(_00819_));
 sky130_fd_sc_hd__o31a_1 _09233_ (.A1(_02210_),
    .A2(_00192_),
    .A3(_00366_),
    .B1(_00819_),
    .X(_00820_));
 sky130_fd_sc_hd__or3_2 _09234_ (.A(_01292_),
    .B(_00532_),
    .C(_00820_),
    .X(_00821_));
 sky130_fd_sc_hd__o21ai_2 _09235_ (.A1(_01292_),
    .A2(_00532_),
    .B1(_00820_),
    .Y(_00822_));
 sky130_fd_sc_hd__and2_1 _09236_ (.A(_00821_),
    .B(_00822_),
    .X(_00824_));
 sky130_fd_sc_hd__and3_1 _09237_ (.A(_00592_),
    .B(_00618_),
    .C(_00619_),
    .X(_00825_));
 sky130_fd_sc_hd__a21oi_1 _09238_ (.A1(_00622_),
    .A2(_00592_),
    .B1(_00590_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _09239_ (.A(_00633_),
    .B(_00634_),
    .Y(_00827_));
 sky130_fd_sc_hd__o41ai_1 _09240_ (.A1(_01292_),
    .A2(_00333_),
    .A3(_00366_),
    .A4(_00497_),
    .B1(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hd__o21ai_1 _09241_ (.A1(_00501_),
    .A2(_00615_),
    .B1(_00613_),
    .Y(_00829_));
 sky130_fd_sc_hd__nand2_1 _09242_ (.A(_00614_),
    .B(_00617_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand4_2 _09243_ (.A(_00613_),
    .B(_00635_),
    .C(_00827_),
    .D(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__and3_1 _09244_ (.A(_00828_),
    .B(_00829_),
    .C(_00614_),
    .X(_00832_));
 sky130_fd_sc_hd__nand3_1 _09245_ (.A(_00828_),
    .B(_00829_),
    .C(_00614_),
    .Y(_00833_));
 sky130_fd_sc_hd__o221ai_4 _09246_ (.A1(_02790_),
    .A2(net163),
    .B1(_00063_),
    .B2(_00066_),
    .C1(_00070_),
    .Y(_00835_));
 sky130_fd_sc_hd__o221ai_2 _09247_ (.A1(_03435_),
    .A2(_03457_),
    .B1(_07537_),
    .B2(_00321_),
    .C1(_07536_),
    .Y(_00836_));
 sky130_fd_sc_hd__a32oi_4 _09248_ (.A1(_03555_),
    .A2(_07536_),
    .A3(_07538_),
    .B1(_07440_),
    .B2(_04726_),
    .Y(_00837_));
 sky130_fd_sc_hd__o21ai_1 _09249_ (.A1(_04715_),
    .A2(_07441_),
    .B1(_00836_),
    .Y(_00838_));
 sky130_fd_sc_hd__nand4_2 _09250_ (.A(_00596_),
    .B(_07538_),
    .C(_07536_),
    .D(_03555_),
    .Y(_00839_));
 sky130_fd_sc_hd__o21ai_1 _09251_ (.A1(_03544_),
    .A2(net150),
    .B1(_00596_),
    .Y(_00840_));
 sky130_fd_sc_hd__nand4_2 _09252_ (.A(_03555_),
    .B(_07536_),
    .C(_07538_),
    .D(_00597_),
    .Y(_00841_));
 sky130_fd_sc_hd__o211ai_4 _09253_ (.A1(net159),
    .A2(net148),
    .B1(_00840_),
    .C1(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__nand4_4 _09254_ (.A(_02866_),
    .B(_00072_),
    .C(_00838_),
    .D(_00839_),
    .Y(_00843_));
 sky130_fd_sc_hd__o32a_1 _09255_ (.A1(net158),
    .A2(_07189_),
    .A3(_00597_),
    .B1(net150),
    .B2(net159),
    .X(_00844_));
 sky130_fd_sc_hd__a31o_1 _09256_ (.A1(_02866_),
    .A2(_07540_),
    .A3(_00602_),
    .B1(_00600_),
    .X(_00846_));
 sky130_fd_sc_hd__a21oi_1 _09257_ (.A1(_00842_),
    .A2(_00843_),
    .B1(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__o2bb2ai_2 _09258_ (.A1_N(_00842_),
    .A2_N(_00843_),
    .B1(_00844_),
    .B2(_00601_),
    .Y(_00848_));
 sky130_fd_sc_hd__o2111ai_4 _09259_ (.A1(_00595_),
    .A2(_00600_),
    .B1(_00602_),
    .C1(_00842_),
    .D1(_00843_),
    .Y(_00849_));
 sky130_fd_sc_hd__a2bb2o_1 _09260_ (.A1_N(_00493_),
    .A2_N(_00609_),
    .B1(_00848_),
    .B2(_00849_),
    .X(_00850_));
 sky130_fd_sc_hd__nand3b_1 _09261_ (.A_N(_00611_),
    .B(_00848_),
    .C(_00849_),
    .Y(_00851_));
 sky130_fd_sc_hd__a211o_1 _09262_ (.A1(_00848_),
    .A2(_00849_),
    .B1(_00493_),
    .C1(_00609_),
    .X(_00852_));
 sky130_fd_sc_hd__o211ai_2 _09263_ (.A1(_00493_),
    .A2(_00609_),
    .B1(_00848_),
    .C1(_00849_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_1 _09264_ (.A(_00852_),
    .B(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__a22o_1 _09265_ (.A1(_00831_),
    .A2(_00833_),
    .B1(_00852_),
    .B2(_00853_),
    .X(_00855_));
 sky130_fd_sc_hd__nand4_1 _09266_ (.A(_00831_),
    .B(_00833_),
    .C(_00852_),
    .D(_00853_),
    .Y(_00857_));
 sky130_fd_sc_hd__a22o_1 _09267_ (.A1(_00831_),
    .A2(_00833_),
    .B1(_00850_),
    .B2(_00851_),
    .X(_00858_));
 sky130_fd_sc_hd__nand4_1 _09268_ (.A(_00831_),
    .B(_00833_),
    .C(_00850_),
    .D(_00851_),
    .Y(_00859_));
 sky130_fd_sc_hd__o211a_1 _09269_ (.A1(_00590_),
    .A2(_00825_),
    .B1(_00855_),
    .C1(_00857_),
    .X(_00860_));
 sky130_fd_sc_hd__o211ai_1 _09270_ (.A1(_00590_),
    .A2(_00825_),
    .B1(_00855_),
    .C1(_00857_),
    .Y(_00861_));
 sky130_fd_sc_hd__nand3_1 _09271_ (.A(_00826_),
    .B(_00858_),
    .C(_00859_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(_00861_),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__a21oi_1 _09273_ (.A1(_00821_),
    .A2(_00822_),
    .B1(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__a21o_1 _09274_ (.A1(_00821_),
    .A2(_00822_),
    .B1(_00863_),
    .X(_00865_));
 sky130_fd_sc_hd__nand2_1 _09275_ (.A(_00824_),
    .B(_00863_),
    .Y(_00866_));
 sky130_fd_sc_hd__a31o_1 _09276_ (.A1(_00821_),
    .A2(_00822_),
    .A3(_00862_),
    .B1(_00860_),
    .X(_00868_));
 sky130_fd_sc_hd__a31oi_1 _09277_ (.A1(_00821_),
    .A2(_00822_),
    .A3(_00863_),
    .B1(_00864_),
    .Y(_00869_));
 sky130_fd_sc_hd__a21bo_1 _09278_ (.A1(_00632_),
    .A2(_00641_),
    .B1_N(_00631_),
    .X(_00870_));
 sky130_fd_sc_hd__nand3_1 _09279_ (.A(_00865_),
    .B(_00866_),
    .C(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hd__a21o_1 _09280_ (.A1(_00865_),
    .A2(_00866_),
    .B1(_00870_),
    .X(_00872_));
 sky130_fd_sc_hd__nand2_2 _09281_ (.A(_00871_),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__o211ai_1 _09282_ (.A1(_00483_),
    .A2(_00542_),
    .B1(_00647_),
    .C1(_00650_),
    .Y(_00874_));
 sky130_fd_sc_hd__a22o_1 _09283_ (.A1(_00644_),
    .A2(_00646_),
    .B1(_00651_),
    .B2(_00647_),
    .X(_00875_));
 sky130_fd_sc_hd__xor2_4 _09284_ (.A(_00873_),
    .B(_00875_),
    .X(_00876_));
 sky130_fd_sc_hd__xnor2_2 _09285_ (.A(_00818_),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__xor2_4 _09286_ (.A(_00818_),
    .B(_00876_),
    .X(_00879_));
 sky130_fd_sc_hd__nand2_2 _09287_ (.A(_00877_),
    .B(_00751_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_2 _09288_ (.A(_00879_),
    .B(_00752_),
    .Y(_00881_));
 sky130_fd_sc_hd__o211ai_4 _09289_ (.A1(_00550_),
    .A2(_00553_),
    .B1(_00721_),
    .C1(_00723_),
    .Y(_00882_));
 sky130_fd_sc_hd__o211ai_2 _09290_ (.A1(_00719_),
    .A2(_00584_),
    .B1(_00552_),
    .C1(_00724_),
    .Y(_00883_));
 sky130_fd_sc_hd__a22o_2 _09291_ (.A1(_00880_),
    .A2(_00881_),
    .B1(_00882_),
    .B2(_00720_),
    .X(_00884_));
 sky130_fd_sc_hd__o2111ai_4 _09292_ (.A1(_00584_),
    .A2(_00719_),
    .B1(_00880_),
    .C1(_00881_),
    .D1(_00882_),
    .Y(_00885_));
 sky130_fd_sc_hd__o2111a_1 _09293_ (.A1(_00582_),
    .A2(_00746_),
    .B1(_00750_),
    .C1(_00884_),
    .D1(_00885_),
    .X(_00886_));
 sky130_fd_sc_hd__o2111ai_4 _09294_ (.A1(_00582_),
    .A2(_00746_),
    .B1(_00750_),
    .C1(_00884_),
    .D1(_00885_),
    .Y(_00887_));
 sky130_fd_sc_hd__a22oi_4 _09295_ (.A1(_00749_),
    .A2(_00750_),
    .B1(_00884_),
    .B2(_00885_),
    .Y(_00888_));
 sky130_fd_sc_hd__nor2_2 _09296_ (.A(net7),
    .B(net8),
    .Y(_00890_));
 sky130_fd_sc_hd__or2_2 _09297_ (.A(net7),
    .B(net8),
    .X(_00891_));
 sky130_fd_sc_hd__nand4_4 _09298_ (.A(net160),
    .B(_00524_),
    .C(_00890_),
    .D(_00540_),
    .Y(_00892_));
 sky130_fd_sc_hd__a41oi_4 _09299_ (.A1(net160),
    .A2(_00524_),
    .A3(_00890_),
    .A4(_00540_),
    .B1(_00321_),
    .Y(_00893_));
 sky130_fd_sc_hd__o311a_2 _09300_ (.A1(_00185_),
    .A2(_00525_),
    .A3(_00891_),
    .B1(_00605_),
    .C1(net174),
    .X(_00894_));
 sky130_fd_sc_hd__nand2_2 _09301_ (.A(_00893_),
    .B(_00605_),
    .Y(_00895_));
 sky130_fd_sc_hd__a21oi_4 _09302_ (.A1(_00892_),
    .A2(net174),
    .B1(_00605_),
    .Y(_00896_));
 sky130_fd_sc_hd__a21o_1 _09303_ (.A1(_00892_),
    .A2(net174),
    .B1(_00605_),
    .X(_00897_));
 sky130_fd_sc_hd__o311a_4 _09304_ (.A1(_00185_),
    .A2(_00525_),
    .A3(_00891_),
    .B1(net9),
    .C1(net174),
    .X(_00898_));
 sky130_fd_sc_hd__nand2_8 _09305_ (.A(net9),
    .B(_00893_),
    .Y(_00899_));
 sky130_fd_sc_hd__a21oi_4 _09306_ (.A1(_00892_),
    .A2(net174),
    .B1(net9),
    .Y(_00901_));
 sky130_fd_sc_hd__a21o_4 _09307_ (.A1(_00892_),
    .A2(net174),
    .B1(net9),
    .X(_00902_));
 sky130_fd_sc_hd__nand2_8 _09308_ (.A(_00899_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand2_8 _09309_ (.A(_00895_),
    .B(_00897_),
    .Y(_00904_));
 sky130_fd_sc_hd__and3_1 _09310_ (.A(_00911_),
    .B(_00899_),
    .C(_00902_),
    .X(_00905_));
 sky130_fd_sc_hd__or4_4 _09311_ (.A(_00310_),
    .B(_00900_),
    .C(_00570_),
    .D(_00903_),
    .X(_00906_));
 sky130_fd_sc_hd__a32o_1 _09312_ (.A1(net33),
    .A2(_00899_),
    .A3(_00902_),
    .B1(_00569_),
    .B2(_00911_),
    .X(_00907_));
 sky130_fd_sc_hd__nand2_1 _09313_ (.A(_00906_),
    .B(_00907_),
    .Y(_00908_));
 sky130_fd_sc_hd__o21ai_2 _09314_ (.A1(_00886_),
    .A2(_00888_),
    .B1(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand3_2 _09315_ (.A(_00887_),
    .B(_00906_),
    .C(_00907_),
    .Y(_00910_));
 sky130_fd_sc_hd__o21ai_1 _09316_ (.A1(_00888_),
    .A2(_00910_),
    .B1(_00909_),
    .Y(_00912_));
 sky130_fd_sc_hd__o211ai_4 _09317_ (.A1(_00910_),
    .A2(_00888_),
    .B1(_00735_),
    .C1(_00909_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_1 _09318_ (.A(_00735_),
    .B(_00912_),
    .Y(_00914_));
 sky130_fd_sc_hd__xnor2_1 _09319_ (.A(_00733_),
    .B(_00914_),
    .Y(net73));
 sky130_fd_sc_hd__o32a_1 _09320_ (.A1(_00562_),
    .A2(_00730_),
    .A3(_00914_),
    .B1(_00823_),
    .B2(_00812_),
    .X(_00915_));
 sky130_fd_sc_hd__nand2_1 _09321_ (.A(_00817_),
    .B(_00876_),
    .Y(_00916_));
 sky130_fd_sc_hd__o21a_2 _09322_ (.A1(_00756_),
    .A2(_00815_),
    .B1(_00916_),
    .X(_00917_));
 sky130_fd_sc_hd__o21ai_2 _09323_ (.A1(_00756_),
    .A2(_00815_),
    .B1(_00916_),
    .Y(_00918_));
 sky130_fd_sc_hd__o32a_1 _09324_ (.A1(_06331_),
    .A2(_07146_),
    .A3(_07168_),
    .B1(net153),
    .B2(_05327_),
    .X(_00919_));
 sky130_fd_sc_hd__and4_1 _09325_ (.A(_06341_),
    .B(_07200_),
    .C(_07370_),
    .D(_05316_),
    .X(_00920_));
 sky130_fd_sc_hd__a2bb2o_1 _09326_ (.A1_N(_00919_),
    .A2_N(_00920_),
    .B1(_05436_),
    .B2(_07440_),
    .X(_00922_));
 sky130_fd_sc_hd__or4_1 _09327_ (.A(_05425_),
    .B(_00920_),
    .C(_07441_),
    .D(_00919_),
    .X(_00923_));
 sky130_fd_sc_hd__a21oi_1 _09328_ (.A1(_00922_),
    .A2(_00923_),
    .B1(_00755_),
    .Y(_00924_));
 sky130_fd_sc_hd__and3_1 _09329_ (.A(_00923_),
    .B(_00755_),
    .C(_00922_),
    .X(_00925_));
 sky130_fd_sc_hd__nor2_1 _09330_ (.A(_00924_),
    .B(_00925_),
    .Y(_00926_));
 sky130_fd_sc_hd__a31o_1 _09331_ (.A1(_04255_),
    .A2(_07370_),
    .A3(_00798_),
    .B1(_00799_),
    .X(_00927_));
 sky130_fd_sc_hd__inv_2 _09332_ (.A(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand3_1 _09333_ (.A(_00781_),
    .B(_00786_),
    .C(_00927_),
    .Y(_00929_));
 sky130_fd_sc_hd__and3_1 _09334_ (.A(_01969_),
    .B(_00271_),
    .C(_00273_),
    .X(_00930_));
 sky130_fd_sc_hd__or3_1 _09335_ (.A(_01958_),
    .B(_00270_),
    .C(_00272_),
    .X(_00931_));
 sky130_fd_sc_hd__and3_1 _09336_ (.A(_01499_),
    .B(_00425_),
    .C(_00427_),
    .X(_00933_));
 sky130_fd_sc_hd__a32o_1 _09337_ (.A1(net164),
    .A2(_00271_),
    .A3(_00273_),
    .B1(_00775_),
    .B2(_00774_),
    .X(_00934_));
 sky130_fd_sc_hd__nand2_1 _09338_ (.A(_00934_),
    .B(_00933_),
    .Y(_00935_));
 sky130_fd_sc_hd__a32o_1 _09339_ (.A1(_01499_),
    .A2(_00425_),
    .A3(_00427_),
    .B1(_00775_),
    .B2(_00774_),
    .X(_00936_));
 sky130_fd_sc_hd__nand2_1 _09340_ (.A(_00936_),
    .B(_00930_),
    .Y(_00937_));
 sky130_fd_sc_hd__a22oi_1 _09341_ (.A1(_00934_),
    .A2(_00933_),
    .B1(_00930_),
    .B2(_00936_),
    .Y(_00938_));
 sky130_fd_sc_hd__a31o_1 _09342_ (.A1(_01969_),
    .A2(_00271_),
    .A3(_00273_),
    .B1(_00936_),
    .X(_00939_));
 sky130_fd_sc_hd__a2bb2oi_1 _09343_ (.A1_N(_00931_),
    .A2_N(_00935_),
    .B1(_00939_),
    .B2(_00938_),
    .Y(_00940_));
 sky130_fd_sc_hd__o211a_1 _09344_ (.A1(_00667_),
    .A2(_00779_),
    .B1(_00783_),
    .C1(_00928_),
    .X(_00941_));
 sky130_fd_sc_hd__o211ai_1 _09345_ (.A1(_00667_),
    .A2(_00779_),
    .B1(_00783_),
    .C1(_00928_),
    .Y(_00942_));
 sky130_fd_sc_hd__o21a_1 _09346_ (.A1(_00940_),
    .A2(_00941_),
    .B1(_00929_),
    .X(_00944_));
 sky130_fd_sc_hd__nand3b_1 _09347_ (.A_N(_00940_),
    .B(_00942_),
    .C(_00929_),
    .Y(_00945_));
 sky130_fd_sc_hd__a21bo_1 _09348_ (.A1(_00929_),
    .A2(_00942_),
    .B1_N(_00940_),
    .X(_00946_));
 sky130_fd_sc_hd__o211a_1 _09349_ (.A1(_00786_),
    .A2(_00779_),
    .B1(_00768_),
    .C1(_00789_),
    .X(_00947_));
 sky130_fd_sc_hd__o21ai_1 _09350_ (.A1(_00766_),
    .A2(_00790_),
    .B1(_00768_),
    .Y(_00948_));
 sky130_fd_sc_hd__o2bb2ai_2 _09351_ (.A1_N(_00945_),
    .A2_N(_00946_),
    .B1(_00947_),
    .B2(_00766_),
    .Y(_00949_));
 sky130_fd_sc_hd__and3_1 _09352_ (.A(_00948_),
    .B(_00946_),
    .C(_00945_),
    .X(_00950_));
 sky130_fd_sc_hd__nand3_1 _09353_ (.A(_00948_),
    .B(_00946_),
    .C(_00945_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand2_1 _09354_ (.A(_00949_),
    .B(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__or3_2 _09355_ (.A(_04244_),
    .B(_07508_),
    .C(_07510_),
    .X(_00953_));
 sky130_fd_sc_hd__and3_1 _09356_ (.A(_03917_),
    .B(_00146_),
    .C(_00148_),
    .X(_00955_));
 sky130_fd_sc_hd__o32a_1 _09357_ (.A1(_02636_),
    .A2(_00145_),
    .A3(_00147_),
    .B1(_03906_),
    .B2(_00009_),
    .X(_00956_));
 sky130_fd_sc_hd__a31o_1 _09358_ (.A1(_02647_),
    .A2(_00010_),
    .A3(_00955_),
    .B1(_00956_),
    .X(_00957_));
 sky130_fd_sc_hd__xor2_2 _09359_ (.A(_00953_),
    .B(_00957_),
    .X(_00958_));
 sky130_fd_sc_hd__inv_2 _09360_ (.A(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__and3_2 _09361_ (.A(_00949_),
    .B(_00951_),
    .C(_00959_),
    .X(_00960_));
 sky130_fd_sc_hd__a21oi_1 _09362_ (.A1(_00949_),
    .A2(_00951_),
    .B1(_00959_),
    .Y(_00961_));
 sky130_fd_sc_hd__a21boi_2 _09363_ (.A1(_00797_),
    .A2(_00803_),
    .B1_N(_00796_),
    .Y(_00962_));
 sky130_fd_sc_hd__o21ai_4 _09364_ (.A1(_00960_),
    .A2(_00961_),
    .B1(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__a21o_1 _09365_ (.A1(_00952_),
    .A2(_00958_),
    .B1(_00962_),
    .X(_00964_));
 sky130_fd_sc_hd__a31o_1 _09366_ (.A1(_00949_),
    .A2(_00951_),
    .A3(_00959_),
    .B1(_00964_),
    .X(_00966_));
 sky130_fd_sc_hd__o21ai_1 _09367_ (.A1(_00960_),
    .A2(_00964_),
    .B1(_00963_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand3_2 _09368_ (.A(_00709_),
    .B(_00809_),
    .C(_00811_),
    .Y(_00968_));
 sky130_fd_sc_hd__o211ai_2 _09369_ (.A1(_00806_),
    .A2(_00760_),
    .B1(_00708_),
    .C1(_00810_),
    .Y(_00969_));
 sky130_fd_sc_hd__a22o_1 _09370_ (.A1(_00963_),
    .A2(_00966_),
    .B1(_00969_),
    .B2(_00809_),
    .X(_00970_));
 sky130_fd_sc_hd__a21o_1 _09371_ (.A1(_00808_),
    .A2(_00968_),
    .B1(_00967_),
    .X(_00971_));
 sky130_fd_sc_hd__a21o_1 _09372_ (.A1(_00809_),
    .A2(_00969_),
    .B1(_00967_),
    .X(_00972_));
 sky130_fd_sc_hd__a22o_1 _09373_ (.A1(_00963_),
    .A2(_00966_),
    .B1(_00968_),
    .B2(_00808_),
    .X(_00973_));
 sky130_fd_sc_hd__o211ai_1 _09374_ (.A1(_00924_),
    .A2(_00925_),
    .B1(_00970_),
    .C1(_00971_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand3_2 _09375_ (.A(_00973_),
    .B(_00926_),
    .C(_00972_),
    .Y(_00975_));
 sky130_fd_sc_hd__nand2_1 _09376_ (.A(_00974_),
    .B(_00975_),
    .Y(_00977_));
 sky130_fd_sc_hd__a32o_1 _09377_ (.A1(_00367_),
    .A2(_02199_),
    .A3(_00193_),
    .B1(_00533_),
    .B2(_01303_),
    .X(_00978_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(_00819_),
    .B(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__o21ai_1 _09379_ (.A1(_00493_),
    .A2(_00609_),
    .B1(_00849_),
    .Y(_00980_));
 sky130_fd_sc_hd__o211ai_2 _09380_ (.A1(_00611_),
    .A2(_00847_),
    .B1(_00849_),
    .C1(_00979_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand4_2 _09381_ (.A(_00819_),
    .B(_00848_),
    .C(_00978_),
    .D(_00980_),
    .Y(_00982_));
 sky130_fd_sc_hd__a21oi_2 _09382_ (.A1(_00597_),
    .A2(_00836_),
    .B1(_00835_),
    .Y(_00983_));
 sky130_fd_sc_hd__o221a_1 _09383_ (.A1(_04638_),
    .A2(_04649_),
    .B1(_07537_),
    .B2(_00321_),
    .C1(_07536_),
    .X(_00984_));
 sky130_fd_sc_hd__o22ai_4 _09384_ (.A1(_04715_),
    .A2(net150),
    .B1(_00835_),
    .B2(_00837_),
    .Y(_00985_));
 sky130_fd_sc_hd__o21ai_4 _09385_ (.A1(_00598_),
    .A2(_00983_),
    .B1(_00984_),
    .Y(_00986_));
 sky130_fd_sc_hd__a22oi_1 _09386_ (.A1(_03555_),
    .A2(_00072_),
    .B1(_00985_),
    .B2(_00986_),
    .Y(_00988_));
 sky130_fd_sc_hd__and4_1 _09387_ (.A(_03555_),
    .B(_00072_),
    .C(_00985_),
    .D(_00986_),
    .X(_00989_));
 sky130_fd_sc_hd__a211o_1 _09388_ (.A1(_00985_),
    .A2(_00986_),
    .B1(_03544_),
    .C1(net148),
    .X(_00990_));
 sky130_fd_sc_hd__o221ai_2 _09389_ (.A1(_03544_),
    .A2(net148),
    .B1(_00983_),
    .B2(_00984_),
    .C1(_00986_),
    .Y(_00991_));
 sky130_fd_sc_hd__nor2_1 _09390_ (.A(_00988_),
    .B(_00989_),
    .Y(_00992_));
 sky130_fd_sc_hd__o211a_1 _09391_ (.A1(_00988_),
    .A2(_00989_),
    .B1(_00981_),
    .C1(_00982_),
    .X(_00993_));
 sky130_fd_sc_hd__a22oi_2 _09392_ (.A1(_00981_),
    .A2(_00982_),
    .B1(_00990_),
    .B2(_00991_),
    .Y(_00994_));
 sky130_fd_sc_hd__a31o_1 _09393_ (.A1(_00831_),
    .A2(_00850_),
    .A3(_00851_),
    .B1(_00832_),
    .X(_00995_));
 sky130_fd_sc_hd__o21ai_1 _09394_ (.A1(_00993_),
    .A2(_00994_),
    .B1(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hd__a2111o_1 _09395_ (.A1(_00854_),
    .A2(_00831_),
    .B1(_00832_),
    .C1(_00993_),
    .D1(_00994_),
    .X(_00997_));
 sky130_fd_sc_hd__and3_1 _09396_ (.A(_00367_),
    .B(_02899_),
    .C(_00193_),
    .X(_00999_));
 sky130_fd_sc_hd__o32a_1 _09397_ (.A1(_02122_),
    .A2(_00361_),
    .A3(_00363_),
    .B1(net159),
    .B2(_00192_),
    .X(_01000_));
 sky130_fd_sc_hd__o32ai_1 _09398_ (.A1(_02122_),
    .A2(_00361_),
    .A3(_00363_),
    .B1(net159),
    .B2(_00192_),
    .Y(_01001_));
 sky130_fd_sc_hd__o22ai_1 _09399_ (.A1(_01620_),
    .A2(_00532_),
    .B1(_00999_),
    .B2(_01000_),
    .Y(_01002_));
 sky130_fd_sc_hd__or4_1 _09400_ (.A(_01620_),
    .B(_00532_),
    .C(_00999_),
    .D(_01000_),
    .X(_01003_));
 sky130_fd_sc_hd__nand2_1 _09401_ (.A(_01002_),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__nand3_1 _09402_ (.A(_00996_),
    .B(_00997_),
    .C(_01004_),
    .Y(_01005_));
 sky130_fd_sc_hd__a21o_1 _09403_ (.A1(_00996_),
    .A2(_00997_),
    .B1(_01004_),
    .X(_01006_));
 sky130_fd_sc_hd__a221o_1 _09404_ (.A1(_00824_),
    .A2(_00862_),
    .B1(_01005_),
    .B2(_01006_),
    .C1(_00860_),
    .X(_01007_));
 sky130_fd_sc_hd__nand3_1 _09405_ (.A(_01006_),
    .B(_00868_),
    .C(_01005_),
    .Y(_01008_));
 sky130_fd_sc_hd__nand2_2 _09406_ (.A(_01007_),
    .B(_01008_),
    .Y(_01010_));
 sky130_fd_sc_hd__o211ai_1 _09407_ (.A1(_00586_),
    .A2(_00645_),
    .B1(_00871_),
    .C1(_00874_),
    .Y(_01011_));
 sky130_fd_sc_hd__o21a_1 _09408_ (.A1(_00869_),
    .A2(_00870_),
    .B1(_01011_),
    .X(_01012_));
 sky130_fd_sc_hd__o211ai_1 _09409_ (.A1(_00869_),
    .A2(_00870_),
    .B1(_01008_),
    .C1(_01011_),
    .Y(_01013_));
 sky130_fd_sc_hd__xor2_4 _09410_ (.A(_01010_),
    .B(_01012_),
    .X(_01014_));
 sky130_fd_sc_hd__nand2_1 _09411_ (.A(_00977_),
    .B(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__or2_1 _09412_ (.A(_00977_),
    .B(_01014_),
    .X(_01016_));
 sky130_fd_sc_hd__and2_2 _09413_ (.A(_01015_),
    .B(_01016_),
    .X(_01017_));
 sky130_fd_sc_hd__nand2_2 _09414_ (.A(_01015_),
    .B(_01016_),
    .Y(_01018_));
 sky130_fd_sc_hd__a22o_1 _09415_ (.A1(_00816_),
    .A2(_00916_),
    .B1(_01015_),
    .B2(_01016_),
    .X(_01019_));
 sky130_fd_sc_hd__nand2_2 _09416_ (.A(_00917_),
    .B(_01017_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _09417_ (.A(_01019_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__o211ai_4 _09418_ (.A1(_00585_),
    .A2(_00718_),
    .B1(_00881_),
    .C1(_00883_),
    .Y(_01023_));
 sky130_fd_sc_hd__o211ai_4 _09419_ (.A1(_00584_),
    .A2(_00719_),
    .B1(_00880_),
    .C1(_00882_),
    .Y(_01024_));
 sky130_fd_sc_hd__o211ai_1 _09420_ (.A1(_00751_),
    .A2(_00877_),
    .B1(_01022_),
    .C1(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__o2111ai_1 _09421_ (.A1(_00752_),
    .A2(_00879_),
    .B1(_01019_),
    .C1(_01021_),
    .D1(_01023_),
    .Y(_01026_));
 sky130_fd_sc_hd__o211ai_1 _09422_ (.A1(_00879_),
    .A2(_00752_),
    .B1(_01023_),
    .C1(_01022_),
    .Y(_01027_));
 sky130_fd_sc_hd__o2111ai_1 _09423_ (.A1(_00751_),
    .A2(_00877_),
    .B1(_01019_),
    .C1(_01021_),
    .D1(_01024_),
    .Y(_01028_));
 sky130_fd_sc_hd__nor2_4 _09424_ (.A(net40),
    .B(net41),
    .Y(_01029_));
 sky130_fd_sc_hd__or2_2 _09425_ (.A(net40),
    .B(net41),
    .X(_01030_));
 sky130_fd_sc_hd__nand4b_4 _09426_ (.A_N(_00143_),
    .B(_00573_),
    .C(_01029_),
    .D(_00551_),
    .Y(_01032_));
 sky130_fd_sc_hd__a21oi_4 _09427_ (.A1(_01032_),
    .A2(net173),
    .B1(net42),
    .Y(_01033_));
 sky130_fd_sc_hd__a21o_4 _09428_ (.A1(_01032_),
    .A2(net173),
    .B1(net42),
    .X(_01034_));
 sky130_fd_sc_hd__o311a_4 _09429_ (.A1(net40),
    .A2(net41),
    .A3(_00575_),
    .B1(net42),
    .C1(net173),
    .X(_01035_));
 sky130_fd_sc_hd__o211ai_4 _09430_ (.A1(_00575_),
    .A2(_01030_),
    .B1(net173),
    .C1(net42),
    .Y(_01036_));
 sky130_fd_sc_hd__nand2_8 _09431_ (.A(_01034_),
    .B(_01036_),
    .Y(_01037_));
 sky130_fd_sc_hd__nor2_8 _09432_ (.A(_01033_),
    .B(_01035_),
    .Y(_01038_));
 sky130_fd_sc_hd__a31oi_1 _09433_ (.A1(_01032_),
    .A2(net42),
    .A3(net173),
    .B1(_00288_),
    .Y(_01039_));
 sky130_fd_sc_hd__nand2_2 _09434_ (.A(_01034_),
    .B(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__and3_1 _09435_ (.A(_00745_),
    .B(_01034_),
    .C(_01039_),
    .X(_01041_));
 sky130_fd_sc_hd__xor2_1 _09436_ (.A(_00745_),
    .B(_01040_),
    .X(_01043_));
 sky130_fd_sc_hd__o21ai_1 _09437_ (.A1(net166),
    .A2(_00580_),
    .B1(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__or3_1 _09438_ (.A(_01150_),
    .B(_01161_),
    .C(_01043_),
    .X(_01045_));
 sky130_fd_sc_hd__o31a_1 _09439_ (.A1(_00576_),
    .A2(_00578_),
    .A3(_01045_),
    .B1(_01044_),
    .X(_01046_));
 sky130_fd_sc_hd__nor2_2 _09440_ (.A(_00748_),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__and4_2 _09441_ (.A(net1),
    .B(_01046_),
    .C(_00581_),
    .D(_00745_),
    .X(_01048_));
 sky130_fd_sc_hd__nor2_1 _09442_ (.A(_01047_),
    .B(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__o211ai_2 _09443_ (.A1(_01047_),
    .A2(_01048_),
    .B1(_01027_),
    .C1(_01028_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand3_1 _09444_ (.A(_01025_),
    .B(_01026_),
    .C(_01049_),
    .Y(_01051_));
 sky130_fd_sc_hd__nor2_4 _09445_ (.A(net8),
    .B(net9),
    .Y(_01052_));
 sky130_fd_sc_hd__nand4b_4 _09446_ (.A_N(_00185_),
    .B(_00524_),
    .C(_00890_),
    .D(_00605_),
    .Y(_01053_));
 sky130_fd_sc_hd__a21oi_4 _09447_ (.A1(_01053_),
    .A2(net174),
    .B1(net10),
    .Y(_01054_));
 sky130_fd_sc_hd__a21o_4 _09448_ (.A1(_01053_),
    .A2(net174),
    .B1(net10),
    .X(_01055_));
 sky130_fd_sc_hd__o311a_4 _09449_ (.A1(_00891_),
    .A2(net9),
    .A3(_00526_),
    .B1(net10),
    .C1(net174),
    .X(_01056_));
 sky130_fd_sc_hd__o211ai_4 _09450_ (.A1(net9),
    .A2(_00892_),
    .B1(net10),
    .C1(net174),
    .Y(_01057_));
 sky130_fd_sc_hd__nand2_8 _09451_ (.A(_01055_),
    .B(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__nor2_8 _09452_ (.A(_01054_),
    .B(_01056_),
    .Y(_01059_));
 sky130_fd_sc_hd__o211ai_4 _09453_ (.A1(_01238_),
    .A2(_01249_),
    .B1(net147),
    .C1(net146),
    .Y(_01060_));
 sky130_fd_sc_hd__a32o_1 _09454_ (.A1(_00911_),
    .A2(_00899_),
    .A3(_00902_),
    .B1(_00569_),
    .B2(_01303_),
    .X(_01061_));
 sky130_fd_sc_hd__nand4_2 _09455_ (.A(_00569_),
    .B(_00904_),
    .C(_00911_),
    .D(_01303_),
    .Y(_01062_));
 sky130_fd_sc_hd__o2bb2a_1 _09456_ (.A1_N(_01061_),
    .A2_N(_01062_),
    .B1(_00310_),
    .B2(_01058_),
    .X(_01064_));
 sky130_fd_sc_hd__and4_1 _09457_ (.A(_01061_),
    .B(net33),
    .C(net141),
    .D(_01062_),
    .X(_01065_));
 sky130_fd_sc_hd__o32a_1 _09458_ (.A1(_00900_),
    .A2(_00903_),
    .A3(_00571_),
    .B1(_01065_),
    .B2(_01064_),
    .X(_01066_));
 sky130_fd_sc_hd__o2111a_1 _09459_ (.A1(_01292_),
    .A2(net141),
    .B1(_00569_),
    .C1(net33),
    .D1(_00905_),
    .X(_01067_));
 sky130_fd_sc_hd__nor3_2 _09460_ (.A(_01065_),
    .B(_00906_),
    .C(_01064_),
    .Y(_01068_));
 sky130_fd_sc_hd__nor2_1 _09461_ (.A(_01066_),
    .B(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand3_1 _09462_ (.A(_01050_),
    .B(_01051_),
    .C(_01069_),
    .Y(_01070_));
 sky130_fd_sc_hd__o2bb2ai_2 _09463_ (.A1_N(_01050_),
    .A2_N(_01051_),
    .B1(_01066_),
    .B2(_01068_),
    .Y(_01071_));
 sky130_fd_sc_hd__a21oi_2 _09464_ (.A1(_00887_),
    .A2(_00908_),
    .B1(_00888_),
    .Y(_01072_));
 sky130_fd_sc_hd__and3_1 _09465_ (.A(_01070_),
    .B(_01071_),
    .C(_01072_),
    .X(_01073_));
 sky130_fd_sc_hd__nand3_2 _09466_ (.A(_01070_),
    .B(_01071_),
    .C(_01072_),
    .Y(_01075_));
 sky130_fd_sc_hd__a21oi_2 _09467_ (.A1(_01070_),
    .A2(_01071_),
    .B1(_01072_),
    .Y(_01076_));
 sky130_fd_sc_hd__nor2_1 _09468_ (.A(_01073_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__xor2_1 _09469_ (.A(_00913_),
    .B(_01077_),
    .X(_01078_));
 sky130_fd_sc_hd__xnor2_1 _09470_ (.A(_00915_),
    .B(_01078_),
    .Y(net74));
 sky130_fd_sc_hd__or4b_4 _09471_ (.A(_00562_),
    .B(_00730_),
    .C(_00914_),
    .D_N(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__o21a_1 _09472_ (.A1(_00913_),
    .A2(_01076_),
    .B1(_01075_),
    .X(_01080_));
 sky130_fd_sc_hd__o221a_1 _09473_ (.A1(_00321_),
    .A2(_07537_),
    .B1(_05370_),
    .B2(_05359_),
    .C1(_07536_),
    .X(_01081_));
 sky130_fd_sc_hd__o32a_1 _09474_ (.A1(_07508_),
    .A2(_07510_),
    .A3(_05327_),
    .B1(_07189_),
    .B2(net153),
    .X(_01082_));
 sky130_fd_sc_hd__and3_1 _09475_ (.A(_07513_),
    .B(_05316_),
    .C(_07200_),
    .X(_01083_));
 sky130_fd_sc_hd__a21oi_1 _09476_ (.A1(_01083_),
    .A2(net151),
    .B1(_01082_),
    .Y(_01085_));
 sky130_fd_sc_hd__and3_1 _09477_ (.A(_01085_),
    .B(_06341_),
    .C(_07440_),
    .X(_01086_));
 sky130_fd_sc_hd__a31o_1 _09478_ (.A1(_06341_),
    .A2(_07436_),
    .A3(net154),
    .B1(_01085_),
    .X(_01087_));
 sky130_fd_sc_hd__and2b_1 _09479_ (.A_N(_01086_),
    .B(_01087_),
    .X(_01088_));
 sky130_fd_sc_hd__xnor2_1 _09480_ (.A(_01081_),
    .B(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__nor4_1 _09481_ (.A(_05327_),
    .B(net153),
    .C(_00754_),
    .D(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__or4_1 _09482_ (.A(_05327_),
    .B(net153),
    .C(_00754_),
    .D(_01089_),
    .X(_01091_));
 sky130_fd_sc_hd__o31a_1 _09483_ (.A1(_05327_),
    .A2(net153),
    .A3(_00754_),
    .B1(_01089_),
    .X(_01092_));
 sky130_fd_sc_hd__or2_1 _09484_ (.A(_01090_),
    .B(_01092_),
    .X(_01093_));
 sky130_fd_sc_hd__a21boi_2 _09485_ (.A1(_00755_),
    .A2(_00922_),
    .B1_N(_00923_),
    .Y(_01094_));
 sky130_fd_sc_hd__xnor2_1 _09486_ (.A(_01093_),
    .B(_01094_),
    .Y(_01096_));
 sky130_fd_sc_hd__or4_1 _09487_ (.A(_01958_),
    .B(_02636_),
    .C(_00274_),
    .D(_00428_),
    .X(_01097_));
 sky130_fd_sc_hd__o32a_1 _09488_ (.A1(_02636_),
    .A2(_00270_),
    .A3(_00272_),
    .B1(_00428_),
    .B2(_01958_),
    .X(_01098_));
 sky130_fd_sc_hd__a32o_1 _09489_ (.A1(_01969_),
    .A2(_00425_),
    .A3(_00427_),
    .B1(_02647_),
    .B2(_00275_),
    .X(_01099_));
 sky130_fd_sc_hd__a311o_1 _09490_ (.A1(_02647_),
    .A2(_00429_),
    .A3(_00930_),
    .B1(_00955_),
    .C1(_01098_),
    .X(_01100_));
 sky130_fd_sc_hd__a211o_1 _09491_ (.A1(_01097_),
    .A2(_01099_),
    .B1(_03906_),
    .C1(net143),
    .X(_01101_));
 sky130_fd_sc_hd__nand2_1 _09492_ (.A(_01100_),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__o32a_1 _09493_ (.A1(_03906_),
    .A2(net143),
    .A3(_00664_),
    .B1(_00953_),
    .B2(_00956_),
    .X(_01103_));
 sky130_fd_sc_hd__a21o_1 _09494_ (.A1(_00935_),
    .A2(_00937_),
    .B1(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__nand2_1 _09495_ (.A(_00938_),
    .B(_01103_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand4_1 _09496_ (.A(_01100_),
    .B(_01101_),
    .C(_01104_),
    .D(_01105_),
    .Y(_01107_));
 sky130_fd_sc_hd__a22o_1 _09497_ (.A1(_01100_),
    .A2(_01101_),
    .B1(_01104_),
    .B2(_01105_),
    .X(_01108_));
 sky130_fd_sc_hd__a21boi_2 _09498_ (.A1(_01102_),
    .A2(_01105_),
    .B1_N(_01104_),
    .Y(_01109_));
 sky130_fd_sc_hd__and3_1 _09499_ (.A(_00944_),
    .B(_01107_),
    .C(_01108_),
    .X(_01110_));
 sky130_fd_sc_hd__o2111ai_1 _09500_ (.A1(_00940_),
    .A2(_00941_),
    .B1(_01107_),
    .C1(_01108_),
    .D1(_00929_),
    .Y(_01111_));
 sky130_fd_sc_hd__a21o_1 _09501_ (.A1(_01107_),
    .A2(_01108_),
    .B1(_00944_),
    .X(_01112_));
 sky130_fd_sc_hd__a22oi_1 _09502_ (.A1(_04255_),
    .A2(_00010_),
    .B1(_01111_),
    .B2(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__o2111ai_1 _09503_ (.A1(_00003_),
    .A2(_00004_),
    .B1(_01111_),
    .C1(_01112_),
    .D1(_04255_),
    .Y(_01114_));
 sky130_fd_sc_hd__and2b_2 _09504_ (.A_N(_01113_),
    .B(_01114_),
    .X(_01115_));
 sky130_fd_sc_hd__inv_2 _09505_ (.A(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__a21o_2 _09506_ (.A1(_00949_),
    .A2(_00958_),
    .B1(_00950_),
    .X(_01118_));
 sky130_fd_sc_hd__inv_2 _09507_ (.A(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand2_1 _09508_ (.A(_01115_),
    .B(_01118_),
    .Y(_01120_));
 sky130_fd_sc_hd__a211o_1 _09509_ (.A1(_00958_),
    .A2(_00949_),
    .B1(_00950_),
    .C1(_01115_),
    .X(_01121_));
 sky130_fd_sc_hd__o211ai_2 _09510_ (.A1(_00759_),
    .A2(_00807_),
    .B1(_00963_),
    .C1(_00969_),
    .Y(_01122_));
 sky130_fd_sc_hd__o211ai_2 _09511_ (.A1(_00964_),
    .A2(_00960_),
    .B1(_00808_),
    .C1(_00968_),
    .Y(_01123_));
 sky130_fd_sc_hd__a22o_1 _09512_ (.A1(_01120_),
    .A2(_01121_),
    .B1(_01123_),
    .B2(_00963_),
    .X(_01124_));
 sky130_fd_sc_hd__nand4_1 _09513_ (.A(_00963_),
    .B(_01120_),
    .C(_01121_),
    .D(_01123_),
    .Y(_01125_));
 sky130_fd_sc_hd__a21oi_1 _09514_ (.A1(_01124_),
    .A2(_01125_),
    .B1(_01096_),
    .Y(_01126_));
 sky130_fd_sc_hd__a21o_1 _09515_ (.A1(_01124_),
    .A2(_01125_),
    .B1(_01096_),
    .X(_01127_));
 sky130_fd_sc_hd__nand3_1 _09516_ (.A(_01124_),
    .B(_01125_),
    .C(_01096_),
    .Y(_01129_));
 sky130_fd_sc_hd__a21boi_1 _09517_ (.A1(_00996_),
    .A2(_01004_),
    .B1_N(_00997_),
    .Y(_01130_));
 sky130_fd_sc_hd__o2111ai_4 _09518_ (.A1(_00299_),
    .A2(_03511_),
    .B1(_00072_),
    .C1(_00985_),
    .D1(_03490_),
    .Y(_01131_));
 sky130_fd_sc_hd__o32a_1 _09519_ (.A1(_02910_),
    .A2(_00192_),
    .A3(_00366_),
    .B1(_00532_),
    .B2(_01620_),
    .X(_01132_));
 sky130_fd_sc_hd__o211a_1 _09520_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_00533_),
    .C1(_01001_),
    .X(_01133_));
 sky130_fd_sc_hd__o211ai_2 _09521_ (.A1(_01000_),
    .A2(_01132_),
    .B1(_01131_),
    .C1(_00986_),
    .Y(_01134_));
 sky130_fd_sc_hd__o2bb2ai_1 _09522_ (.A1_N(_00986_),
    .A2_N(_01131_),
    .B1(_01133_),
    .B2(_00999_),
    .Y(_01135_));
 sky130_fd_sc_hd__and3_1 _09523_ (.A(_02866_),
    .B(_00362_),
    .C(_00364_),
    .X(_01136_));
 sky130_fd_sc_hd__a32o_1 _09524_ (.A1(net156),
    .A2(_00189_),
    .A3(_00191_),
    .B1(_04726_),
    .B2(_00072_),
    .X(_01137_));
 sky130_fd_sc_hd__or3_1 _09525_ (.A(_04671_),
    .B(_04693_),
    .C(_00190_),
    .X(_01138_));
 sky130_fd_sc_hd__and4_1 _09526_ (.A(net156),
    .B(_04726_),
    .C(_00072_),
    .D(_00193_),
    .X(_01140_));
 sky130_fd_sc_hd__or4_1 _09527_ (.A(_03544_),
    .B(_04715_),
    .C(net148),
    .D(_00192_),
    .X(_01141_));
 sky130_fd_sc_hd__a32o_1 _09528_ (.A1(_02866_),
    .A2(_00362_),
    .A3(_00364_),
    .B1(_01137_),
    .B2(_01141_),
    .X(_01142_));
 sky130_fd_sc_hd__nand4_1 _09529_ (.A(_02866_),
    .B(_00367_),
    .C(_01137_),
    .D(_01141_),
    .Y(_01143_));
 sky130_fd_sc_hd__a22o_1 _09530_ (.A1(_01134_),
    .A2(_01135_),
    .B1(_01142_),
    .B2(_01143_),
    .X(_01144_));
 sky130_fd_sc_hd__nand4_1 _09531_ (.A(_01134_),
    .B(_01135_),
    .C(_01142_),
    .D(_01143_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand2_1 _09532_ (.A(_01144_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__a21boi_1 _09533_ (.A1(_00992_),
    .A2(_00981_),
    .B1_N(_00982_),
    .Y(_01147_));
 sky130_fd_sc_hd__or2_1 _09534_ (.A(_01146_),
    .B(_01147_),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_01146_),
    .B(_01147_),
    .Y(_01149_));
 sky130_fd_sc_hd__nand2_1 _09536_ (.A(_01148_),
    .B(_01149_),
    .Y(_01151_));
 sky130_fd_sc_hd__o31a_1 _09537_ (.A1(_02079_),
    .A2(_02100_),
    .A3(_00532_),
    .B1(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__a211oi_1 _09538_ (.A1(_02046_),
    .A2(_02068_),
    .B1(_00532_),
    .C1(_01151_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor2_1 _09539_ (.A(_01152_),
    .B(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand2_1 _09540_ (.A(_01154_),
    .B(_01130_),
    .Y(_01155_));
 sky130_fd_sc_hd__or2_1 _09541_ (.A(_01130_),
    .B(_01154_),
    .X(_01156_));
 sky130_fd_sc_hd__nand2_1 _09542_ (.A(_01155_),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(_01007_),
    .B(_01013_),
    .Y(_01158_));
 sky130_fd_sc_hd__xnor2_2 _09544_ (.A(_01157_),
    .B(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__a21o_1 _09545_ (.A1(_01127_),
    .A2(_01129_),
    .B1(_01159_),
    .X(_01160_));
 sky130_fd_sc_hd__nand2_1 _09546_ (.A(_01129_),
    .B(_01159_),
    .Y(_01162_));
 sky130_fd_sc_hd__o21a_2 _09547_ (.A1(_01126_),
    .A2(_01162_),
    .B1(_01160_),
    .X(_01163_));
 sky130_fd_sc_hd__a21boi_4 _09548_ (.A1(_00975_),
    .A2(_01014_),
    .B1_N(_00974_),
    .Y(_01164_));
 sky130_fd_sc_hd__nand2_4 _09549_ (.A(_01163_),
    .B(_01164_),
    .Y(_01165_));
 sky130_fd_sc_hd__or2_2 _09550_ (.A(_01164_),
    .B(_01163_),
    .X(_01166_));
 sky130_fd_sc_hd__nand2_1 _09551_ (.A(_01165_),
    .B(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__o211ai_4 _09552_ (.A1(_00751_),
    .A2(_00877_),
    .B1(_01021_),
    .C1(_01024_),
    .Y(_01168_));
 sky130_fd_sc_hd__o211ai_4 _09553_ (.A1(_00752_),
    .A2(_00879_),
    .B1(_01019_),
    .C1(_01023_),
    .Y(_01169_));
 sky130_fd_sc_hd__o211ai_2 _09554_ (.A1(_00917_),
    .A2(_01017_),
    .B1(_01167_),
    .C1(_01168_),
    .Y(_01170_));
 sky130_fd_sc_hd__o2111ai_2 _09555_ (.A1(_00918_),
    .A2(_01018_),
    .B1(_01165_),
    .C1(_01166_),
    .D1(_01169_),
    .Y(_01171_));
 sky130_fd_sc_hd__o2111ai_1 _09556_ (.A1(_00917_),
    .A2(_01017_),
    .B1(_01165_),
    .C1(_01166_),
    .D1(_01168_),
    .Y(_01173_));
 sky130_fd_sc_hd__o211ai_1 _09557_ (.A1(_00918_),
    .A2(_01018_),
    .B1(_01167_),
    .C1(_01169_),
    .Y(_01174_));
 sky130_fd_sc_hd__o2111ai_1 _09558_ (.A1(net164),
    .A2(_01040_),
    .B1(_00581_),
    .C1(net1),
    .D1(_00745_),
    .Y(_01175_));
 sky130_fd_sc_hd__o31a_2 _09559_ (.A1(net166),
    .A2(_00580_),
    .A3(_01043_),
    .B1(_01175_),
    .X(_01176_));
 sky130_fd_sc_hd__and3_1 _09560_ (.A(_01499_),
    .B(_00577_),
    .C(_00579_),
    .X(_01177_));
 sky130_fd_sc_hd__nor2_1 _09561_ (.A(net41),
    .B(net42),
    .Y(_01178_));
 sky130_fd_sc_hd__nor3_4 _09562_ (.A(_01030_),
    .B(net42),
    .C(_00575_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand4b_4 _09563_ (.A_N(_00263_),
    .B(_00573_),
    .C(_01029_),
    .D(_00616_),
    .Y(_01180_));
 sky130_fd_sc_hd__o311a_4 _09564_ (.A1(_01030_),
    .A2(net42),
    .A3(_00575_),
    .B1(_00638_),
    .C1(net173),
    .X(_01181_));
 sky130_fd_sc_hd__a21oi_4 _09565_ (.A1(_01180_),
    .A2(net173),
    .B1(_00638_),
    .Y(_01182_));
 sky130_fd_sc_hd__a21oi_4 _09566_ (.A1(_01180_),
    .A2(net173),
    .B1(net43),
    .Y(_01184_));
 sky130_fd_sc_hd__o21ai_4 _09567_ (.A1(_00299_),
    .A2(_01179_),
    .B1(_00638_),
    .Y(_01185_));
 sky130_fd_sc_hd__o311a_4 _09568_ (.A1(_01030_),
    .A2(net42),
    .A3(_00575_),
    .B1(net43),
    .C1(net173),
    .X(_01186_));
 sky130_fd_sc_hd__o211ai_4 _09569_ (.A1(net42),
    .A2(_01032_),
    .B1(net43),
    .C1(net173),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_8 _09570_ (.A(_01185_),
    .B(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__nor2_8 _09571_ (.A(_01184_),
    .B(_01186_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand3_4 _09572_ (.A(_01185_),
    .B(_01187_),
    .C(net1),
    .Y(_01190_));
 sky130_fd_sc_hd__o21ai_2 _09573_ (.A1(_00987_),
    .A2(_01037_),
    .B1(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__o22ai_4 _09574_ (.A1(net172),
    .A2(_00943_),
    .B1(_01181_),
    .B2(_01182_),
    .Y(_01192_));
 sky130_fd_sc_hd__or4_1 _09575_ (.A(_00987_),
    .B(_01184_),
    .C(_01186_),
    .D(_01040_),
    .X(_01193_));
 sky130_fd_sc_hd__o21ai_1 _09576_ (.A1(_01040_),
    .A2(_01192_),
    .B1(_01191_),
    .Y(_01195_));
 sky130_fd_sc_hd__o2111a_1 _09577_ (.A1(_01040_),
    .A2(_01192_),
    .B1(_00743_),
    .C1(_01191_),
    .D1(net164),
    .X(_01196_));
 sky130_fd_sc_hd__o2111ai_4 _09578_ (.A1(_01040_),
    .A2(_01192_),
    .B1(_00743_),
    .C1(_01191_),
    .D1(net164),
    .Y(_01197_));
 sky130_fd_sc_hd__o31a_1 _09579_ (.A1(_01150_),
    .A2(_01161_),
    .A3(_00744_),
    .B1(_01195_),
    .X(_01198_));
 sky130_fd_sc_hd__o21ai_2 _09580_ (.A1(net166),
    .A2(_00744_),
    .B1(_01195_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _09581_ (.A(_01197_),
    .B(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__a32o_1 _09582_ (.A1(_01499_),
    .A2(_00577_),
    .A3(_00579_),
    .B1(_01197_),
    .B2(_01199_),
    .X(_01201_));
 sky130_fd_sc_hd__o2111ai_4 _09583_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_00581_),
    .C1(_01197_),
    .D1(_01199_),
    .Y(_01202_));
 sky130_fd_sc_hd__a311o_2 _09584_ (.A1(_01499_),
    .A2(_00577_),
    .A3(_00579_),
    .B1(_01196_),
    .C1(_01198_),
    .X(_01203_));
 sky130_fd_sc_hd__nand3_1 _09585_ (.A(_01201_),
    .B(_01202_),
    .C(_01041_),
    .Y(_01204_));
 sky130_fd_sc_hd__a21oi_2 _09586_ (.A1(_01200_),
    .A2(_01177_),
    .B1(_01041_),
    .Y(_01206_));
 sky130_fd_sc_hd__a32oi_4 _09587_ (.A1(_01041_),
    .A2(_01201_),
    .A3(_01202_),
    .B1(_01206_),
    .B2(_01203_),
    .Y(_01207_));
 sky130_fd_sc_hd__xor2_4 _09588_ (.A(_01176_),
    .B(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__nand3_2 _09589_ (.A(_01170_),
    .B(_01171_),
    .C(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand3b_2 _09590_ (.A_N(_01208_),
    .B(_01174_),
    .C(_01173_),
    .Y(_01210_));
 sky130_fd_sc_hd__or2_2 _09591_ (.A(net9),
    .B(net10),
    .X(_01211_));
 sky130_fd_sc_hd__nand4_1 _09592_ (.A(_00359_),
    .B(_00563_),
    .C(_01052_),
    .D(_00627_),
    .Y(_01212_));
 sky130_fd_sc_hd__o21ai_4 _09593_ (.A1(_00892_),
    .A2(_01211_),
    .B1(net174),
    .Y(_01213_));
 sky130_fd_sc_hd__a311o_4 _09594_ (.A1(_00564_),
    .A2(_01052_),
    .A3(_00627_),
    .B1(net11),
    .C1(_00321_),
    .X(_01214_));
 sky130_fd_sc_hd__nand2_4 _09595_ (.A(_01213_),
    .B(net11),
    .Y(_01215_));
 sky130_fd_sc_hd__o311a_4 _09596_ (.A1(_00526_),
    .A2(_00891_),
    .A3(_01211_),
    .B1(net11),
    .C1(net174),
    .X(_01217_));
 sky130_fd_sc_hd__o211ai_4 _09597_ (.A1(_00892_),
    .A2(_01211_),
    .B1(net174),
    .C1(net11),
    .Y(_01218_));
 sky130_fd_sc_hd__a21oi_4 _09598_ (.A1(_01212_),
    .A2(net174),
    .B1(net11),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_8 _09599_ (.A(_00649_),
    .B(_01213_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2_8 _09600_ (.A(_01218_),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_8 _09601_ (.A(_01214_),
    .B(_01215_),
    .Y(_01222_));
 sky130_fd_sc_hd__o211ai_4 _09602_ (.A1(_01532_),
    .A2(_01554_),
    .B1(net147),
    .C1(net146),
    .Y(_01223_));
 sky130_fd_sc_hd__o31a_1 _09603_ (.A1(_01292_),
    .A2(_00898_),
    .A3(_00901_),
    .B1(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__o21ai_1 _09604_ (.A1(_01292_),
    .A2(_00903_),
    .B1(_01223_),
    .Y(_01225_));
 sky130_fd_sc_hd__o211ai_4 _09605_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_00899_),
    .C1(_00902_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _09606_ (.A(_01060_),
    .B(_01226_),
    .Y(_01228_));
 sky130_fd_sc_hd__o32a_1 _09607_ (.A1(_00900_),
    .A2(_01054_),
    .A3(_01056_),
    .B1(_01224_),
    .B2(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__o22ai_1 _09608_ (.A1(_00900_),
    .A2(_01058_),
    .B1(_01224_),
    .B2(_01228_),
    .Y(_01230_));
 sky130_fd_sc_hd__o2111ai_2 _09609_ (.A1(_01060_),
    .A2(_01226_),
    .B1(_01225_),
    .C1(_00911_),
    .D1(net141),
    .Y(_01231_));
 sky130_fd_sc_hd__o2bb2ai_1 _09610_ (.A1_N(_01230_),
    .A2_N(_01231_),
    .B1(_00310_),
    .B2(_01221_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand4_1 _09611_ (.A(_01222_),
    .B(_01230_),
    .C(_01231_),
    .D(net33),
    .Y(_01233_));
 sky130_fd_sc_hd__a21bo_2 _09612_ (.A1(_01232_),
    .A2(_01233_),
    .B1_N(_01062_),
    .X(_01234_));
 sky130_fd_sc_hd__nand3b_2 _09613_ (.A_N(_01062_),
    .B(_01232_),
    .C(_01233_),
    .Y(_01235_));
 sky130_fd_sc_hd__nor2_1 _09614_ (.A(_01065_),
    .B(_01067_),
    .Y(_01236_));
 sky130_fd_sc_hd__a41o_1 _09615_ (.A1(net33),
    .A2(net141),
    .A3(_01061_),
    .A4(_01062_),
    .B1(_01067_),
    .X(_01237_));
 sky130_fd_sc_hd__a21oi_1 _09616_ (.A1(_01234_),
    .A2(_01235_),
    .B1(_01237_),
    .Y(_01239_));
 sky130_fd_sc_hd__and3_1 _09617_ (.A(_01234_),
    .B(_01235_),
    .C(_01237_),
    .X(_01240_));
 sky130_fd_sc_hd__a21oi_1 _09618_ (.A1(_01234_),
    .A2(_01235_),
    .B1(_01236_),
    .Y(_01241_));
 sky130_fd_sc_hd__and3_1 _09619_ (.A(_01234_),
    .B(_01235_),
    .C(_01236_),
    .X(_01242_));
 sky130_fd_sc_hd__nor2_1 _09620_ (.A(_01241_),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__o211a_1 _09621_ (.A1(_01241_),
    .A2(_01242_),
    .B1(_01209_),
    .C1(_01210_),
    .X(_01244_));
 sky130_fd_sc_hd__o211ai_2 _09622_ (.A1(_01241_),
    .A2(_01242_),
    .B1(_01209_),
    .C1(_01210_),
    .Y(_01245_));
 sky130_fd_sc_hd__a21boi_1 _09623_ (.A1(_01209_),
    .A2(_01210_),
    .B1_N(_01243_),
    .Y(_01246_));
 sky130_fd_sc_hd__o2bb2ai_1 _09624_ (.A1_N(_01209_),
    .A2_N(_01210_),
    .B1(_01239_),
    .B2(_01240_),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_1 _09625_ (.A(_01244_),
    .B(_01246_),
    .Y(_01248_));
 sky130_fd_sc_hd__a21bo_2 _09626_ (.A1(_01050_),
    .A2(_01069_),
    .B1_N(_01051_),
    .X(_01250_));
 sky130_fd_sc_hd__nand3_2 _09627_ (.A(_01245_),
    .B(_01247_),
    .C(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__a21o_1 _09628_ (.A1(_01245_),
    .A2(_01247_),
    .B1(_01250_),
    .X(_01252_));
 sky130_fd_sc_hd__nand2_1 _09629_ (.A(_01251_),
    .B(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hd__xor2_2 _09630_ (.A(_01080_),
    .B(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__a21oi_1 _09631_ (.A1(_00845_),
    .A2(_01079_),
    .B1(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__and3_1 _09632_ (.A(_00845_),
    .B(_01079_),
    .C(_01254_),
    .X(_01256_));
 sky130_fd_sc_hd__nor2_1 _09633_ (.A(_01255_),
    .B(_01256_),
    .Y(net75));
 sky130_fd_sc_hd__nor2_1 _09634_ (.A(_01079_),
    .B(_01254_),
    .Y(_01257_));
 sky130_fd_sc_hd__a22oi_4 _09635_ (.A1(_01206_),
    .A2(_01203_),
    .B1(_01176_),
    .B2(_01204_),
    .Y(_01258_));
 sky130_fd_sc_hd__a31o_1 _09636_ (.A1(_01499_),
    .A2(_00581_),
    .A3(_01199_),
    .B1(_01196_),
    .X(_01260_));
 sky130_fd_sc_hd__and3_1 _09637_ (.A(_01969_),
    .B(_00577_),
    .C(_00579_),
    .X(_01261_));
 sky130_fd_sc_hd__and3_1 _09638_ (.A(_01499_),
    .B(_00739_),
    .C(_00740_),
    .X(_01262_));
 sky130_fd_sc_hd__and3_1 _09639_ (.A(net164),
    .B(_01034_),
    .C(_01036_),
    .X(_01263_));
 sky130_fd_sc_hd__nor2_2 _09640_ (.A(net42),
    .B(net43),
    .Y(_01264_));
 sky130_fd_sc_hd__nand4b_4 _09641_ (.A_N(_00263_),
    .B(_00573_),
    .C(_01029_),
    .D(_01264_),
    .Y(_01265_));
 sky130_fd_sc_hd__o211ai_4 _09642_ (.A1(net43),
    .A2(_01180_),
    .B1(_00660_),
    .C1(net173),
    .Y(_01266_));
 sky130_fd_sc_hd__a21o_4 _09643_ (.A1(_01265_),
    .A2(net173),
    .B1(_00660_),
    .X(_01267_));
 sky130_fd_sc_hd__a21oi_1 _09644_ (.A1(_01265_),
    .A2(net173),
    .B1(net45),
    .Y(_01268_));
 sky130_fd_sc_hd__a21o_4 _09645_ (.A1(_01265_),
    .A2(net173),
    .B1(net45),
    .X(_01269_));
 sky130_fd_sc_hd__o211ai_4 _09646_ (.A1(net43),
    .A2(_01180_),
    .B1(net45),
    .C1(net173),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2_8 _09647_ (.A(_01269_),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_8 _09648_ (.A(_01266_),
    .B(_01267_),
    .Y(_01273_));
 sky130_fd_sc_hd__a31oi_1 _09649_ (.A1(_01265_),
    .A2(net45),
    .A3(net173),
    .B1(_00288_),
    .Y(_01274_));
 sky130_fd_sc_hd__a31o_1 _09650_ (.A1(_01265_),
    .A2(net45),
    .A3(net173),
    .B1(_00288_),
    .X(_01275_));
 sky130_fd_sc_hd__o21ai_2 _09651_ (.A1(_01268_),
    .A2(_01275_),
    .B1(_01192_),
    .Y(_01276_));
 sky130_fd_sc_hd__o211ai_4 _09652_ (.A1(net172),
    .A2(_00943_),
    .B1(_01269_),
    .C1(_01271_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand4_2 _09653_ (.A(_01189_),
    .B(_01274_),
    .C(_01269_),
    .D(_00998_),
    .Y(_01278_));
 sky130_fd_sc_hd__o21ai_1 _09654_ (.A1(_01190_),
    .A2(_01277_),
    .B1(_01276_),
    .Y(_01279_));
 sky130_fd_sc_hd__o211a_2 _09655_ (.A1(_01190_),
    .A2(_01277_),
    .B1(_01263_),
    .C1(_01276_),
    .X(_01280_));
 sky130_fd_sc_hd__o2111ai_2 _09656_ (.A1(_01095_),
    .A2(_01117_),
    .B1(_01038_),
    .C1(_01276_),
    .D1(_01278_),
    .Y(_01282_));
 sky130_fd_sc_hd__a2bb2oi_1 _09657_ (.A1_N(net166),
    .A2_N(_01037_),
    .B1(_01276_),
    .B2(_01278_),
    .Y(_01283_));
 sky130_fd_sc_hd__o21ai_1 _09658_ (.A1(net166),
    .A2(_01037_),
    .B1(_01279_),
    .Y(_01284_));
 sky130_fd_sc_hd__o2111ai_1 _09659_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_00743_),
    .C1(_01282_),
    .D1(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__o22ai_1 _09660_ (.A1(_01488_),
    .A2(_00744_),
    .B1(_01280_),
    .B2(_01283_),
    .Y(_01286_));
 sky130_fd_sc_hd__o21ai_1 _09661_ (.A1(_01280_),
    .A2(_01283_),
    .B1(_01262_),
    .Y(_01287_));
 sky130_fd_sc_hd__o211ai_1 _09662_ (.A1(_01488_),
    .A2(_00744_),
    .B1(_01282_),
    .C1(_01284_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand3b_2 _09663_ (.A_N(_01193_),
    .B(_01285_),
    .C(_01286_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand3_2 _09664_ (.A(_01193_),
    .B(_01287_),
    .C(_01288_),
    .Y(_01290_));
 sky130_fd_sc_hd__a21oi_2 _09665_ (.A1(_01289_),
    .A2(_01290_),
    .B1(_01261_),
    .Y(_01291_));
 sky130_fd_sc_hd__a32o_1 _09666_ (.A1(_01936_),
    .A2(_01947_),
    .A3(_00581_),
    .B1(_01289_),
    .B2(_01290_),
    .X(_01293_));
 sky130_fd_sc_hd__o2111a_1 _09667_ (.A1(_01892_),
    .A2(_01914_),
    .B1(_00581_),
    .C1(_01289_),
    .D1(_01290_),
    .X(_01294_));
 sky130_fd_sc_hd__o2111ai_2 _09668_ (.A1(_01892_),
    .A2(_01914_),
    .B1(_00581_),
    .C1(_01289_),
    .D1(_01290_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _09669_ (.A(_01295_),
    .B(_01260_),
    .Y(_01296_));
 sky130_fd_sc_hd__a21oi_1 _09670_ (.A1(_01293_),
    .A2(_01295_),
    .B1(_01260_),
    .Y(_01297_));
 sky130_fd_sc_hd__o21bai_2 _09671_ (.A1(_01291_),
    .A2(_01294_),
    .B1_N(_01260_),
    .Y(_01298_));
 sky130_fd_sc_hd__o21ai_2 _09672_ (.A1(_01291_),
    .A2(_01296_),
    .B1(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__a31oi_1 _09673_ (.A1(_01293_),
    .A2(_01295_),
    .A3(_01260_),
    .B1(_01258_),
    .Y(_01300_));
 sky130_fd_sc_hd__a2bb2oi_4 _09674_ (.A1_N(_01296_),
    .A2_N(_01291_),
    .B1(_01258_),
    .B2(_01298_),
    .Y(_01301_));
 sky130_fd_sc_hd__xnor2_4 _09675_ (.A(_01258_),
    .B(_01299_),
    .Y(_01302_));
 sky130_fd_sc_hd__o21a_2 _09676_ (.A1(_01126_),
    .A2(_01159_),
    .B1(_01129_),
    .X(_01304_));
 sky130_fd_sc_hd__o2bb2ai_1 _09677_ (.A1_N(_01007_),
    .A2_N(_01013_),
    .B1(_01130_),
    .B2(_01154_),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_2 _09678_ (.A(_01155_),
    .B(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__o21ai_1 _09679_ (.A1(_01136_),
    .A2(_01140_),
    .B1(_01137_),
    .Y(_01307_));
 sky130_fd_sc_hd__and3_1 _09680_ (.A(_02866_),
    .B(_00528_),
    .C(_00531_),
    .X(_01308_));
 sky130_fd_sc_hd__or3_1 _09681_ (.A(_03479_),
    .B(_03522_),
    .C(_00363_),
    .X(_01309_));
 sky130_fd_sc_hd__a32o_1 _09682_ (.A1(net156),
    .A2(_00362_),
    .A3(_00364_),
    .B1(_04726_),
    .B2(_00193_),
    .X(_01310_));
 sky130_fd_sc_hd__o41a_1 _09683_ (.A1(_00188_),
    .A2(_00361_),
    .A3(_01138_),
    .A4(_01309_),
    .B1(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__xnor2_1 _09684_ (.A(_01308_),
    .B(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__a21bo_1 _09685_ (.A1(_01142_),
    .A2(_01143_),
    .B1_N(_01135_),
    .X(_01313_));
 sky130_fd_sc_hd__and3b_1 _09686_ (.A_N(_01312_),
    .B(_01313_),
    .C(_01134_),
    .X(_01315_));
 sky130_fd_sc_hd__a21boi_1 _09687_ (.A1(_01134_),
    .A2(_01313_),
    .B1_N(_01312_),
    .Y(_01316_));
 sky130_fd_sc_hd__o21ba_1 _09688_ (.A1(_01307_),
    .A2(_01316_),
    .B1_N(_01315_),
    .X(_01317_));
 sky130_fd_sc_hd__or3_1 _09689_ (.A(_01307_),
    .B(_01315_),
    .C(_01316_),
    .X(_01318_));
 sky130_fd_sc_hd__o21ai_1 _09690_ (.A1(_01315_),
    .A2(_01316_),
    .B1(_01307_),
    .Y(_01319_));
 sky130_fd_sc_hd__a2bb2o_1 _09691_ (.A1_N(_01146_),
    .A2_N(_01147_),
    .B1(_02133_),
    .B2(_00533_),
    .X(_01320_));
 sky130_fd_sc_hd__a22o_1 _09692_ (.A1(_01318_),
    .A2(_01319_),
    .B1(_01320_),
    .B2(_01149_),
    .X(_01321_));
 sky130_fd_sc_hd__o2111ai_1 _09693_ (.A1(_01315_),
    .A2(_01317_),
    .B1(_01319_),
    .C1(_01320_),
    .D1(_01149_),
    .Y(_01322_));
 sky130_fd_sc_hd__and2_1 _09694_ (.A(_01321_),
    .B(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__nand3_1 _09695_ (.A(_01155_),
    .B(_01305_),
    .C(_01322_),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2_2 _09696_ (.A(_01321_),
    .B(_01324_),
    .Y(_01326_));
 sky130_fd_sc_hd__xnor2_4 _09697_ (.A(_01306_),
    .B(_01323_),
    .Y(_01327_));
 sky130_fd_sc_hd__a31o_1 _09698_ (.A1(_05436_),
    .A2(_07540_),
    .A3(_01087_),
    .B1(_01086_),
    .X(_01328_));
 sky130_fd_sc_hd__o221a_1 _09699_ (.A1(_00063_),
    .A2(_00066_),
    .B1(_05359_),
    .B2(_05370_),
    .C1(_00070_),
    .X(_01329_));
 sky130_fd_sc_hd__a32o_1 _09700_ (.A1(_05316_),
    .A2(_00006_),
    .A3(_00008_),
    .B1(_07200_),
    .B2(_07513_),
    .X(_01330_));
 sky130_fd_sc_hd__nand4_4 _09701_ (.A(_07200_),
    .B(_00006_),
    .C(_00008_),
    .D(_05316_),
    .Y(_01331_));
 sky130_fd_sc_hd__o21ai_1 _09702_ (.A1(_07512_),
    .A2(_01331_),
    .B1(_01330_),
    .Y(_01332_));
 sky130_fd_sc_hd__o21a_1 _09703_ (.A1(net153),
    .A2(_07441_),
    .B1(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__o2111a_1 _09704_ (.A1(_01331_),
    .A2(_07512_),
    .B1(_07440_),
    .C1(net151),
    .D1(_01330_),
    .X(_01334_));
 sky130_fd_sc_hd__or3_1 _09705_ (.A(net153),
    .B(_07441_),
    .C(_01332_),
    .X(_01335_));
 sky130_fd_sc_hd__o22ai_1 _09706_ (.A1(_06331_),
    .A2(_07539_),
    .B1(_01333_),
    .B2(_01334_),
    .Y(_01337_));
 sky130_fd_sc_hd__a2111o_1 _09707_ (.A1(_06276_),
    .A2(_06298_),
    .B1(_07539_),
    .C1(_01333_),
    .D1(_01334_),
    .X(_01338_));
 sky130_fd_sc_hd__nand2_1 _09708_ (.A(_01337_),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__a21bo_1 _09709_ (.A1(net151),
    .A2(_01083_),
    .B1_N(_01339_),
    .X(_01340_));
 sky130_fd_sc_hd__or3b_1 _09710_ (.A(_01339_),
    .B(net153),
    .C_N(_01083_),
    .X(_01341_));
 sky130_fd_sc_hd__a21oi_1 _09711_ (.A1(_01340_),
    .A2(_01341_),
    .B1(_01329_),
    .Y(_01342_));
 sky130_fd_sc_hd__and3_1 _09712_ (.A(_01341_),
    .B(_01329_),
    .C(_01340_),
    .X(_01343_));
 sky130_fd_sc_hd__nor2_1 _09713_ (.A(_01342_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2_1 _09714_ (.A(_01344_),
    .B(_01328_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _09715_ (.A(_01328_),
    .B(_01344_),
    .Y(_01346_));
 sky130_fd_sc_hd__xnor2_1 _09716_ (.A(_01328_),
    .B(_01344_),
    .Y(_01348_));
 sky130_fd_sc_hd__o21a_1 _09717_ (.A1(_01092_),
    .A2(_01094_),
    .B1(_01091_),
    .X(_01349_));
 sky130_fd_sc_hd__nor2_1 _09718_ (.A(_01348_),
    .B(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__o211a_1 _09719_ (.A1(_01094_),
    .A2(_01092_),
    .B1(_01091_),
    .C1(_01348_),
    .X(_01351_));
 sky130_fd_sc_hd__o32a_1 _09720_ (.A1(_03906_),
    .A2(_00270_),
    .A3(_00272_),
    .B1(_00428_),
    .B2(_02636_),
    .X(_01352_));
 sky130_fd_sc_hd__and4_1 _09721_ (.A(_02647_),
    .B(_03917_),
    .C(_00275_),
    .D(_00429_),
    .X(_01353_));
 sky130_fd_sc_hd__o32a_2 _09722_ (.A1(_04244_),
    .A2(_00145_),
    .A3(_00147_),
    .B1(_01352_),
    .B2(_01353_),
    .X(_01354_));
 sky130_fd_sc_hd__nor4_2 _09723_ (.A(_04244_),
    .B(net143),
    .C(_01352_),
    .D(_01353_),
    .Y(_01355_));
 sky130_fd_sc_hd__o21a_1 _09724_ (.A1(_01354_),
    .A2(_01355_),
    .B1(_01109_),
    .X(_01356_));
 sky130_fd_sc_hd__nor3_1 _09725_ (.A(_01354_),
    .B(_01355_),
    .C(_01109_),
    .Y(_01357_));
 sky130_fd_sc_hd__or2_1 _09726_ (.A(_01356_),
    .B(_01357_),
    .X(_01359_));
 sky130_fd_sc_hd__o31a_1 _09727_ (.A1(_03906_),
    .A2(net143),
    .A3(_01098_),
    .B1(_01097_),
    .X(_01360_));
 sky130_fd_sc_hd__o311a_1 _09728_ (.A1(_03906_),
    .A2(net143),
    .A3(_01098_),
    .B1(_01359_),
    .C1(_01097_),
    .X(_01361_));
 sky130_fd_sc_hd__nor2_1 _09729_ (.A(_01360_),
    .B(_01359_),
    .Y(_01362_));
 sky130_fd_sc_hd__o31a_1 _09730_ (.A1(_04244_),
    .A2(_00009_),
    .A3(_01110_),
    .B1(_01112_),
    .X(_01363_));
 sky130_fd_sc_hd__or3_2 _09731_ (.A(_01363_),
    .B(_01362_),
    .C(_01361_),
    .X(_01364_));
 sky130_fd_sc_hd__o21ai_2 _09732_ (.A1(_01361_),
    .A2(_01362_),
    .B1(_01363_),
    .Y(_01365_));
 sky130_fd_sc_hd__o211ai_1 _09733_ (.A1(_01116_),
    .A2(_01119_),
    .B1(_01123_),
    .C1(_00963_),
    .Y(_01366_));
 sky130_fd_sc_hd__o221ai_4 _09734_ (.A1(_00960_),
    .A2(_00964_),
    .B1(_01115_),
    .B2(_01118_),
    .C1(_01122_),
    .Y(_01367_));
 sky130_fd_sc_hd__a22o_1 _09735_ (.A1(_01364_),
    .A2(_01365_),
    .B1(_01367_),
    .B2(_01120_),
    .X(_01368_));
 sky130_fd_sc_hd__o2111ai_1 _09736_ (.A1(_01116_),
    .A2(_01119_),
    .B1(_01364_),
    .C1(_01365_),
    .D1(_01367_),
    .Y(_01370_));
 sky130_fd_sc_hd__o211a_2 _09737_ (.A1(_01350_),
    .A2(_01351_),
    .B1(_01368_),
    .C1(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__and2_2 _09738_ (.A(_01371_),
    .B(_01327_),
    .X(_01372_));
 sky130_fd_sc_hd__a211o_1 _09739_ (.A1(_01368_),
    .A2(_01370_),
    .B1(_01350_),
    .C1(_01351_),
    .X(_01373_));
 sky130_fd_sc_hd__nor2_1 _09740_ (.A(_01327_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_01327_),
    .B(_01373_),
    .Y(_01375_));
 sky130_fd_sc_hd__a21o_2 _09742_ (.A1(_01327_),
    .A2(_01373_),
    .B1(_01371_),
    .X(_01376_));
 sky130_fd_sc_hd__a21oi_2 _09743_ (.A1(_01327_),
    .A2(_01373_),
    .B1(_01371_),
    .Y(_01377_));
 sky130_fd_sc_hd__and2b_1 _09744_ (.A_N(_01371_),
    .B(_01373_),
    .X(_01378_));
 sky130_fd_sc_hd__o22ai_4 _09745_ (.A1(_01371_),
    .A2(_01375_),
    .B1(_01327_),
    .B2(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__o21ai_4 _09746_ (.A1(_01374_),
    .A2(_01376_),
    .B1(_01304_),
    .Y(_01381_));
 sky130_fd_sc_hd__o211a_1 _09747_ (.A1(_01126_),
    .A2(_01159_),
    .B1(_01129_),
    .C1(_01379_),
    .X(_01382_));
 sky130_fd_sc_hd__nor2_1 _09748_ (.A(_01304_),
    .B(_01379_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _09749_ (.A(_01382_),
    .B(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__o211ai_4 _09750_ (.A1(_00917_),
    .A2(_01017_),
    .B1(_01166_),
    .C1(_01168_),
    .Y(_01385_));
 sky130_fd_sc_hd__o211ai_4 _09751_ (.A1(_00918_),
    .A2(_01018_),
    .B1(_01165_),
    .C1(_01169_),
    .Y(_01386_));
 sky130_fd_sc_hd__o221ai_4 _09752_ (.A1(_01163_),
    .A2(_01164_),
    .B1(_01382_),
    .B2(_01383_),
    .C1(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__nand3_1 _09753_ (.A(_01165_),
    .B(_01385_),
    .C(_01384_),
    .Y(_01388_));
 sky130_fd_sc_hd__o211ai_1 _09754_ (.A1(_01382_),
    .A2(_01383_),
    .B1(_01385_),
    .C1(_01165_),
    .Y(_01389_));
 sky130_fd_sc_hd__o211ai_1 _09755_ (.A1(_01163_),
    .A2(_01164_),
    .B1(_01384_),
    .C1(_01386_),
    .Y(_01390_));
 sky130_fd_sc_hd__nand2_1 _09756_ (.A(_01387_),
    .B(_01388_),
    .Y(_01391_));
 sky130_fd_sc_hd__nand3b_2 _09757_ (.A_N(_01302_),
    .B(_01387_),
    .C(_01388_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand3_1 _09758_ (.A(_01389_),
    .B(_01390_),
    .C(_01302_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_4 _09759_ (.A(net10),
    .B(net11),
    .Y(_01394_));
 sky130_fd_sc_hd__or2_1 _09760_ (.A(net10),
    .B(net11),
    .X(_01395_));
 sky130_fd_sc_hd__and3_4 _09761_ (.A(_00564_),
    .B(_01052_),
    .C(_01394_),
    .X(_01396_));
 sky130_fd_sc_hd__nand4_4 _09762_ (.A(_00359_),
    .B(_00563_),
    .C(_01052_),
    .D(_01394_),
    .Y(_01397_));
 sky130_fd_sc_hd__a31oi_4 _09763_ (.A1(_00564_),
    .A2(_01052_),
    .A3(_01394_),
    .B1(_00321_),
    .Y(_01398_));
 sky130_fd_sc_hd__a21oi_4 _09764_ (.A1(_01397_),
    .A2(net174),
    .B1(net13),
    .Y(_01399_));
 sky130_fd_sc_hd__a21o_4 _09765_ (.A1(_01397_),
    .A2(net174),
    .B1(net13),
    .X(_01400_));
 sky130_fd_sc_hd__nor2_2 _09766_ (.A(_00321_),
    .B(_00671_),
    .Y(_01402_));
 sky130_fd_sc_hd__nand2_4 _09767_ (.A(net174),
    .B(net13),
    .Y(_01403_));
 sky130_fd_sc_hd__o311a_2 _09768_ (.A1(_01211_),
    .A2(net11),
    .A3(_00892_),
    .B1(net13),
    .C1(net174),
    .X(_01404_));
 sky130_fd_sc_hd__a21oi_4 _09769_ (.A1(_01397_),
    .A2(_01402_),
    .B1(_01399_),
    .Y(_01405_));
 sky130_fd_sc_hd__o21ai_4 _09770_ (.A1(_01396_),
    .A2(_01403_),
    .B1(_01400_),
    .Y(_01406_));
 sky130_fd_sc_hd__o211ai_4 _09771_ (.A1(_00856_),
    .A2(_00878_),
    .B1(net145),
    .C1(_01220_),
    .Y(_01407_));
 sky130_fd_sc_hd__o211ai_4 _09772_ (.A1(net170),
    .A2(_02057_),
    .B1(net147),
    .C1(net146),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_2 _09773_ (.A(_01226_),
    .B(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__o211ai_4 _09774_ (.A1(net170),
    .A2(_02057_),
    .B1(_00899_),
    .C1(_00902_),
    .Y(_01410_));
 sky130_fd_sc_hd__or4_1 _09775_ (.A(_02122_),
    .B(_00898_),
    .C(_00901_),
    .D(_01223_),
    .X(_01411_));
 sky130_fd_sc_hd__o21ai_2 _09776_ (.A1(_01223_),
    .A2(_01410_),
    .B1(_01409_),
    .Y(_01413_));
 sky130_fd_sc_hd__o2111ai_4 _09777_ (.A1(_01223_),
    .A2(_01410_),
    .B1(_01409_),
    .C1(_01303_),
    .D1(net141),
    .Y(_01414_));
 sky130_fd_sc_hd__o31a_1 _09778_ (.A1(_01292_),
    .A2(_01054_),
    .A3(_01056_),
    .B1(_01413_),
    .X(_01415_));
 sky130_fd_sc_hd__o21ai_1 _09779_ (.A1(_01292_),
    .A2(_01058_),
    .B1(_01413_),
    .Y(_01416_));
 sky130_fd_sc_hd__o211ai_1 _09780_ (.A1(_01238_),
    .A2(_01249_),
    .B1(net141),
    .C1(_01413_),
    .Y(_01417_));
 sky130_fd_sc_hd__o221ai_2 _09781_ (.A1(_01223_),
    .A2(_01410_),
    .B1(_01292_),
    .B2(_01058_),
    .C1(_01409_),
    .Y(_01418_));
 sky130_fd_sc_hd__o211ai_1 _09782_ (.A1(_00900_),
    .A2(_01221_),
    .B1(_01417_),
    .C1(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__o2111ai_2 _09783_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_01222_),
    .C1(_01414_),
    .D1(_01416_),
    .Y(_01420_));
 sky130_fd_sc_hd__o211ai_2 _09784_ (.A1(_00900_),
    .A2(_01221_),
    .B1(_01414_),
    .C1(_01416_),
    .Y(_01421_));
 sky130_fd_sc_hd__nand3b_1 _09785_ (.A_N(_01407_),
    .B(_01417_),
    .C(_01418_),
    .Y(_01422_));
 sky130_fd_sc_hd__and3_1 _09786_ (.A(_01419_),
    .B(_01420_),
    .C(_01228_),
    .X(_01424_));
 sky130_fd_sc_hd__nand3_2 _09787_ (.A(_01419_),
    .B(_01420_),
    .C(_01228_),
    .Y(_01425_));
 sky130_fd_sc_hd__o211ai_4 _09788_ (.A1(_01060_),
    .A2(_01226_),
    .B1(_01421_),
    .C1(_01422_),
    .Y(_01426_));
 sky130_fd_sc_hd__o2bb2ai_2 _09789_ (.A1_N(_01425_),
    .A2_N(_01426_),
    .B1(_00310_),
    .B2(_01406_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand4_1 _09790_ (.A(_01425_),
    .B(_01426_),
    .C(net33),
    .D(_01405_),
    .Y(_01428_));
 sky130_fd_sc_hd__o31a_1 _09791_ (.A1(_00310_),
    .A2(_01221_),
    .A3(_01229_),
    .B1(_01231_),
    .X(_01429_));
 sky130_fd_sc_hd__a21boi_2 _09792_ (.A1(_01427_),
    .A2(_01428_),
    .B1_N(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__a41oi_4 _09793_ (.A1(_01425_),
    .A2(_01426_),
    .A3(net33),
    .A4(_01405_),
    .B1(_01429_),
    .Y(_01431_));
 sky130_fd_sc_hd__a21oi_1 _09794_ (.A1(_01427_),
    .A2(_01431_),
    .B1(_01430_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _09795_ (.A(_01235_),
    .B(_01236_),
    .Y(_01433_));
 sky130_fd_sc_hd__a21bo_1 _09796_ (.A1(_01234_),
    .A2(_01237_),
    .B1_N(_01235_),
    .X(_01435_));
 sky130_fd_sc_hd__and2b_1 _09797_ (.A_N(_01432_),
    .B(_01435_),
    .X(_01436_));
 sky130_fd_sc_hd__a211oi_2 _09798_ (.A1(_01427_),
    .A2(_01431_),
    .B1(_01435_),
    .C1(_01430_),
    .Y(_01437_));
 sky130_fd_sc_hd__nor2_1 _09799_ (.A(_01436_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__nand3_1 _09800_ (.A(_01392_),
    .B(_01393_),
    .C(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__o2bb2ai_1 _09801_ (.A1_N(_01392_),
    .A2_N(_01393_),
    .B1(_01436_),
    .B2(_01437_),
    .Y(_01440_));
 sky130_fd_sc_hd__o211ai_1 _09802_ (.A1(_01436_),
    .A2(_01437_),
    .B1(_01392_),
    .C1(_01393_),
    .Y(_01441_));
 sky130_fd_sc_hd__a21bo_1 _09803_ (.A1(_01392_),
    .A2(_01393_),
    .B1_N(_01438_),
    .X(_01442_));
 sky130_fd_sc_hd__nand2_1 _09804_ (.A(_01441_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__a32o_1 _09805_ (.A1(_01170_),
    .A2(_01171_),
    .A3(_01208_),
    .B1(_01210_),
    .B2(_01243_),
    .X(_01444_));
 sky130_fd_sc_hd__a21o_1 _09806_ (.A1(_01439_),
    .A2(_01440_),
    .B1(_01444_),
    .X(_01446_));
 sky130_fd_sc_hd__nand3_2 _09807_ (.A(_01439_),
    .B(_01440_),
    .C(_01444_),
    .Y(_01447_));
 sky130_fd_sc_hd__o211ai_4 _09808_ (.A1(_00913_),
    .A2(_01076_),
    .B1(_01251_),
    .C1(_01075_),
    .Y(_01448_));
 sky130_fd_sc_hd__a22o_1 _09809_ (.A1(_01446_),
    .A2(_01447_),
    .B1(_01448_),
    .B2(_01252_),
    .X(_01449_));
 sky130_fd_sc_hd__o2111ai_4 _09810_ (.A1(_01248_),
    .A2(_01250_),
    .B1(_01446_),
    .C1(_01447_),
    .D1(_01448_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand2_1 _09811_ (.A(_01449_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__a2bb2o_1 _09812_ (.A1_N(_00834_),
    .A2_N(_01257_),
    .B1(_01449_),
    .B2(_01450_),
    .X(_01452_));
 sky130_fd_sc_hd__or3_1 _09813_ (.A(_00834_),
    .B(_01257_),
    .C(_01451_),
    .X(_01453_));
 sky130_fd_sc_hd__and2_1 _09814_ (.A(_01452_),
    .B(_01453_),
    .X(net77));
 sky130_fd_sc_hd__a2bb2o_1 _09815_ (.A1_N(_00812_),
    .A2_N(_00823_),
    .B1(_01257_),
    .B2(_01451_),
    .X(_01454_));
 sky130_fd_sc_hd__a311o_1 _09816_ (.A1(_01389_),
    .A2(_01390_),
    .A3(_01302_),
    .B1(_01436_),
    .C1(_01437_),
    .X(_01456_));
 sky130_fd_sc_hd__or3_1 _09817_ (.A(_04244_),
    .B(_00270_),
    .C(_00272_),
    .X(_01457_));
 sky130_fd_sc_hd__and3_1 _09818_ (.A(_03917_),
    .B(_00425_),
    .C(_00427_),
    .X(_01458_));
 sky130_fd_sc_hd__o32ai_1 _09819_ (.A1(_04244_),
    .A2(net143),
    .A3(_01352_),
    .B1(_00274_),
    .B2(_02636_),
    .Y(_01459_));
 sky130_fd_sc_hd__o32a_1 _09820_ (.A1(_04244_),
    .A2(net143),
    .A3(_01352_),
    .B1(_00428_),
    .B2(_03906_),
    .X(_01460_));
 sky130_fd_sc_hd__a31o_1 _09821_ (.A1(_03917_),
    .A2(_00429_),
    .A3(_01459_),
    .B1(_01460_),
    .X(_01461_));
 sky130_fd_sc_hd__xor2_2 _09822_ (.A(_01457_),
    .B(_01461_),
    .X(_01462_));
 sky130_fd_sc_hd__o32ai_4 _09823_ (.A1(_01109_),
    .A2(_01354_),
    .A3(_01355_),
    .B1(_01356_),
    .B2(_01360_),
    .Y(_01463_));
 sky130_fd_sc_hd__nor2_1 _09824_ (.A(_01462_),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_1 _09825_ (.A(_01462_),
    .B(_01463_),
    .X(_01465_));
 sky130_fd_sc_hd__nand2_1 _09826_ (.A(_01462_),
    .B(_01463_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _09827_ (.A(_01464_),
    .B(_01465_),
    .Y(_01468_));
 sky130_fd_sc_hd__o211ai_1 _09828_ (.A1(_01116_),
    .A2(_01119_),
    .B1(_01364_),
    .C1(_01367_),
    .Y(_01469_));
 sky130_fd_sc_hd__o211ai_2 _09829_ (.A1(_01115_),
    .A2(_01118_),
    .B1(_01365_),
    .C1(_01366_),
    .Y(_01470_));
 sky130_fd_sc_hd__o211ai_2 _09830_ (.A1(_01464_),
    .A2(_01465_),
    .B1(_01470_),
    .C1(_01364_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand3_1 _09831_ (.A(_01365_),
    .B(_01469_),
    .C(_01468_),
    .Y(_01472_));
 sky130_fd_sc_hd__a32o_1 _09832_ (.A1(_06341_),
    .A2(_00068_),
    .A3(_00070_),
    .B1(_07370_),
    .B2(_07540_),
    .X(_01473_));
 sky130_fd_sc_hd__nand4_2 _09833_ (.A(_06341_),
    .B(net151),
    .C(_07540_),
    .D(_00072_),
    .Y(_01474_));
 sky130_fd_sc_hd__nand4_1 _09834_ (.A(_00010_),
    .B(_05316_),
    .C(_07200_),
    .D(_00150_),
    .Y(_01475_));
 sky130_fd_sc_hd__a32o_1 _09835_ (.A1(_07200_),
    .A2(_00006_),
    .A3(_00008_),
    .B1(_00150_),
    .B2(_05316_),
    .X(_01476_));
 sky130_fd_sc_hd__o2bb2a_1 _09836_ (.A1_N(_01475_),
    .A2_N(_01476_),
    .B1(_07441_),
    .B2(_07512_),
    .X(_01478_));
 sky130_fd_sc_hd__a32o_1 _09837_ (.A1(_07436_),
    .A2(net154),
    .A3(_07513_),
    .B1(_01475_),
    .B2(_01476_),
    .X(_01479_));
 sky130_fd_sc_hd__and4_1 _09838_ (.A(_07513_),
    .B(_01475_),
    .C(_01476_),
    .D(_07440_),
    .X(_01480_));
 sky130_fd_sc_hd__o2111ai_1 _09839_ (.A1(_01331_),
    .A2(net143),
    .B1(_07513_),
    .C1(_07440_),
    .D1(_01476_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand4_1 _09840_ (.A(_01473_),
    .B(_01474_),
    .C(_01479_),
    .D(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__o2bb2a_1 _09841_ (.A1_N(_01473_),
    .A2_N(_01474_),
    .B1(_01478_),
    .B2(_01480_),
    .X(_01483_));
 sky130_fd_sc_hd__a22o_1 _09842_ (.A1(_01473_),
    .A2(_01474_),
    .B1(_01479_),
    .B2(_01481_),
    .X(_01484_));
 sky130_fd_sc_hd__or4bb_1 _09843_ (.A(_07512_),
    .B(_01331_),
    .C_N(_01482_),
    .D_N(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__a2bb2o_1 _09844_ (.A1_N(_01331_),
    .A2_N(_07512_),
    .B1(_01484_),
    .B2(_01482_),
    .X(_01486_));
 sky130_fd_sc_hd__o31a_1 _09845_ (.A1(_06331_),
    .A2(_07539_),
    .A3(_01333_),
    .B1(_01335_),
    .X(_01487_));
 sky130_fd_sc_hd__a21bo_1 _09846_ (.A1(_01485_),
    .A2(_01486_),
    .B1_N(_01487_),
    .X(_01489_));
 sky130_fd_sc_hd__nand3b_1 _09847_ (.A_N(_01487_),
    .B(_01486_),
    .C(_01485_),
    .Y(_01490_));
 sky130_fd_sc_hd__a2111oi_1 _09848_ (.A1(_01489_),
    .A2(_01490_),
    .B1(_05425_),
    .C1(_00188_),
    .D1(_00190_),
    .Y(_01491_));
 sky130_fd_sc_hd__o311a_1 _09849_ (.A1(_05425_),
    .A2(_00188_),
    .A3(_00190_),
    .B1(_01489_),
    .C1(_01490_),
    .X(_01492_));
 sky130_fd_sc_hd__a21bo_1 _09850_ (.A1(_01329_),
    .A2(_01340_),
    .B1_N(_01341_),
    .X(_01493_));
 sky130_fd_sc_hd__o21a_1 _09851_ (.A1(_01491_),
    .A2(_01492_),
    .B1(_01493_),
    .X(_01494_));
 sky130_fd_sc_hd__or3_1 _09852_ (.A(_01491_),
    .B(_01492_),
    .C(_01493_),
    .X(_01495_));
 sky130_fd_sc_hd__nand2b_1 _09853_ (.A_N(_01494_),
    .B(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__a21oi_1 _09854_ (.A1(_01345_),
    .A2(_01349_),
    .B1(_01346_),
    .Y(_01497_));
 sky130_fd_sc_hd__and2_1 _09855_ (.A(_01496_),
    .B(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__nor2_1 _09856_ (.A(_01496_),
    .B(_01497_),
    .Y(_01500_));
 sky130_fd_sc_hd__o211ai_2 _09857_ (.A1(_01498_),
    .A2(_01500_),
    .B1(_01471_),
    .C1(_01472_),
    .Y(_01501_));
 sky130_fd_sc_hd__a211o_1 _09858_ (.A1(_01471_),
    .A2(_01472_),
    .B1(_01498_),
    .C1(_01500_),
    .X(_01502_));
 sky130_fd_sc_hd__nand2_2 _09859_ (.A(_01501_),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__a32o_1 _09860_ (.A1(net156),
    .A2(_00189_),
    .A3(_00191_),
    .B1(_01308_),
    .B2(_01310_),
    .X(_01504_));
 sky130_fd_sc_hd__and3_1 _09861_ (.A(_04726_),
    .B(_00367_),
    .C(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__a32o_1 _09862_ (.A1(_04726_),
    .A2(_00362_),
    .A3(_00364_),
    .B1(_01308_),
    .B2(_01310_),
    .X(_01506_));
 sky130_fd_sc_hd__inv_2 _09863_ (.A(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__o32a_1 _09864_ (.A1(_03479_),
    .A2(_03522_),
    .A3(_00532_),
    .B1(_01505_),
    .B2(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__nor4_1 _09865_ (.A(_03544_),
    .B(_00532_),
    .C(_01505_),
    .D(_01507_),
    .Y(_01509_));
 sky130_fd_sc_hd__o21ai_1 _09866_ (.A1(_01508_),
    .A2(_01509_),
    .B1(_01317_),
    .Y(_01511_));
 sky130_fd_sc_hd__or3_1 _09867_ (.A(_01508_),
    .B(_01509_),
    .C(_01317_),
    .X(_01512_));
 sky130_fd_sc_hd__inv_2 _09868_ (.A(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_2 _09869_ (.A(_01511_),
    .B(_01512_),
    .Y(_01514_));
 sky130_fd_sc_hd__xor2_4 _09870_ (.A(_01326_),
    .B(_01514_),
    .X(_01515_));
 sky130_fd_sc_hd__xor2_4 _09871_ (.A(_01503_),
    .B(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__xnor2_2 _09872_ (.A(_01503_),
    .B(_01515_),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _09873_ (.A(_01377_),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__nand2_2 _09874_ (.A(_01376_),
    .B(_01516_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _09875_ (.A(_01518_),
    .B(_01519_),
    .Y(_01520_));
 sky130_fd_sc_hd__o211ai_4 _09876_ (.A1(_01381_),
    .A2(_01372_),
    .B1(_01165_),
    .C1(_01385_),
    .Y(_01522_));
 sky130_fd_sc_hd__o211ai_2 _09877_ (.A1(_01379_),
    .A2(_01304_),
    .B1(_01166_),
    .C1(_01386_),
    .Y(_01523_));
 sky130_fd_sc_hd__o211ai_1 _09878_ (.A1(_01304_),
    .A2(_01379_),
    .B1(_01520_),
    .C1(_01522_),
    .Y(_01524_));
 sky130_fd_sc_hd__o2111ai_1 _09879_ (.A1(_01372_),
    .A2(_01381_),
    .B1(_01518_),
    .C1(_01519_),
    .D1(_01523_),
    .Y(_01525_));
 sky130_fd_sc_hd__o2111ai_1 _09880_ (.A1(_01304_),
    .A2(_01379_),
    .B1(_01518_),
    .C1(_01519_),
    .D1(_01522_),
    .Y(_01526_));
 sky130_fd_sc_hd__o211ai_1 _09881_ (.A1(_01381_),
    .A2(_01372_),
    .B1(_01523_),
    .C1(_01520_),
    .Y(_01527_));
 sky130_fd_sc_hd__a21bo_1 _09882_ (.A1(_01261_),
    .A2(_01290_),
    .B1_N(_01289_),
    .X(_01528_));
 sky130_fd_sc_hd__and3_1 _09883_ (.A(_02647_),
    .B(_00577_),
    .C(_00579_),
    .X(_01529_));
 sky130_fd_sc_hd__and3_2 _09884_ (.A(_01262_),
    .B(_01038_),
    .C(_01969_),
    .X(_01530_));
 sky130_fd_sc_hd__o32a_2 _09885_ (.A1(_01488_),
    .A2(_01033_),
    .A3(_01035_),
    .B1(_01958_),
    .B2(_00744_),
    .X(_01531_));
 sky130_fd_sc_hd__a31oi_2 _09886_ (.A1(_01969_),
    .A2(_01038_),
    .A3(_01262_),
    .B1(_01531_),
    .Y(_01533_));
 sky130_fd_sc_hd__nor2_2 _09887_ (.A(net43),
    .B(net45),
    .Y(_01534_));
 sky130_fd_sc_hd__nand4b_4 _09888_ (.A_N(_00575_),
    .B(_01029_),
    .C(_01264_),
    .D(_00660_),
    .Y(_01535_));
 sky130_fd_sc_hd__o21ai_1 _09889_ (.A1(net45),
    .A2(_01265_),
    .B1(net173),
    .Y(_01536_));
 sky130_fd_sc_hd__nor2_4 _09890_ (.A(_00299_),
    .B(_00682_),
    .Y(_01537_));
 sky130_fd_sc_hd__o21a_4 _09891_ (.A1(net45),
    .A2(_01265_),
    .B1(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__o21ai_4 _09892_ (.A1(net45),
    .A2(_01265_),
    .B1(_01537_),
    .Y(_01539_));
 sky130_fd_sc_hd__a21oi_4 _09893_ (.A1(_01535_),
    .A2(net173),
    .B1(net46),
    .Y(_01540_));
 sky130_fd_sc_hd__a21o_4 _09894_ (.A1(_01535_),
    .A2(net173),
    .B1(net46),
    .X(_01541_));
 sky130_fd_sc_hd__nand2_8 _09895_ (.A(_01539_),
    .B(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__a21oi_4 _09896_ (.A1(_01535_),
    .A2(_01537_),
    .B1(_01540_),
    .Y(_01544_));
 sky130_fd_sc_hd__nand3_2 _09897_ (.A(_01541_),
    .B(net1),
    .C(_01539_),
    .Y(_01545_));
 sky130_fd_sc_hd__o31ai_4 _09898_ (.A1(_00288_),
    .A2(_01538_),
    .A3(_01540_),
    .B1(_01277_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand4_2 _09899_ (.A(_01273_),
    .B(_01539_),
    .C(_01541_),
    .D(_02177_),
    .Y(_01547_));
 sky130_fd_sc_hd__o221a_1 _09900_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01181_),
    .B2(_01182_),
    .C1(_01172_),
    .X(_01548_));
 sky130_fd_sc_hd__a22oi_4 _09901_ (.A1(net164),
    .A2(_01189_),
    .B1(_01546_),
    .B2(_01547_),
    .Y(_01549_));
 sky130_fd_sc_hd__a32o_1 _09902_ (.A1(net164),
    .A2(_01185_),
    .A3(_01187_),
    .B1(_01546_),
    .B2(_01547_),
    .X(_01550_));
 sky130_fd_sc_hd__o311a_1 _09903_ (.A1(_02188_),
    .A2(_01272_),
    .A3(_01542_),
    .B1(_01546_),
    .C1(_01548_),
    .X(_01551_));
 sky130_fd_sc_hd__nand4_1 _09904_ (.A(net164),
    .B(_01189_),
    .C(_01546_),
    .D(_01547_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand3_4 _09905_ (.A(_01550_),
    .B(_01552_),
    .C(_01533_),
    .Y(_01553_));
 sky130_fd_sc_hd__o22a_1 _09906_ (.A1(_01530_),
    .A2(_01531_),
    .B1(_01549_),
    .B2(_01551_),
    .X(_01555_));
 sky130_fd_sc_hd__o22ai_4 _09907_ (.A1(_01530_),
    .A2(_01531_),
    .B1(_01549_),
    .B2(_01551_),
    .Y(_01556_));
 sky130_fd_sc_hd__o2bb2ai_4 _09908_ (.A1_N(_01553_),
    .A2_N(_01556_),
    .B1(_01190_),
    .B2(_01277_),
    .Y(_01557_));
 sky130_fd_sc_hd__nand3b_4 _09909_ (.A_N(_01278_),
    .B(_01553_),
    .C(_01556_),
    .Y(_01558_));
 sky130_fd_sc_hd__o32a_1 _09910_ (.A1(net166),
    .A2(_01037_),
    .A3(_01279_),
    .B1(_01488_),
    .B2(_00744_),
    .X(_01559_));
 sky130_fd_sc_hd__and3_1 _09911_ (.A(_01499_),
    .B(_01284_),
    .C(_00743_),
    .X(_01560_));
 sky130_fd_sc_hd__a31o_1 _09912_ (.A1(_01499_),
    .A2(_01284_),
    .A3(_00743_),
    .B1(_01280_),
    .X(_01561_));
 sky130_fd_sc_hd__o211a_1 _09913_ (.A1(_01280_),
    .A2(_01560_),
    .B1(_01558_),
    .C1(_01557_),
    .X(_01562_));
 sky130_fd_sc_hd__o211ai_4 _09914_ (.A1(_01280_),
    .A2(_01560_),
    .B1(_01558_),
    .C1(_01557_),
    .Y(_01563_));
 sky130_fd_sc_hd__a21oi_2 _09915_ (.A1(_01557_),
    .A2(_01558_),
    .B1(_01561_),
    .Y(_01564_));
 sky130_fd_sc_hd__o2bb2ai_2 _09916_ (.A1_N(_01557_),
    .A2_N(_01558_),
    .B1(_01559_),
    .B2(_01283_),
    .Y(_01566_));
 sky130_fd_sc_hd__a21oi_2 _09917_ (.A1(_01563_),
    .A2(_01566_),
    .B1(_01529_),
    .Y(_01567_));
 sky130_fd_sc_hd__o22ai_1 _09918_ (.A1(_02636_),
    .A2(_00580_),
    .B1(_01562_),
    .B2(_01564_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand3_1 _09919_ (.A(_01566_),
    .B(_01529_),
    .C(_01563_),
    .Y(_01569_));
 sky130_fd_sc_hd__a21boi_1 _09920_ (.A1(_01563_),
    .A2(_01566_),
    .B1_N(_01529_),
    .Y(_01570_));
 sky130_fd_sc_hd__o311a_1 _09921_ (.A1(_02636_),
    .A2(_00576_),
    .A3(_00578_),
    .B1(_01563_),
    .C1(_01566_),
    .X(_01571_));
 sky130_fd_sc_hd__nand2_1 _09922_ (.A(_01569_),
    .B(_01528_),
    .Y(_01572_));
 sky130_fd_sc_hd__a21oi_1 _09923_ (.A1(_01568_),
    .A2(_01569_),
    .B1(_01528_),
    .Y(_01573_));
 sky130_fd_sc_hd__o21ba_2 _09924_ (.A1(_01567_),
    .A2(_01572_),
    .B1_N(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__xor2_1 _09925_ (.A(_01301_),
    .B(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__xnor2_1 _09926_ (.A(_01301_),
    .B(_01574_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand3_1 _09927_ (.A(_01524_),
    .B(_01525_),
    .C(_01575_),
    .Y(_01578_));
 sky130_fd_sc_hd__nand3_1 _09928_ (.A(_01526_),
    .B(_01527_),
    .C(_01577_),
    .Y(_01579_));
 sky130_fd_sc_hd__a31o_1 _09929_ (.A1(net33),
    .A2(_01405_),
    .A3(_01426_),
    .B1(_01424_),
    .X(_01580_));
 sky130_fd_sc_hd__nor4_4 _09930_ (.A(net9),
    .B(_01395_),
    .C(net13),
    .D(_00892_),
    .Y(_01581_));
 sky130_fd_sc_hd__nand4_4 _09931_ (.A(_00564_),
    .B(_01052_),
    .C(_01394_),
    .D(_00671_),
    .Y(_01582_));
 sky130_fd_sc_hd__a41o_1 _09932_ (.A1(_00564_),
    .A2(_01052_),
    .A3(_01394_),
    .A4(_00671_),
    .B1(_00321_),
    .X(_01583_));
 sky130_fd_sc_hd__o311a_4 _09933_ (.A1(_01395_),
    .A2(net13),
    .A3(_01053_),
    .B1(net14),
    .C1(net174),
    .X(_01584_));
 sky130_fd_sc_hd__o211ai_4 _09934_ (.A1(net13),
    .A2(_01397_),
    .B1(net14),
    .C1(net174),
    .Y(_01585_));
 sky130_fd_sc_hd__a21oi_4 _09935_ (.A1(_01582_),
    .A2(net174),
    .B1(net14),
    .Y(_01586_));
 sky130_fd_sc_hd__a21o_4 _09936_ (.A1(_01582_),
    .A2(net174),
    .B1(net14),
    .X(_01588_));
 sky130_fd_sc_hd__nand2_8 _09937_ (.A(_01585_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_8 _09938_ (.A(_01584_),
    .B(_01586_),
    .Y(_01590_));
 sky130_fd_sc_hd__and3_1 _09939_ (.A(_01588_),
    .B(net33),
    .C(_01585_),
    .X(_01591_));
 sky130_fd_sc_hd__o32a_1 _09940_ (.A1(_01292_),
    .A2(_01058_),
    .A3(_01413_),
    .B1(_01221_),
    .B2(_00900_),
    .X(_01592_));
 sky130_fd_sc_hd__o21ai_1 _09941_ (.A1(_01407_),
    .A2(_01415_),
    .B1(_01414_),
    .Y(_01593_));
 sky130_fd_sc_hd__o211ai_2 _09942_ (.A1(_01238_),
    .A2(_01249_),
    .B1(net145),
    .C1(_01220_),
    .Y(_01594_));
 sky130_fd_sc_hd__a21oi_2 _09943_ (.A1(_01397_),
    .A2(_01402_),
    .B1(_00900_),
    .Y(_01595_));
 sky130_fd_sc_hd__o21ai_4 _09944_ (.A1(net13),
    .A2(_01398_),
    .B1(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__nand2_1 _09945_ (.A(_01594_),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__o221ai_4 _09946_ (.A1(_01238_),
    .A2(_01249_),
    .B1(_01396_),
    .B2(_01403_),
    .C1(_01400_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand4_2 _09947_ (.A(_01222_),
    .B(_01595_),
    .C(_01400_),
    .D(_01303_),
    .Y(_01600_));
 sky130_fd_sc_hd__o21ai_1 _09948_ (.A1(_01407_),
    .A2(_01599_),
    .B1(_01597_),
    .Y(_01601_));
 sky130_fd_sc_hd__o211ai_4 _09949_ (.A1(net168),
    .A2(net163),
    .B1(_00899_),
    .C1(_00902_),
    .Y(_01602_));
 sky130_fd_sc_hd__a211o_2 _09950_ (.A1(_00895_),
    .A2(_00897_),
    .B1(net159),
    .C1(_01408_),
    .X(_01603_));
 sky130_fd_sc_hd__o211ai_4 _09951_ (.A1(_02790_),
    .A2(net163),
    .B1(net147),
    .C1(net146),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_2 _09952_ (.A(_01410_),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__o2bb2ai_1 _09953_ (.A1_N(_01410_),
    .A2_N(_01604_),
    .B1(_01602_),
    .B2(_01408_),
    .Y(_01606_));
 sky130_fd_sc_hd__o21ai_1 _09954_ (.A1(_01620_),
    .A2(_01058_),
    .B1(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__o2111ai_4 _09955_ (.A1(_01408_),
    .A2(_01602_),
    .B1(_01605_),
    .C1(net141),
    .D1(_01631_),
    .Y(_01608_));
 sky130_fd_sc_hd__o211ai_2 _09956_ (.A1(_01532_),
    .A2(_01554_),
    .B1(net141),
    .C1(_01606_),
    .Y(_01610_));
 sky130_fd_sc_hd__o221ai_4 _09957_ (.A1(_01408_),
    .A2(_01602_),
    .B1(_01620_),
    .B2(_01058_),
    .C1(_01605_),
    .Y(_01611_));
 sky130_fd_sc_hd__o2111ai_4 _09958_ (.A1(_01407_),
    .A2(_01599_),
    .B1(_01607_),
    .C1(_01608_),
    .D1(_01597_),
    .Y(_01612_));
 sky130_fd_sc_hd__nand3_4 _09959_ (.A(_01601_),
    .B(_01610_),
    .C(_01611_),
    .Y(_01613_));
 sky130_fd_sc_hd__o211ai_2 _09960_ (.A1(_01226_),
    .A2(_01408_),
    .B1(_01612_),
    .C1(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__a21o_1 _09961_ (.A1(_01612_),
    .A2(_01613_),
    .B1(_01411_),
    .X(_01615_));
 sky130_fd_sc_hd__nand3b_1 _09962_ (.A_N(_01411_),
    .B(_01612_),
    .C(_01613_),
    .Y(_01616_));
 sky130_fd_sc_hd__o2bb2ai_1 _09963_ (.A1_N(_01612_),
    .A2_N(_01613_),
    .B1(_01226_),
    .B2(_01408_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand3_1 _09964_ (.A(_01617_),
    .B(_01593_),
    .C(_01616_),
    .Y(_01618_));
 sky130_fd_sc_hd__o211ai_2 _09965_ (.A1(_01415_),
    .A2(_01592_),
    .B1(_01614_),
    .C1(_01615_),
    .Y(_01619_));
 sky130_fd_sc_hd__nand3_1 _09966_ (.A(_01615_),
    .B(_01593_),
    .C(_01614_),
    .Y(_01621_));
 sky130_fd_sc_hd__o211ai_1 _09967_ (.A1(_01415_),
    .A2(_01592_),
    .B1(_01616_),
    .C1(_01617_),
    .Y(_01622_));
 sky130_fd_sc_hd__o211ai_1 _09968_ (.A1(_01589_),
    .A2(_00310_),
    .B1(_01622_),
    .C1(_01621_),
    .Y(_01623_));
 sky130_fd_sc_hd__nand3_1 _09969_ (.A(_01619_),
    .B(_01591_),
    .C(_01618_),
    .Y(_01624_));
 sky130_fd_sc_hd__o211ai_1 _09970_ (.A1(_00310_),
    .A2(_01589_),
    .B1(_01618_),
    .C1(_01619_),
    .Y(_01625_));
 sky130_fd_sc_hd__nand4_1 _09971_ (.A(_01621_),
    .B(net33),
    .C(_01590_),
    .D(_01622_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _09972_ (.A(_01625_),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__nand3_1 _09973_ (.A(_01623_),
    .B(_01624_),
    .C(_01580_),
    .Y(_01628_));
 sky130_fd_sc_hd__a311o_1 _09974_ (.A1(net33),
    .A2(_01426_),
    .A3(_01405_),
    .B1(_01424_),
    .C1(_01627_),
    .X(_01629_));
 sky130_fd_sc_hd__nand2_1 _09975_ (.A(_01628_),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__a22oi_2 _09976_ (.A1(_01234_),
    .A2(_01433_),
    .B1(_01431_),
    .B2(_01427_),
    .Y(_01632_));
 sky130_fd_sc_hd__o2bb2a_1 _09977_ (.A1_N(_01628_),
    .A2_N(_01629_),
    .B1(_01632_),
    .B2(_01430_),
    .X(_01633_));
 sky130_fd_sc_hd__nor3_1 _09978_ (.A(_01430_),
    .B(_01632_),
    .C(_01630_),
    .Y(_01634_));
 sky130_fd_sc_hd__or2_1 _09979_ (.A(_01633_),
    .B(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__nand3b_1 _09980_ (.A_N(_01635_),
    .B(_01579_),
    .C(_01578_),
    .Y(_01636_));
 sky130_fd_sc_hd__o2bb2ai_1 _09981_ (.A1_N(_01578_),
    .A2_N(_01579_),
    .B1(_01633_),
    .B2(_01634_),
    .Y(_01637_));
 sky130_fd_sc_hd__o2111ai_2 _09982_ (.A1(_01302_),
    .A2(_01391_),
    .B1(_01456_),
    .C1(_01636_),
    .D1(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__a22o_1 _09983_ (.A1(_01392_),
    .A2(_01456_),
    .B1(_01636_),
    .B2(_01637_),
    .X(_01639_));
 sky130_fd_sc_hd__nand2_1 _09984_ (.A(_01638_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__o211ai_2 _09985_ (.A1(_01248_),
    .A2(_01250_),
    .B1(_01447_),
    .C1(_01448_),
    .Y(_01641_));
 sky130_fd_sc_hd__o21ai_2 _09986_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_01641_),
    .Y(_01643_));
 sky130_fd_sc_hd__xnor2_2 _09987_ (.A(_01640_),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__xnor2_1 _09988_ (.A(_01454_),
    .B(_01644_),
    .Y(net78));
 sky130_fd_sc_hd__a2111oi_4 _09989_ (.A1(_01449_),
    .A2(_01450_),
    .B1(_01644_),
    .C1(_01254_),
    .D1(_01079_),
    .Y(_01645_));
 sky130_fd_sc_hd__a32o_1 _09990_ (.A1(_01524_),
    .A2(_01525_),
    .A3(_01575_),
    .B1(_01579_),
    .B2(_01635_),
    .X(_01646_));
 sky130_fd_sc_hd__a31o_1 _09991_ (.A1(_01544_),
    .A2(_02177_),
    .A3(_01273_),
    .B1(_01548_),
    .X(_01647_));
 sky130_fd_sc_hd__a21oi_2 _09992_ (.A1(_01546_),
    .A2(_01647_),
    .B1(_01530_),
    .Y(_01648_));
 sky130_fd_sc_hd__and3_1 _09993_ (.A(_01647_),
    .B(_01530_),
    .C(_01546_),
    .X(_01649_));
 sky130_fd_sc_hd__nand3_2 _09994_ (.A(_01647_),
    .B(_01530_),
    .C(_01546_),
    .Y(_01650_));
 sky130_fd_sc_hd__and3_2 _09995_ (.A(_01499_),
    .B(_01185_),
    .C(_01187_),
    .X(_01651_));
 sky130_fd_sc_hd__or3_1 _09996_ (.A(_01488_),
    .B(_01184_),
    .C(_01186_),
    .X(_01653_));
 sky130_fd_sc_hd__o2bb2ai_2 _09997_ (.A1_N(_01537_),
    .A2_N(_01535_),
    .B1(_00943_),
    .B2(net172),
    .Y(_01654_));
 sky130_fd_sc_hd__a21oi_1 _09998_ (.A1(_00682_),
    .A2(_01536_),
    .B1(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand4_4 _09999_ (.A(_00738_),
    .B(_01178_),
    .C(_01534_),
    .D(_00682_),
    .Y(_01656_));
 sky130_fd_sc_hd__a41o_1 _10000_ (.A1(_00738_),
    .A2(_01178_),
    .A3(_01534_),
    .A4(_00682_),
    .B1(_00299_),
    .X(_01657_));
 sky130_fd_sc_hd__a21oi_4 _10001_ (.A1(_01656_),
    .A2(net173),
    .B1(net47),
    .Y(_01658_));
 sky130_fd_sc_hd__a21o_4 _10002_ (.A1(_01656_),
    .A2(net173),
    .B1(net47),
    .X(_01659_));
 sky130_fd_sc_hd__o311a_4 _10003_ (.A1(net45),
    .A2(net46),
    .A3(_01265_),
    .B1(net47),
    .C1(net173),
    .X(_01660_));
 sky130_fd_sc_hd__o211ai_4 _10004_ (.A1(net46),
    .A2(_01535_),
    .B1(net47),
    .C1(net173),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_8 _10005_ (.A(_01659_),
    .B(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__nor2_8 _10006_ (.A(_01658_),
    .B(_01660_),
    .Y(_01664_));
 sky130_fd_sc_hd__nand3_2 _10007_ (.A(_01659_),
    .B(net140),
    .C(net1),
    .Y(_01665_));
 sky130_fd_sc_hd__o21ai_4 _10008_ (.A1(_01540_),
    .A2(_01654_),
    .B1(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__o211ai_4 _10009_ (.A1(_00921_),
    .A2(_00943_),
    .B1(_01659_),
    .C1(net140),
    .Y(_01667_));
 sky130_fd_sc_hd__and3_1 _10010_ (.A(_01664_),
    .B(_01655_),
    .C(net1),
    .X(_01668_));
 sky130_fd_sc_hd__nand4_4 _10011_ (.A(net1),
    .B(_01655_),
    .C(_01659_),
    .D(net140),
    .Y(_01669_));
 sky130_fd_sc_hd__and3_1 _10012_ (.A(net164),
    .B(_01269_),
    .C(_01271_),
    .X(_01670_));
 sky130_fd_sc_hd__a22oi_4 _10013_ (.A1(net164),
    .A2(_01273_),
    .B1(_01666_),
    .B2(_01669_),
    .Y(_01671_));
 sky130_fd_sc_hd__a32o_2 _10014_ (.A1(net164),
    .A2(_01269_),
    .A3(_01271_),
    .B1(_01666_),
    .B2(_01669_),
    .X(_01672_));
 sky130_fd_sc_hd__o311a_1 _10015_ (.A1(_00987_),
    .A2(_01545_),
    .A3(_01662_),
    .B1(_01670_),
    .C1(_01666_),
    .X(_01673_));
 sky130_fd_sc_hd__o2111ai_4 _10016_ (.A1(_01545_),
    .A2(_01667_),
    .B1(_01666_),
    .C1(net164),
    .D1(_01273_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand3_1 _10017_ (.A(_01672_),
    .B(_01675_),
    .C(_01651_),
    .Y(_01676_));
 sky130_fd_sc_hd__o22ai_2 _10018_ (.A1(_01488_),
    .A2(_01188_),
    .B1(_01671_),
    .B2(_01673_),
    .Y(_01677_));
 sky130_fd_sc_hd__o21ai_2 _10019_ (.A1(_01671_),
    .A2(_01673_),
    .B1(_01651_),
    .Y(_01678_));
 sky130_fd_sc_hd__o211ai_4 _10020_ (.A1(_01488_),
    .A2(_01188_),
    .B1(_01672_),
    .C1(_01675_),
    .Y(_01679_));
 sky130_fd_sc_hd__o211ai_4 _10021_ (.A1(_01648_),
    .A2(_01649_),
    .B1(_01678_),
    .C1(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__nand4b_4 _10022_ (.A_N(_01648_),
    .B(_01650_),
    .C(_01676_),
    .D(_01677_),
    .Y(_01681_));
 sky130_fd_sc_hd__o31a_1 _10023_ (.A1(_00288_),
    .A2(_01192_),
    .A3(_01272_),
    .B1(_01553_),
    .X(_01682_));
 sky130_fd_sc_hd__o21ai_2 _10024_ (.A1(_01190_),
    .A2(_01277_),
    .B1(_01553_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand4_4 _10025_ (.A(_01556_),
    .B(_01680_),
    .C(_01681_),
    .D(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__inv_2 _10026_ (.A(_01684_),
    .Y(_01686_));
 sky130_fd_sc_hd__o2bb2ai_4 _10027_ (.A1_N(_01680_),
    .A2_N(_01681_),
    .B1(_01682_),
    .B2(_01555_),
    .Y(_01687_));
 sky130_fd_sc_hd__nor4_4 _10028_ (.A(_01958_),
    .B(_02636_),
    .C(_00744_),
    .D(_01037_),
    .Y(_01688_));
 sky130_fd_sc_hd__o32a_4 _10029_ (.A1(_01958_),
    .A2(_01033_),
    .A3(_01035_),
    .B1(_02636_),
    .B2(_00744_),
    .X(_01689_));
 sky130_fd_sc_hd__o32a_1 _10030_ (.A1(_03906_),
    .A2(_00576_),
    .A3(_00578_),
    .B1(_01688_),
    .B2(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__nor4_1 _10031_ (.A(_03906_),
    .B(_00580_),
    .C(_01688_),
    .D(_01689_),
    .Y(_01691_));
 sky130_fd_sc_hd__o211a_1 _10032_ (.A1(_01688_),
    .A2(_01689_),
    .B1(_03917_),
    .C1(_00581_),
    .X(_01692_));
 sky130_fd_sc_hd__a311oi_4 _10033_ (.A1(_03917_),
    .A2(_00577_),
    .A3(_00579_),
    .B1(_01688_),
    .C1(_01689_),
    .Y(_01693_));
 sky130_fd_sc_hd__o2bb2ai_4 _10034_ (.A1_N(_01684_),
    .A2_N(_01687_),
    .B1(_01692_),
    .B2(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__o211ai_4 _10035_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01684_),
    .C1(_01687_),
    .Y(_01695_));
 sky130_fd_sc_hd__and2_1 _10036_ (.A(_01694_),
    .B(_01695_),
    .X(_01697_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(_01694_),
    .B(_01695_),
    .Y(_01698_));
 sky130_fd_sc_hd__o31a_1 _10038_ (.A1(_02636_),
    .A2(_00576_),
    .A3(_00578_),
    .B1(_01563_),
    .X(_01699_));
 sky130_fd_sc_hd__a211oi_2 _10039_ (.A1(_02592_),
    .A2(_02603_),
    .B1(_00580_),
    .C1(_01564_),
    .Y(_01700_));
 sky130_fd_sc_hd__o31a_1 _10040_ (.A1(_02636_),
    .A2(_00580_),
    .A3(_01564_),
    .B1(_01563_),
    .X(_01701_));
 sky130_fd_sc_hd__inv_2 _10041_ (.A(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__o2bb2ai_4 _10042_ (.A1_N(_01694_),
    .A2_N(_01695_),
    .B1(_01700_),
    .B2(_01562_),
    .Y(_01703_));
 sky130_fd_sc_hd__o211ai_4 _10043_ (.A1(_01564_),
    .A2(_01699_),
    .B1(_01695_),
    .C1(_01694_),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_2 _10044_ (.A(_01703_),
    .B(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__o22ai_2 _10045_ (.A1(_01297_),
    .A2(_01300_),
    .B1(_01567_),
    .B2(_01572_),
    .Y(_01706_));
 sky130_fd_sc_hd__o22a_1 _10046_ (.A1(_01567_),
    .A2(_01572_),
    .B1(_01301_),
    .B2(_01573_),
    .X(_01708_));
 sky130_fd_sc_hd__xor2_4 _10047_ (.A(_01705_),
    .B(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__a31o_1 _10048_ (.A1(net156),
    .A2(_00533_),
    .A3(_01506_),
    .B1(_01505_),
    .X(_01710_));
 sky130_fd_sc_hd__and3_1 _10049_ (.A(_04726_),
    .B(_00533_),
    .C(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__a31o_1 _10050_ (.A1(_04682_),
    .A2(_04704_),
    .A3(_00533_),
    .B1(_01710_),
    .X(_01712_));
 sky130_fd_sc_hd__and2b_1 _10051_ (.A_N(_01711_),
    .B(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__a31o_2 _10052_ (.A1(_01321_),
    .A2(_01324_),
    .A3(_01511_),
    .B1(_01513_),
    .X(_01714_));
 sky130_fd_sc_hd__xor2_4 _10053_ (.A(_01713_),
    .B(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__o21ai_1 _10054_ (.A1(_05425_),
    .A2(_00192_),
    .B1(_01490_),
    .Y(_01716_));
 sky130_fd_sc_hd__nand2_1 _10055_ (.A(_01489_),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__a2bb2o_1 _10056_ (.A1_N(net143),
    .A2_N(_01331_),
    .B1(_07440_),
    .B2(_07513_),
    .X(_01719_));
 sky130_fd_sc_hd__a21bo_1 _10057_ (.A1(_01476_),
    .A2(_01719_),
    .B1_N(_01474_),
    .X(_01720_));
 sky130_fd_sc_hd__nand3b_1 _10058_ (.A_N(_01474_),
    .B(_01476_),
    .C(_01719_),
    .Y(_01721_));
 sky130_fd_sc_hd__nand2_1 _10059_ (.A(_01720_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__a32o_1 _10060_ (.A1(_05316_),
    .A2(_00271_),
    .A3(_00273_),
    .B1(_07200_),
    .B2(_00150_),
    .X(_01723_));
 sky130_fd_sc_hd__nand4_1 _10061_ (.A(_00271_),
    .B(_05316_),
    .C(_07200_),
    .D(_00273_),
    .Y(_01724_));
 sky130_fd_sc_hd__and4_1 _10062_ (.A(_07200_),
    .B(_00150_),
    .C(_00275_),
    .D(_05316_),
    .X(_01725_));
 sky130_fd_sc_hd__nand4_2 _10063_ (.A(_07200_),
    .B(_00150_),
    .C(_00275_),
    .D(_05316_),
    .Y(_01726_));
 sky130_fd_sc_hd__o2111a_1 _10064_ (.A1(_01724_),
    .A2(net143),
    .B1(_00010_),
    .C1(_07440_),
    .D1(_01723_),
    .X(_01727_));
 sky130_fd_sc_hd__o2111ai_1 _10065_ (.A1(_01724_),
    .A2(net143),
    .B1(_00010_),
    .C1(_07440_),
    .D1(_01723_),
    .Y(_01728_));
 sky130_fd_sc_hd__a22oi_1 _10066_ (.A1(_07440_),
    .A2(_00010_),
    .B1(_01723_),
    .B2(_01726_),
    .Y(_01730_));
 sky130_fd_sc_hd__a32o_1 _10067_ (.A1(_07436_),
    .A2(net154),
    .A3(_00010_),
    .B1(_01723_),
    .B2(_01726_),
    .X(_01731_));
 sky130_fd_sc_hd__o22ai_1 _10068_ (.A1(_07512_),
    .A2(_07539_),
    .B1(_01727_),
    .B2(_01730_),
    .Y(_01732_));
 sky130_fd_sc_hd__o2111ai_1 _10069_ (.A1(_07506_),
    .A2(_07507_),
    .B1(_07540_),
    .C1(_01728_),
    .D1(_01731_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand2_1 _10070_ (.A(_01732_),
    .B(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__xnor2_1 _10071_ (.A(_01722_),
    .B(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__o31a_1 _10072_ (.A1(_07512_),
    .A2(_01331_),
    .A3(_01483_),
    .B1(_01482_),
    .X(_01736_));
 sky130_fd_sc_hd__xor2_1 _10073_ (.A(_01735_),
    .B(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__and4_1 _10074_ (.A(_06341_),
    .B(net151),
    .C(_00072_),
    .D(_00193_),
    .X(_01738_));
 sky130_fd_sc_hd__or4_1 _10075_ (.A(_06331_),
    .B(net153),
    .C(net148),
    .D(_00192_),
    .X(_01739_));
 sky130_fd_sc_hd__a32o_1 _10076_ (.A1(_06341_),
    .A2(_00189_),
    .A3(_00191_),
    .B1(net151),
    .B2(_00072_),
    .X(_01741_));
 sky130_fd_sc_hd__a32o_1 _10077_ (.A1(_05436_),
    .A2(_00362_),
    .A3(_00364_),
    .B1(_01739_),
    .B2(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__or4b_1 _10078_ (.A(_05425_),
    .B(_00366_),
    .C(_01738_),
    .D_N(_01741_),
    .X(_01743_));
 sky130_fd_sc_hd__nand2_1 _10079_ (.A(_01742_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__xnor2_1 _10080_ (.A(_01737_),
    .B(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__nand3_1 _10081_ (.A(_01745_),
    .B(_01716_),
    .C(_01489_),
    .Y(_01746_));
 sky130_fd_sc_hd__a21oi_1 _10082_ (.A1(_01489_),
    .A2(_01716_),
    .B1(_01745_),
    .Y(_01747_));
 sky130_fd_sc_hd__xnor2_1 _10083_ (.A(_01717_),
    .B(_01745_),
    .Y(_01748_));
 sky130_fd_sc_hd__a21oi_1 _10084_ (.A1(_01495_),
    .A2(_01497_),
    .B1(_01494_),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_1 _10085_ (.A(_01749_),
    .B(_01748_),
    .Y(_01750_));
 sky130_fd_sc_hd__and2_1 _10086_ (.A(_01748_),
    .B(_01749_),
    .X(_01752_));
 sky130_fd_sc_hd__a2bb2o_1 _10087_ (.A1_N(_01457_),
    .A2_N(_01460_),
    .B1(_01458_),
    .B2(_01459_),
    .X(_01753_));
 sky130_fd_sc_hd__a31o_1 _10088_ (.A1(_04222_),
    .A2(_04233_),
    .A3(_00429_),
    .B1(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__or3b_1 _10089_ (.A(_04244_),
    .B(_00428_),
    .C_N(_01753_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _10090_ (.A(_01754_),
    .B(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__nand3_1 _10091_ (.A(_01364_),
    .B(_01467_),
    .C(_01470_),
    .Y(_01757_));
 sky130_fd_sc_hd__o211ai_1 _10092_ (.A1(_01462_),
    .A2(_01463_),
    .B1(_01469_),
    .C1(_01365_),
    .Y(_01758_));
 sky130_fd_sc_hd__o211ai_2 _10093_ (.A1(_01462_),
    .A2(_01463_),
    .B1(_01756_),
    .C1(_01757_),
    .Y(_01759_));
 sky130_fd_sc_hd__nand4_1 _10094_ (.A(_01467_),
    .B(_01754_),
    .C(_01755_),
    .D(_01758_),
    .Y(_01760_));
 sky130_fd_sc_hd__and4bb_1 _10095_ (.A_N(_01750_),
    .B_N(_01752_),
    .C(_01759_),
    .D(_01760_),
    .X(_01761_));
 sky130_fd_sc_hd__a2bb2oi_2 _10096_ (.A1_N(_01750_),
    .A2_N(_01752_),
    .B1(_01759_),
    .B2(_01760_),
    .Y(_01763_));
 sky130_fd_sc_hd__or2_1 _10097_ (.A(_01715_),
    .B(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__o21ai_1 _10098_ (.A1(_01761_),
    .A2(_01763_),
    .B1(_01715_),
    .Y(_01765_));
 sky130_fd_sc_hd__o21a_2 _10099_ (.A1(_01761_),
    .A2(_01764_),
    .B1(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__nand2_1 _10100_ (.A(_01502_),
    .B(_01515_),
    .Y(_01767_));
 sky130_fd_sc_hd__and2_2 _10101_ (.A(_01501_),
    .B(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__a21o_1 _10102_ (.A1(_01501_),
    .A2(_01767_),
    .B1(_01766_),
    .X(_01769_));
 sky130_fd_sc_hd__nand2_2 _10103_ (.A(_01766_),
    .B(_01768_),
    .Y(_01770_));
 sky130_fd_sc_hd__and2_1 _10104_ (.A(_01769_),
    .B(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__nand2_1 _10105_ (.A(_01769_),
    .B(_01770_),
    .Y(_01772_));
 sky130_fd_sc_hd__o211ai_4 _10106_ (.A1(_01304_),
    .A2(_01379_),
    .B1(_01519_),
    .C1(_01522_),
    .Y(_01774_));
 sky130_fd_sc_hd__o211ai_2 _10107_ (.A1(_01372_),
    .A2(_01381_),
    .B1(_01518_),
    .C1(_01523_),
    .Y(_01775_));
 sky130_fd_sc_hd__o211ai_1 _10108_ (.A1(_01377_),
    .A2(_01517_),
    .B1(_01772_),
    .C1(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__o211ai_1 _10109_ (.A1(_01376_),
    .A2(_01516_),
    .B1(_01771_),
    .C1(_01774_),
    .Y(_01777_));
 sky130_fd_sc_hd__o2111ai_1 _10110_ (.A1(_01377_),
    .A2(_01517_),
    .B1(_01769_),
    .C1(_01770_),
    .D1(_01775_),
    .Y(_01778_));
 sky130_fd_sc_hd__o211ai_1 _10111_ (.A1(_01376_),
    .A2(_01516_),
    .B1(_01772_),
    .C1(_01774_),
    .Y(_01779_));
 sky130_fd_sc_hd__nand3b_2 _10112_ (.A_N(_01709_),
    .B(_01776_),
    .C(_01777_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand3_2 _10113_ (.A(_01778_),
    .B(_01779_),
    .C(_01709_),
    .Y(_01781_));
 sky130_fd_sc_hd__inv_2 _10114_ (.A(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__o21ai_2 _10115_ (.A1(_01226_),
    .A2(_01408_),
    .B1(_01612_),
    .Y(_01783_));
 sky130_fd_sc_hd__nand2_1 _10116_ (.A(_01613_),
    .B(_01783_),
    .Y(_01785_));
 sky130_fd_sc_hd__o2111ai_4 _10117_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_01055_),
    .C1(_01057_),
    .D1(_01605_),
    .Y(_01786_));
 sky130_fd_sc_hd__o211a_1 _10118_ (.A1(_01594_),
    .A2(_01596_),
    .B1(_01603_),
    .C1(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__o211ai_2 _10119_ (.A1(_01594_),
    .A2(_01596_),
    .B1(_01603_),
    .C1(_01786_),
    .Y(_01788_));
 sky130_fd_sc_hd__a21oi_4 _10120_ (.A1(_01603_),
    .A2(_01786_),
    .B1(_01600_),
    .Y(_01789_));
 sky130_fd_sc_hd__a21o_1 _10121_ (.A1(_01603_),
    .A2(_01786_),
    .B1(_01600_),
    .X(_01790_));
 sky130_fd_sc_hd__o211ai_4 _10122_ (.A1(_01532_),
    .A2(_01554_),
    .B1(net145),
    .C1(_01220_),
    .Y(_01791_));
 sky130_fd_sc_hd__a22oi_2 _10123_ (.A1(_03446_),
    .A2(_03468_),
    .B1(_00567_),
    .B2(_00568_),
    .Y(_01792_));
 sky130_fd_sc_hd__o211ai_4 _10124_ (.A1(_03435_),
    .A2(_03457_),
    .B1(net147),
    .C1(net146),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_2 _10125_ (.A(_01602_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__o21ai_1 _10126_ (.A1(net9),
    .A2(_00893_),
    .B1(net156),
    .Y(_01796_));
 sky130_fd_sc_hd__o211ai_4 _10127_ (.A1(_03435_),
    .A2(_03457_),
    .B1(_00899_),
    .C1(_00902_),
    .Y(_01797_));
 sky130_fd_sc_hd__and3_1 _10128_ (.A(_01792_),
    .B(_00904_),
    .C(_02866_),
    .X(_01798_));
 sky130_fd_sc_hd__nand3_1 _10129_ (.A(_01792_),
    .B(_00904_),
    .C(_02866_),
    .Y(_01799_));
 sky130_fd_sc_hd__o21ai_1 _10130_ (.A1(_01604_),
    .A2(_01797_),
    .B1(_01794_),
    .Y(_01800_));
 sky130_fd_sc_hd__o211a_1 _10131_ (.A1(net170),
    .A2(_02057_),
    .B1(_01055_),
    .C1(_01057_),
    .X(_01801_));
 sky130_fd_sc_hd__a22oi_2 _10132_ (.A1(_02133_),
    .A2(net141),
    .B1(_01794_),
    .B2(_01799_),
    .Y(_01802_));
 sky130_fd_sc_hd__o21ai_4 _10133_ (.A1(_02122_),
    .A2(_01058_),
    .B1(_01800_),
    .Y(_01803_));
 sky130_fd_sc_hd__o311a_1 _10134_ (.A1(net158),
    .A2(_01604_),
    .A3(_00903_),
    .B1(_01801_),
    .C1(_01794_),
    .X(_01804_));
 sky130_fd_sc_hd__o211ai_4 _10135_ (.A1(_01604_),
    .A2(_01797_),
    .B1(_01794_),
    .C1(_01801_),
    .Y(_01805_));
 sky130_fd_sc_hd__o22ai_2 _10136_ (.A1(_01620_),
    .A2(_01221_),
    .B1(_01802_),
    .B2(_01804_),
    .Y(_01807_));
 sky130_fd_sc_hd__o2111ai_4 _10137_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_01222_),
    .C1(_01803_),
    .D1(_01805_),
    .Y(_01808_));
 sky130_fd_sc_hd__o21bai_2 _10138_ (.A1(_01802_),
    .A2(_01804_),
    .B1_N(_01791_),
    .Y(_01809_));
 sky130_fd_sc_hd__o211ai_2 _10139_ (.A1(_01620_),
    .A2(_01221_),
    .B1(_01803_),
    .C1(_01805_),
    .Y(_01810_));
 sky130_fd_sc_hd__nand2_1 _10140_ (.A(_01809_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__o211ai_2 _10141_ (.A1(_01787_),
    .A2(_01789_),
    .B1(_01809_),
    .C1(_01810_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand4_2 _10142_ (.A(_01788_),
    .B(_01790_),
    .C(_01807_),
    .D(_01808_),
    .Y(_01813_));
 sky130_fd_sc_hd__o211ai_1 _10143_ (.A1(_01787_),
    .A2(_01789_),
    .B1(_01807_),
    .C1(_01808_),
    .Y(_01814_));
 sky130_fd_sc_hd__nand4_1 _10144_ (.A(_01788_),
    .B(_01790_),
    .C(_01809_),
    .D(_01810_),
    .Y(_01815_));
 sky130_fd_sc_hd__nand3_2 _10145_ (.A(_01785_),
    .B(_01814_),
    .C(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand4_4 _10146_ (.A(_01613_),
    .B(_01783_),
    .C(_01812_),
    .D(_01813_),
    .Y(_01818_));
 sky130_fd_sc_hd__inv_2 _10147_ (.A(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__o211ai_4 _10148_ (.A1(net14),
    .A2(_01582_),
    .B1(net15),
    .C1(net174),
    .Y(_01820_));
 sky130_fd_sc_hd__o211ai_4 _10149_ (.A1(_00321_),
    .A2(_00693_),
    .B1(_00715_),
    .C1(_01583_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_8 _10150_ (.A(_01820_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__and2_4 _10151_ (.A(_01820_),
    .B(_01821_),
    .X(_01823_));
 sky130_fd_sc_hd__and3_1 _10152_ (.A(_01821_),
    .B(net33),
    .C(_01820_),
    .X(_01824_));
 sky130_fd_sc_hd__nand3_1 _10153_ (.A(_01821_),
    .B(net33),
    .C(_01820_),
    .Y(_01825_));
 sky130_fd_sc_hd__o211ai_2 _10154_ (.A1(_01238_),
    .A2(_01249_),
    .B1(_01585_),
    .C1(_01588_),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _10155_ (.A(_01596_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__o32a_1 _10156_ (.A1(_00900_),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01292_),
    .B2(_01406_),
    .X(_01829_));
 sky130_fd_sc_hd__a32o_1 _10157_ (.A1(_00911_),
    .A2(_01585_),
    .A3(_01588_),
    .B1(_01405_),
    .B2(_01303_),
    .X(_01830_));
 sky130_fd_sc_hd__o211a_1 _10158_ (.A1(_01827_),
    .A2(_01829_),
    .B1(net33),
    .C1(_01823_),
    .X(_01831_));
 sky130_fd_sc_hd__o311a_1 _10159_ (.A1(_01292_),
    .A2(_01589_),
    .A3(_01596_),
    .B1(_01825_),
    .C1(_01830_),
    .X(_01832_));
 sky130_fd_sc_hd__or2_1 _10160_ (.A(_01831_),
    .B(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__nor2_1 _10161_ (.A(_01831_),
    .B(_01832_),
    .Y(_01834_));
 sky130_fd_sc_hd__a21oi_1 _10162_ (.A1(_01816_),
    .A2(_01818_),
    .B1(_01833_),
    .Y(_01835_));
 sky130_fd_sc_hd__and3_1 _10163_ (.A(_01833_),
    .B(_01818_),
    .C(_01816_),
    .X(_01836_));
 sky130_fd_sc_hd__nand3_1 _10164_ (.A(_01816_),
    .B(_01818_),
    .C(_01834_),
    .Y(_01837_));
 sky130_fd_sc_hd__o2bb2ai_1 _10165_ (.A1_N(_01816_),
    .A2_N(_01818_),
    .B1(_01831_),
    .B2(_01832_),
    .Y(_01838_));
 sky130_fd_sc_hd__a21boi_2 _10166_ (.A1(_01619_),
    .A2(_01591_),
    .B1_N(_01618_),
    .Y(_01840_));
 sky130_fd_sc_hd__and3_1 _10167_ (.A(_01837_),
    .B(_01838_),
    .C(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__nand3_1 _10168_ (.A(_01837_),
    .B(_01838_),
    .C(_01840_),
    .Y(_01842_));
 sky130_fd_sc_hd__a21oi_1 _10169_ (.A1(_01837_),
    .A2(_01838_),
    .B1(_01840_),
    .Y(_01843_));
 sky130_fd_sc_hd__o21ai_1 _10170_ (.A1(_01430_),
    .A2(_01632_),
    .B1(_01628_),
    .Y(_01844_));
 sky130_fd_sc_hd__o21ai_1 _10171_ (.A1(_01580_),
    .A2(_01627_),
    .B1(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__o21a_1 _10172_ (.A1(_01841_),
    .A2(_01843_),
    .B1(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__nor3_1 _10173_ (.A(_01841_),
    .B(_01843_),
    .C(_01845_),
    .Y(_01847_));
 sky130_fd_sc_hd__or2_1 _10174_ (.A(_01846_),
    .B(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__a21oi_1 _10175_ (.A1(_01780_),
    .A2(_01781_),
    .B1(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__a21o_1 _10176_ (.A1(_01780_),
    .A2(_01781_),
    .B1(_01848_),
    .X(_01850_));
 sky130_fd_sc_hd__and3_1 _10177_ (.A(_01780_),
    .B(_01781_),
    .C(_01848_),
    .X(_01851_));
 sky130_fd_sc_hd__o211ai_1 _10178_ (.A1(_01846_),
    .A2(_01847_),
    .B1(_01780_),
    .C1(_01781_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _10179_ (.A(_01849_),
    .B(_01851_),
    .Y(_01853_));
 sky130_fd_sc_hd__a21o_1 _10180_ (.A1(_01850_),
    .A2(_01852_),
    .B1(_01646_),
    .X(_01854_));
 sky130_fd_sc_hd__nand3_1 _10181_ (.A(_01646_),
    .B(_01850_),
    .C(_01852_),
    .Y(_01855_));
 sky130_fd_sc_hd__o211ai_1 _10182_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_01638_),
    .C1(_01641_),
    .Y(_01856_));
 sky130_fd_sc_hd__a21bo_1 _10183_ (.A1(_01643_),
    .A2(_01639_),
    .B1_N(_01638_),
    .X(_01857_));
 sky130_fd_sc_hd__a21oi_1 _10184_ (.A1(_01854_),
    .A2(_01855_),
    .B1(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__and3_1 _10185_ (.A(_01857_),
    .B(_01855_),
    .C(_01854_),
    .X(_01859_));
 sky130_fd_sc_hd__or2_1 _10186_ (.A(_01858_),
    .B(_01859_),
    .X(_01861_));
 sky130_fd_sc_hd__or4_1 _10187_ (.A(_00834_),
    .B(_01645_),
    .C(_01858_),
    .D(_01859_),
    .X(_01862_));
 sky130_fd_sc_hd__o21ai_1 _10188_ (.A1(_00834_),
    .A2(_01645_),
    .B1(_01861_),
    .Y(_01863_));
 sky130_fd_sc_hd__and2_1 _10189_ (.A(_01862_),
    .B(_01863_),
    .X(net79));
 sky130_fd_sc_hd__a2bb2o_1 _10190_ (.A1_N(_00812_),
    .A2_N(_00823_),
    .B1(_01645_),
    .B2(_01861_),
    .X(_01864_));
 sky130_fd_sc_hd__o311ai_4 _10191_ (.A1(_01528_),
    .A2(_01570_),
    .A3(_01571_),
    .B1(_01704_),
    .C1(_01706_),
    .Y(_01865_));
 sky130_fd_sc_hd__o221ai_2 _10192_ (.A1(_01567_),
    .A2(_01572_),
    .B1(_01301_),
    .B2(_01573_),
    .C1(_01703_),
    .Y(_01866_));
 sky130_fd_sc_hd__o21a_1 _10193_ (.A1(_01692_),
    .A2(_01693_),
    .B1(_01687_),
    .X(_01867_));
 sky130_fd_sc_hd__nor2_1 _10194_ (.A(_01686_),
    .B(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__a31oi_2 _10195_ (.A1(_01650_),
    .A2(_01678_),
    .A3(_01679_),
    .B1(_01648_),
    .Y(_01869_));
 sky130_fd_sc_hd__and3_1 _10196_ (.A(_01969_),
    .B(_01269_),
    .C(_01271_),
    .X(_01871_));
 sky130_fd_sc_hd__or3_2 _10197_ (.A(_01958_),
    .B(_01184_),
    .C(_01186_),
    .X(_01872_));
 sky130_fd_sc_hd__o32a_1 _10198_ (.A1(_01958_),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_01272_),
    .B2(_01488_),
    .X(_01873_));
 sky130_fd_sc_hd__a21oi_2 _10199_ (.A1(_01651_),
    .A2(_01871_),
    .B1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__and3_1 _10200_ (.A(net164),
    .B(_01539_),
    .C(_01541_),
    .X(_01875_));
 sky130_fd_sc_hd__a221o_1 _10201_ (.A1(_01106_),
    .A2(_01128_),
    .B1(_01535_),
    .B2(_01537_),
    .C1(_01540_),
    .X(_01876_));
 sky130_fd_sc_hd__a41oi_4 _10202_ (.A1(_01179_),
    .A2(_01534_),
    .A3(_00682_),
    .A4(_00704_),
    .B1(_00299_),
    .Y(_01877_));
 sky130_fd_sc_hd__o311a_2 _10203_ (.A1(net46),
    .A2(net47),
    .A3(_01535_),
    .B1(net48),
    .C1(net173),
    .X(_01878_));
 sky130_fd_sc_hd__o211ai_4 _10204_ (.A1(net47),
    .A2(_01656_),
    .B1(net48),
    .C1(net173),
    .Y(_01879_));
 sky130_fd_sc_hd__o211ai_4 _10205_ (.A1(_00299_),
    .A2(_00704_),
    .B1(_00726_),
    .C1(_01657_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_8 _10206_ (.A(_01879_),
    .B(net134),
    .Y(_01882_));
 sky130_fd_sc_hd__and2_4 _10207_ (.A(_01879_),
    .B(net134),
    .X(_01883_));
 sky130_fd_sc_hd__nand3_1 _10208_ (.A(_01880_),
    .B(net1),
    .C(net135),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_2 _10209_ (.A(_01667_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__o211ai_4 _10210_ (.A1(_00921_),
    .A2(_00943_),
    .B1(net135),
    .C1(_01880_),
    .Y(_01886_));
 sky130_fd_sc_hd__o2111ai_4 _10211_ (.A1(_00921_),
    .A2(_00943_),
    .B1(net1),
    .C1(net135),
    .D1(_01880_),
    .Y(_01887_));
 sky130_fd_sc_hd__o2bb2ai_1 _10212_ (.A1_N(_01667_),
    .A2_N(_01884_),
    .B1(_01662_),
    .B2(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__o21ai_2 _10213_ (.A1(net166),
    .A2(_01542_),
    .B1(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__o211ai_4 _10214_ (.A1(_01665_),
    .A2(_01886_),
    .B1(_01875_),
    .C1(_01885_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _10215_ (.A(_01888_),
    .B(_01875_),
    .Y(_01891_));
 sky130_fd_sc_hd__o211ai_2 _10216_ (.A1(_01887_),
    .A2(_01662_),
    .B1(_01876_),
    .C1(_01885_),
    .Y(_01893_));
 sky130_fd_sc_hd__a21oi_1 _10217_ (.A1(_01889_),
    .A2(_01890_),
    .B1(_01874_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand3b_4 _10218_ (.A_N(_01874_),
    .B(_01891_),
    .C(_01893_),
    .Y(_01895_));
 sky130_fd_sc_hd__nand3_2 _10219_ (.A(_01889_),
    .B(_01890_),
    .C(_01874_),
    .Y(_01896_));
 sky130_fd_sc_hd__o211ai_1 _10220_ (.A1(_01545_),
    .A2(_01667_),
    .B1(_01895_),
    .C1(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__a21o_1 _10221_ (.A1(_01895_),
    .A2(_01896_),
    .B1(_01669_),
    .X(_01898_));
 sky130_fd_sc_hd__o2bb2ai_2 _10222_ (.A1_N(_01895_),
    .A2_N(_01896_),
    .B1(_01545_),
    .B2(_01667_),
    .Y(_01899_));
 sky130_fd_sc_hd__nand3_2 _10223_ (.A(_01895_),
    .B(_01896_),
    .C(_01668_),
    .Y(_01900_));
 sky130_fd_sc_hd__a2111oi_4 _10224_ (.A1(_03862_),
    .A2(_03873_),
    .B1(_00576_),
    .C1(_00578_),
    .D1(_01689_),
    .Y(_01901_));
 sky130_fd_sc_hd__a21oi_1 _10225_ (.A1(_03917_),
    .A2(_00581_),
    .B1(_01688_),
    .Y(_01902_));
 sky130_fd_sc_hd__a31o_1 _10226_ (.A1(_01666_),
    .A2(_01669_),
    .A3(_01670_),
    .B1(_01651_),
    .X(_01904_));
 sky130_fd_sc_hd__o221a_2 _10227_ (.A1(_01689_),
    .A2(_01902_),
    .B1(_01653_),
    .B2(_01671_),
    .C1(_01675_),
    .X(_01905_));
 sky130_fd_sc_hd__a211o_1 _10228_ (.A1(_01672_),
    .A2(_01904_),
    .B1(_01901_),
    .C1(_01688_),
    .X(_01906_));
 sky130_fd_sc_hd__o211a_2 _10229_ (.A1(_01688_),
    .A2(_01901_),
    .B1(_01904_),
    .C1(_01672_),
    .X(_01907_));
 sky130_fd_sc_hd__o211ai_4 _10230_ (.A1(_01688_),
    .A2(_01901_),
    .B1(_01904_),
    .C1(_01672_),
    .Y(_01908_));
 sky130_fd_sc_hd__nor2_1 _10231_ (.A(_01905_),
    .B(_01907_),
    .Y(_01909_));
 sky130_fd_sc_hd__nand4_1 _10232_ (.A(_01899_),
    .B(_01900_),
    .C(_01906_),
    .D(_01908_),
    .Y(_01910_));
 sky130_fd_sc_hd__o211ai_1 _10233_ (.A1(_01905_),
    .A2(_01907_),
    .B1(_01897_),
    .C1(_01898_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand3_1 _10234_ (.A(_01909_),
    .B(_01898_),
    .C(_01897_),
    .Y(_01912_));
 sky130_fd_sc_hd__o211ai_2 _10235_ (.A1(_01905_),
    .A2(_01907_),
    .B1(_01899_),
    .C1(_01900_),
    .Y(_01913_));
 sky130_fd_sc_hd__nand3_2 _10236_ (.A(_01911_),
    .B(_01869_),
    .C(_01910_),
    .Y(_01915_));
 sky130_fd_sc_hd__nand3b_4 _10237_ (.A_N(_01869_),
    .B(_01912_),
    .C(_01913_),
    .Y(_01916_));
 sky130_fd_sc_hd__o32a_4 _10238_ (.A1(_02636_),
    .A2(_01033_),
    .A3(_01035_),
    .B1(_03906_),
    .B2(_00744_),
    .X(_01917_));
 sky130_fd_sc_hd__and3_1 _10239_ (.A(_03917_),
    .B(_01034_),
    .C(_01036_),
    .X(_01918_));
 sky130_fd_sc_hd__and3_2 _10240_ (.A(_01918_),
    .B(_02647_),
    .C(_00743_),
    .X(_01919_));
 sky130_fd_sc_hd__o32a_1 _10241_ (.A1(_04244_),
    .A2(_00576_),
    .A3(_00578_),
    .B1(_01917_),
    .B2(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__a2111oi_2 _10242_ (.A1(_04201_),
    .A2(_04212_),
    .B1(_00580_),
    .C1(_01917_),
    .D1(_01919_),
    .Y(_01921_));
 sky130_fd_sc_hd__o211a_1 _10243_ (.A1(_01917_),
    .A2(_01919_),
    .B1(_04255_),
    .C1(_00581_),
    .X(_01922_));
 sky130_fd_sc_hd__a311oi_2 _10244_ (.A1(_04222_),
    .A2(_04233_),
    .A3(_00581_),
    .B1(_01917_),
    .C1(_01919_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_1 _10245_ (.A(_01920_),
    .B(_01921_),
    .Y(_01924_));
 sky130_fd_sc_hd__o211ai_2 _10246_ (.A1(_01920_),
    .A2(_01921_),
    .B1(_01915_),
    .C1(_01916_),
    .Y(_01926_));
 sky130_fd_sc_hd__o2bb2ai_1 _10247_ (.A1_N(_01915_),
    .A2_N(_01916_),
    .B1(_01922_),
    .B2(_01923_),
    .Y(_01927_));
 sky130_fd_sc_hd__o211ai_2 _10248_ (.A1(_01922_),
    .A2(_01923_),
    .B1(_01915_),
    .C1(_01916_),
    .Y(_01928_));
 sky130_fd_sc_hd__o2bb2ai_1 _10249_ (.A1_N(_01915_),
    .A2_N(_01916_),
    .B1(_01920_),
    .B2(_01921_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand3_4 _10250_ (.A(_01868_),
    .B(_01926_),
    .C(_01927_),
    .Y(_01930_));
 sky130_fd_sc_hd__o211ai_4 _10251_ (.A1(_01686_),
    .A2(_01867_),
    .B1(_01928_),
    .C1(_01929_),
    .Y(_01931_));
 sky130_fd_sc_hd__a22oi_2 _10252_ (.A1(_01703_),
    .A2(_01865_),
    .B1(_01930_),
    .B2(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__o211ai_2 _10253_ (.A1(_01702_),
    .A2(_01698_),
    .B1(_01930_),
    .C1(_01866_),
    .Y(_01933_));
 sky130_fd_sc_hd__o211ai_4 _10254_ (.A1(_01701_),
    .A2(_01697_),
    .B1(_01931_),
    .C1(_01865_),
    .Y(_01934_));
 sky130_fd_sc_hd__a41oi_4 _10255_ (.A1(_01703_),
    .A2(_01865_),
    .A3(_01930_),
    .A4(_01931_),
    .B1(_01932_),
    .Y(_01935_));
 sky130_fd_sc_hd__o21bai_4 _10256_ (.A1(_01715_),
    .A2(_01763_),
    .B1_N(_01761_),
    .Y(_01937_));
 sky130_fd_sc_hd__inv_2 _10257_ (.A(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__a31o_1 _10258_ (.A1(_05436_),
    .A2(_00367_),
    .A3(_01741_),
    .B1(_01738_),
    .X(_01939_));
 sky130_fd_sc_hd__a31o_1 _10259_ (.A1(_07509_),
    .A2(_07511_),
    .A3(_07540_),
    .B1(_01727_),
    .X(_01940_));
 sky130_fd_sc_hd__and3_1 _10260_ (.A(_01731_),
    .B(_01939_),
    .C(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__a311o_1 _10261_ (.A1(_07513_),
    .A2(_07540_),
    .A3(_01731_),
    .B1(_01939_),
    .C1(_01727_),
    .X(_01942_));
 sky130_fd_sc_hd__nand2b_1 _10262_ (.A_N(_01941_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__or4_2 _10263_ (.A(_07512_),
    .B(_07539_),
    .C(_00009_),
    .D(_00071_),
    .X(_01944_));
 sky130_fd_sc_hd__a32o_1 _10264_ (.A1(_07540_),
    .A2(_00006_),
    .A3(_00008_),
    .B1(_00072_),
    .B2(_07513_),
    .X(_01945_));
 sky130_fd_sc_hd__and4_1 _10265_ (.A(_07200_),
    .B(_00275_),
    .C(_00429_),
    .D(_05316_),
    .X(_01946_));
 sky130_fd_sc_hd__nand4_1 _10266_ (.A(_07200_),
    .B(_00275_),
    .C(_00429_),
    .D(_05316_),
    .Y(_01948_));
 sky130_fd_sc_hd__a32o_1 _10267_ (.A1(_05316_),
    .A2(_00425_),
    .A3(_00427_),
    .B1(_07200_),
    .B2(_00275_),
    .X(_01949_));
 sky130_fd_sc_hd__a32o_1 _10268_ (.A1(_07436_),
    .A2(net154),
    .A3(_00150_),
    .B1(_01948_),
    .B2(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__nand4_1 _10269_ (.A(_00150_),
    .B(_01948_),
    .C(_01949_),
    .D(_07440_),
    .Y(_01951_));
 sky130_fd_sc_hd__a22o_1 _10270_ (.A1(_01944_),
    .A2(_01945_),
    .B1(_01950_),
    .B2(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__nand4_2 _10271_ (.A(_01944_),
    .B(_01945_),
    .C(_01950_),
    .D(_01951_),
    .Y(_01953_));
 sky130_fd_sc_hd__a21oi_1 _10272_ (.A1(_01952_),
    .A2(_01953_),
    .B1(_01725_),
    .Y(_01954_));
 sky130_fd_sc_hd__and3_1 _10273_ (.A(_01952_),
    .B(_01953_),
    .C(_01725_),
    .X(_01955_));
 sky130_fd_sc_hd__nor2_1 _10274_ (.A(_01954_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__nand2_1 _10275_ (.A(_01943_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__o21bai_2 _10276_ (.A1(_01954_),
    .A2(_01955_),
    .B1_N(_01943_),
    .Y(_01959_));
 sky130_fd_sc_hd__a21bo_1 _10277_ (.A1(_01721_),
    .A2(_01734_),
    .B1_N(_01720_),
    .X(_01960_));
 sky130_fd_sc_hd__nand3_1 _10278_ (.A(_01957_),
    .B(_01959_),
    .C(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__a21oi_1 _10279_ (.A1(_01957_),
    .A2(_01959_),
    .B1(_01960_),
    .Y(_01962_));
 sky130_fd_sc_hd__a21o_1 _10280_ (.A1(_01957_),
    .A2(_01959_),
    .B1(_01960_),
    .X(_01963_));
 sky130_fd_sc_hd__nand2_1 _10281_ (.A(_01961_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__o32a_1 _10282_ (.A1(_06331_),
    .A2(_00361_),
    .A3(_00363_),
    .B1(net153),
    .B2(_00192_),
    .X(_01965_));
 sky130_fd_sc_hd__a32o_1 _10283_ (.A1(_06341_),
    .A2(_00362_),
    .A3(_00364_),
    .B1(net151),
    .B2(_00193_),
    .X(_01966_));
 sky130_fd_sc_hd__or4_1 _10284_ (.A(_06331_),
    .B(net153),
    .C(_00192_),
    .D(_00366_),
    .X(_01967_));
 sky130_fd_sc_hd__a211o_1 _10285_ (.A1(_01966_),
    .A2(_01967_),
    .B1(_05425_),
    .C1(_00532_),
    .X(_01968_));
 sky130_fd_sc_hd__o211ai_1 _10286_ (.A1(_05425_),
    .A2(_00532_),
    .B1(_01966_),
    .C1(_01967_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _10287_ (.A(_01968_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__xnor2_1 _10288_ (.A(_01964_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__a21o_1 _10289_ (.A1(_01735_),
    .A2(_01736_),
    .B1(_01744_),
    .X(_01973_));
 sky130_fd_sc_hd__o21ai_1 _10290_ (.A1(_01735_),
    .A2(_01736_),
    .B1(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(_01972_),
    .B(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__or2_1 _10292_ (.A(_01974_),
    .B(_01972_),
    .X(_01976_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(_01975_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__o21ai_1 _10294_ (.A1(_01747_),
    .A2(_01749_),
    .B1(_01746_),
    .Y(_01978_));
 sky130_fd_sc_hd__xnor2_1 _10295_ (.A(_01977_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand3_1 _10296_ (.A(_01467_),
    .B(_01755_),
    .C(_01758_),
    .Y(_01981_));
 sky130_fd_sc_hd__nand3_1 _10297_ (.A(_01979_),
    .B(_01981_),
    .C(_01754_),
    .Y(_01982_));
 sky130_fd_sc_hd__a21oi_1 _10298_ (.A1(_01754_),
    .A2(_01981_),
    .B1(_01979_),
    .Y(_01983_));
 sky130_fd_sc_hd__a21o_1 _10299_ (.A1(_01754_),
    .A2(_01981_),
    .B1(_01979_),
    .X(_01984_));
 sky130_fd_sc_hd__a21oi_2 _10300_ (.A1(_01714_),
    .A2(_01712_),
    .B1(_01711_),
    .Y(_01985_));
 sky130_fd_sc_hd__and3_2 _10301_ (.A(_01982_),
    .B(_01984_),
    .C(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__a21oi_1 _10302_ (.A1(_01982_),
    .A2(_01984_),
    .B1(_01985_),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2_1 _10303_ (.A(_01986_),
    .B(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__or2_1 _10304_ (.A(_01986_),
    .B(_01987_),
    .X(_01989_));
 sky130_fd_sc_hd__o21ai_2 _10305_ (.A1(_01986_),
    .A2(_01987_),
    .B1(_01938_),
    .Y(_01990_));
 sky130_fd_sc_hd__or2_2 _10306_ (.A(_01938_),
    .B(_01987_),
    .X(_01992_));
 sky130_fd_sc_hd__a31o_1 _10307_ (.A1(_01982_),
    .A2(_01984_),
    .A3(_01985_),
    .B1(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__o21ai_1 _10308_ (.A1(_01986_),
    .A2(_01992_),
    .B1(_01990_),
    .Y(_01994_));
 sky130_fd_sc_hd__o221ai_4 _10309_ (.A1(_01376_),
    .A2(_01516_),
    .B1(_01766_),
    .B2(_01768_),
    .C1(_01774_),
    .Y(_01995_));
 sky130_fd_sc_hd__o211ai_2 _10310_ (.A1(_01377_),
    .A2(_01517_),
    .B1(_01770_),
    .C1(_01775_),
    .Y(_01996_));
 sky130_fd_sc_hd__nand3_1 _10311_ (.A(_01770_),
    .B(_01994_),
    .C(_01995_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand4_1 _10312_ (.A(_01769_),
    .B(_01990_),
    .C(_01993_),
    .D(_01996_),
    .Y(_01998_));
 sky130_fd_sc_hd__o2111ai_1 _10313_ (.A1(_01992_),
    .A2(_01986_),
    .B1(_01770_),
    .C1(_01990_),
    .D1(_01995_),
    .Y(_01999_));
 sky130_fd_sc_hd__o211ai_1 _10314_ (.A1(_01766_),
    .A2(_01768_),
    .B1(_01994_),
    .C1(_01996_),
    .Y(_02000_));
 sky130_fd_sc_hd__nand3b_2 _10315_ (.A_N(_01935_),
    .B(_01999_),
    .C(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__nand3_1 _10316_ (.A(_01998_),
    .B(_01935_),
    .C(_01997_),
    .Y(_02003_));
 sky130_fd_sc_hd__o21a_1 _10317_ (.A1(_01831_),
    .A2(_01832_),
    .B1(_01816_),
    .X(_02004_));
 sky130_fd_sc_hd__and3_1 _10318_ (.A(_01788_),
    .B(_01807_),
    .C(_01808_),
    .X(_02005_));
 sky130_fd_sc_hd__o21ai_1 _10319_ (.A1(_01789_),
    .A2(_01811_),
    .B1(_01788_),
    .Y(_02006_));
 sky130_fd_sc_hd__o21ai_1 _10320_ (.A1(_01596_),
    .A2(_01826_),
    .B1(_01825_),
    .Y(_02007_));
 sky130_fd_sc_hd__o21ai_2 _10321_ (.A1(_01620_),
    .A2(_01221_),
    .B1(_01805_),
    .Y(_02008_));
 sky130_fd_sc_hd__o2111a_1 _10322_ (.A1(_01824_),
    .A2(_01827_),
    .B1(_01830_),
    .C1(_02008_),
    .D1(_01803_),
    .X(_02009_));
 sky130_fd_sc_hd__o2111ai_2 _10323_ (.A1(_01824_),
    .A2(_01827_),
    .B1(_01830_),
    .C1(_02008_),
    .D1(_01803_),
    .Y(_02010_));
 sky130_fd_sc_hd__a22oi_2 _10324_ (.A1(_01830_),
    .A2(_02007_),
    .B1(_02008_),
    .B2(_01803_),
    .Y(_02011_));
 sky130_fd_sc_hd__a22o_1 _10325_ (.A1(_01830_),
    .A2(_02007_),
    .B1(_02008_),
    .B2(_01803_),
    .X(_02012_));
 sky130_fd_sc_hd__a21oi_1 _10326_ (.A1(_01397_),
    .A2(_01402_),
    .B1(_01620_),
    .Y(_02014_));
 sky130_fd_sc_hd__o21ai_2 _10327_ (.A1(net13),
    .A2(_01398_),
    .B1(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__o31ai_2 _10328_ (.A1(_02122_),
    .A2(_01217_),
    .A3(_01219_),
    .B1(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__o221ai_4 _10329_ (.A1(net170),
    .A2(_02057_),
    .B1(_01396_),
    .B2(_01403_),
    .C1(_01400_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand4_1 _10330_ (.A(_01222_),
    .B(_02014_),
    .C(_01400_),
    .D(_02133_),
    .Y(_02018_));
 sky130_fd_sc_hd__o21ai_1 _10331_ (.A1(_01791_),
    .A2(_02017_),
    .B1(_02016_),
    .Y(_02019_));
 sky130_fd_sc_hd__o211ai_2 _10332_ (.A1(_04638_),
    .A2(_04649_),
    .B1(net147),
    .C1(net146),
    .Y(_02020_));
 sky130_fd_sc_hd__o21ai_4 _10333_ (.A1(_00898_),
    .A2(_01796_),
    .B1(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__o211ai_4 _10334_ (.A1(_04638_),
    .A2(_04649_),
    .B1(_00899_),
    .C1(_00902_),
    .Y(_02022_));
 sky130_fd_sc_hd__and3_1 _10335_ (.A(_01792_),
    .B(_00904_),
    .C(_04726_),
    .X(_02023_));
 sky130_fd_sc_hd__o2bb2ai_1 _10336_ (.A1_N(_01797_),
    .A2_N(_02020_),
    .B1(_02022_),
    .B2(_01793_),
    .Y(_02025_));
 sky130_fd_sc_hd__o21ai_1 _10337_ (.A1(net159),
    .A2(_01058_),
    .B1(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__o2111ai_1 _10338_ (.A1(_01793_),
    .A2(_02022_),
    .B1(_02021_),
    .C1(_02866_),
    .D1(net141),
    .Y(_02027_));
 sky130_fd_sc_hd__o211ai_2 _10339_ (.A1(net168),
    .A2(net163),
    .B1(net141),
    .C1(_02025_),
    .Y(_02028_));
 sky130_fd_sc_hd__o221ai_4 _10340_ (.A1(_01793_),
    .A2(_02022_),
    .B1(net159),
    .B2(_01058_),
    .C1(_02021_),
    .Y(_02029_));
 sky130_fd_sc_hd__a22oi_2 _10341_ (.A1(_02016_),
    .A2(_02018_),
    .B1(_02026_),
    .B2(_02027_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand3_2 _10342_ (.A(_02019_),
    .B(_02028_),
    .C(_02029_),
    .Y(_02031_));
 sky130_fd_sc_hd__a21oi_1 _10343_ (.A1(_02028_),
    .A2(_02029_),
    .B1(_02019_),
    .Y(_02032_));
 sky130_fd_sc_hd__a21o_2 _10344_ (.A1(_02028_),
    .A2(_02029_),
    .B1(_02019_),
    .X(_02033_));
 sky130_fd_sc_hd__o211ai_2 _10345_ (.A1(_01602_),
    .A2(_01793_),
    .B1(_02031_),
    .C1(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__o21ai_2 _10346_ (.A1(_02030_),
    .A2(_02032_),
    .B1(_01798_),
    .Y(_02036_));
 sky130_fd_sc_hd__o21ai_1 _10347_ (.A1(_02030_),
    .A2(_02032_),
    .B1(_01799_),
    .Y(_02037_));
 sky130_fd_sc_hd__nand3_1 _10348_ (.A(_02033_),
    .B(_01798_),
    .C(_02031_),
    .Y(_02038_));
 sky130_fd_sc_hd__o211ai_1 _10349_ (.A1(_02009_),
    .A2(_02011_),
    .B1(_02037_),
    .C1(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand4_1 _10350_ (.A(_02010_),
    .B(_02012_),
    .C(_02034_),
    .D(_02036_),
    .Y(_02040_));
 sky130_fd_sc_hd__o211ai_2 _10351_ (.A1(_02009_),
    .A2(_02011_),
    .B1(_02034_),
    .C1(_02036_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand4_1 _10352_ (.A(_02010_),
    .B(_02012_),
    .C(_02037_),
    .D(_02038_),
    .Y(_02042_));
 sky130_fd_sc_hd__o211ai_4 _10353_ (.A1(_01789_),
    .A2(_02005_),
    .B1(_02041_),
    .C1(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__nand3_2 _10354_ (.A(_02040_),
    .B(_02006_),
    .C(_02039_),
    .Y(_02044_));
 sky130_fd_sc_hd__nor2_4 _10355_ (.A(net14),
    .B(net15),
    .Y(_02045_));
 sky130_fd_sc_hd__or2_2 _10356_ (.A(net14),
    .B(net15),
    .X(_02047_));
 sky130_fd_sc_hd__nand4b_4 _10357_ (.A_N(_01053_),
    .B(_01394_),
    .C(_02045_),
    .D(_00671_),
    .Y(_02048_));
 sky130_fd_sc_hd__a21oi_4 _10358_ (.A1(_02048_),
    .A2(net174),
    .B1(net16),
    .Y(_02049_));
 sky130_fd_sc_hd__a21o_4 _10359_ (.A1(_02048_),
    .A2(net174),
    .B1(net16),
    .X(_02050_));
 sky130_fd_sc_hd__o311a_4 _10360_ (.A1(_02047_),
    .A2(net13),
    .A3(_01397_),
    .B1(net16),
    .C1(net174),
    .X(_02051_));
 sky130_fd_sc_hd__o211ai_4 _10361_ (.A1(_01582_),
    .A2(_02047_),
    .B1(net174),
    .C1(net16),
    .Y(_02052_));
 sky130_fd_sc_hd__nand2_8 _10362_ (.A(_02050_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__nor2_8 _10363_ (.A(_02049_),
    .B(_02051_),
    .Y(_02054_));
 sky130_fd_sc_hd__o21ai_2 _10364_ (.A1(_00900_),
    .A2(_01822_),
    .B1(_01826_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand4_4 _10365_ (.A(_00911_),
    .B(_01303_),
    .C(_01590_),
    .D(_01823_),
    .Y(_02056_));
 sky130_fd_sc_hd__o2bb2a_1 _10366_ (.A1_N(_02055_),
    .A2_N(_02056_),
    .B1(_00310_),
    .B2(_02053_),
    .X(_02058_));
 sky130_fd_sc_hd__and4_1 _10367_ (.A(_02054_),
    .B(_02055_),
    .C(_02056_),
    .D(net33),
    .X(_02059_));
 sky130_fd_sc_hd__nor2_1 _10368_ (.A(_02058_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__or2_1 _10369_ (.A(_02058_),
    .B(_02059_),
    .X(_02061_));
 sky130_fd_sc_hd__a21oi_2 _10370_ (.A1(_02043_),
    .A2(_02044_),
    .B1(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__o211a_1 _10371_ (.A1(_02058_),
    .A2(_02059_),
    .B1(_02043_),
    .C1(_02044_),
    .X(_02063_));
 sky130_fd_sc_hd__a311o_1 _10372_ (.A1(_02043_),
    .A2(_02044_),
    .A3(_02061_),
    .B1(_02004_),
    .C1(_01819_),
    .X(_02064_));
 sky130_fd_sc_hd__nor2_1 _10373_ (.A(_02062_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__o22a_1 _10374_ (.A1(_01819_),
    .A2(_02004_),
    .B1(_02062_),
    .B2(_02063_),
    .X(_02066_));
 sky130_fd_sc_hd__o22ai_1 _10375_ (.A1(_01819_),
    .A2(_02004_),
    .B1(_02062_),
    .B2(_02063_),
    .Y(_02067_));
 sky130_fd_sc_hd__o211ai_2 _10376_ (.A1(_01580_),
    .A2(_01627_),
    .B1(_01842_),
    .C1(_01844_),
    .Y(_02069_));
 sky130_fd_sc_hd__o31a_1 _10377_ (.A1(_01835_),
    .A2(_01836_),
    .A3(_01840_),
    .B1(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__o21a_1 _10378_ (.A1(_02065_),
    .A2(_02066_),
    .B1(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__nor3_1 _10379_ (.A(_02070_),
    .B(_02066_),
    .C(_02065_),
    .Y(_02072_));
 sky130_fd_sc_hd__nor2_1 _10380_ (.A(_02071_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__o2bb2ai_1 _10381_ (.A1_N(_02001_),
    .A2_N(_02003_),
    .B1(_02071_),
    .B2(_02072_),
    .Y(_02074_));
 sky130_fd_sc_hd__a311o_1 _10382_ (.A1(_01997_),
    .A2(_01998_),
    .A3(_01935_),
    .B1(_02071_),
    .C1(_02072_),
    .X(_02075_));
 sky130_fd_sc_hd__nand3_1 _10383_ (.A(_02001_),
    .B(_02003_),
    .C(_02073_),
    .Y(_02076_));
 sky130_fd_sc_hd__and2b_1 _10384_ (.A_N(_01848_),
    .B(_01780_),
    .X(_02077_));
 sky130_fd_sc_hd__a211o_1 _10385_ (.A1(_02074_),
    .A2(_02076_),
    .B1(_02077_),
    .C1(_01782_),
    .X(_02078_));
 sky130_fd_sc_hd__o211ai_2 _10386_ (.A1(_01782_),
    .A2(_02077_),
    .B1(_02076_),
    .C1(_02074_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand3_1 _10387_ (.A(_01639_),
    .B(_01855_),
    .C(_01856_),
    .Y(_02081_));
 sky130_fd_sc_hd__and4_1 _10388_ (.A(_01854_),
    .B(_02078_),
    .C(_02080_),
    .D(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__a22oi_1 _10389_ (.A1(_02078_),
    .A2(_02080_),
    .B1(_02081_),
    .B2(_01854_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_1 _10390_ (.A(_02082_),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__xor2_1 _10391_ (.A(_01864_),
    .B(_02084_),
    .X(net80));
 sky130_fd_sc_hd__and3_1 _10392_ (.A(_01645_),
    .B(_01861_),
    .C(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__or3_4 _10393_ (.A(_05327_),
    .B(_00576_),
    .C(_00578_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_4 _10394_ (.A(net47),
    .B(net48),
    .Y(_02087_));
 sky130_fd_sc_hd__or2_2 _10395_ (.A(net47),
    .B(net48),
    .X(_02088_));
 sky130_fd_sc_hd__nor4_4 _10396_ (.A(net45),
    .B(_02088_),
    .C(net46),
    .D(_01265_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand4_4 _10397_ (.A(_01179_),
    .B(_01534_),
    .C(_02087_),
    .D(_00682_),
    .Y(_02091_));
 sky130_fd_sc_hd__a21oi_4 _10398_ (.A1(_02091_),
    .A2(net173),
    .B1(net49),
    .Y(_02092_));
 sky130_fd_sc_hd__a21o_2 _10399_ (.A1(_02091_),
    .A2(net173),
    .B1(net49),
    .X(_02093_));
 sky130_fd_sc_hd__o311a_4 _10400_ (.A1(_02088_),
    .A2(net46),
    .A3(_01535_),
    .B1(net49),
    .C1(net173),
    .X(_02094_));
 sky130_fd_sc_hd__or3b_4 _10401_ (.A(_00299_),
    .B(_02090_),
    .C_N(net49),
    .X(_02095_));
 sky130_fd_sc_hd__or2_4 _10402_ (.A(_02092_),
    .B(_02094_),
    .X(_02096_));
 sky130_fd_sc_hd__nor2_8 _10403_ (.A(_02092_),
    .B(_02094_),
    .Y(_02097_));
 sky130_fd_sc_hd__or3_4 _10404_ (.A(_00288_),
    .B(_02092_),
    .C(_02094_),
    .X(_02098_));
 sky130_fd_sc_hd__and3_1 _10405_ (.A(_01651_),
    .B(_01871_),
    .C(_01918_),
    .X(_02099_));
 sky130_fd_sc_hd__or4b_1 _10406_ (.A(_03906_),
    .B(_01037_),
    .C(_01653_),
    .D_N(_01871_),
    .X(_02101_));
 sky130_fd_sc_hd__a31o_1 _10407_ (.A1(_01651_),
    .A2(_01273_),
    .A3(_01969_),
    .B1(_01918_),
    .X(_02102_));
 sky130_fd_sc_hd__o2bb2a_1 _10408_ (.A1_N(_02101_),
    .A2_N(_02102_),
    .B1(_04244_),
    .B2(_00744_),
    .X(_02103_));
 sky130_fd_sc_hd__and4_1 _10409_ (.A(_04255_),
    .B(_02101_),
    .C(_02102_),
    .D(_00743_),
    .X(_02104_));
 sky130_fd_sc_hd__nor2_2 _10410_ (.A(_02103_),
    .B(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__and3_1 _10411_ (.A(_01899_),
    .B(_01900_),
    .C(_01906_),
    .X(_02106_));
 sky130_fd_sc_hd__nand3_1 _10412_ (.A(_01899_),
    .B(_01900_),
    .C(_01906_),
    .Y(_02107_));
 sky130_fd_sc_hd__a21oi_2 _10413_ (.A1(_01899_),
    .A2(_01900_),
    .B1(_01907_),
    .Y(_02108_));
 sky130_fd_sc_hd__a2111oi_4 _10414_ (.A1(_04201_),
    .A2(_04212_),
    .B1(_00576_),
    .C1(_00578_),
    .D1(_01917_),
    .Y(_02109_));
 sky130_fd_sc_hd__nor2_1 _10415_ (.A(_01919_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__a31oi_2 _10416_ (.A1(_01889_),
    .A2(_01890_),
    .A3(_01874_),
    .B1(_01668_),
    .Y(_02112_));
 sky130_fd_sc_hd__a31o_1 _10417_ (.A1(_01889_),
    .A2(_01890_),
    .A3(_01874_),
    .B1(_01668_),
    .X(_02113_));
 sky130_fd_sc_hd__o211a_1 _10418_ (.A1(_01919_),
    .A2(_02109_),
    .B1(_02113_),
    .C1(_01895_),
    .X(_02114_));
 sky130_fd_sc_hd__o211ai_4 _10419_ (.A1(_01919_),
    .A2(_02109_),
    .B1(_02113_),
    .C1(_01895_),
    .Y(_02115_));
 sky130_fd_sc_hd__o21ai_4 _10420_ (.A1(_01894_),
    .A2(_02112_),
    .B1(_02110_),
    .Y(_02116_));
 sky130_fd_sc_hd__a22o_2 _10421_ (.A1(_02592_),
    .A2(_02603_),
    .B1(_01266_),
    .B2(_01267_),
    .X(_02117_));
 sky130_fd_sc_hd__and3_1 _10422_ (.A(_02647_),
    .B(_01185_),
    .C(_01187_),
    .X(_02118_));
 sky130_fd_sc_hd__nor4_2 _10423_ (.A(_01958_),
    .B(_02636_),
    .C(_01188_),
    .D(_01272_),
    .Y(_02119_));
 sky130_fd_sc_hd__or4_2 _10424_ (.A(_01958_),
    .B(_02636_),
    .C(_01188_),
    .D(_01272_),
    .X(_02120_));
 sky130_fd_sc_hd__o32a_1 _10425_ (.A1(_02636_),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_01272_),
    .B2(_01958_),
    .X(_02121_));
 sky130_fd_sc_hd__nor2_1 _10426_ (.A(_02119_),
    .B(_02121_),
    .Y(_02123_));
 sky130_fd_sc_hd__and3_1 _10427_ (.A(net164),
    .B(_01659_),
    .C(net140),
    .X(_02124_));
 sky130_fd_sc_hd__o2111ai_2 _10428_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01172_),
    .C1(_01659_),
    .D1(net140),
    .Y(_02125_));
 sky130_fd_sc_hd__o21ai_4 _10429_ (.A1(net166),
    .A2(_01662_),
    .B1(_01886_),
    .Y(_02126_));
 sky130_fd_sc_hd__o211ai_4 _10430_ (.A1(_01095_),
    .A2(_01117_),
    .B1(net135),
    .C1(_01880_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _10431_ (.A(_01667_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__o2bb2ai_1 _10432_ (.A1_N(_01886_),
    .A2_N(_02125_),
    .B1(_02127_),
    .B2(_01667_),
    .Y(_02129_));
 sky130_fd_sc_hd__and3_1 _10433_ (.A(_01499_),
    .B(_01539_),
    .C(_01541_),
    .X(_02130_));
 sky130_fd_sc_hd__a221o_1 _10434_ (.A1(_01434_),
    .A2(_01455_),
    .B1(_01535_),
    .B2(_01537_),
    .C1(_01540_),
    .X(_02131_));
 sky130_fd_sc_hd__o21ai_2 _10435_ (.A1(_01488_),
    .A2(_01542_),
    .B1(_02129_),
    .Y(_02132_));
 sky130_fd_sc_hd__o211ai_2 _10436_ (.A1(_01667_),
    .A2(_02127_),
    .B1(_02130_),
    .C1(_02126_),
    .Y(_02134_));
 sky130_fd_sc_hd__o221ai_4 _10437_ (.A1(_01488_),
    .A2(_01542_),
    .B1(_01667_),
    .B2(_02127_),
    .C1(_02126_),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _10438_ (.A(_02129_),
    .B(_02130_),
    .Y(_02136_));
 sky130_fd_sc_hd__o211a_1 _10439_ (.A1(_02119_),
    .A2(_02121_),
    .B1(_02135_),
    .C1(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__o211ai_4 _10440_ (.A1(_02119_),
    .A2(_02121_),
    .B1(_02135_),
    .C1(_02136_),
    .Y(_02138_));
 sky130_fd_sc_hd__nand3_2 _10441_ (.A(_02132_),
    .B(_02134_),
    .C(_02123_),
    .Y(_02139_));
 sky130_fd_sc_hd__o2bb2a_1 _10442_ (.A1_N(_01875_),
    .A2_N(_01885_),
    .B1(_01887_),
    .B2(_01662_),
    .X(_02140_));
 sky130_fd_sc_hd__a2bb2o_2 _10443_ (.A1_N(_01662_),
    .A2_N(_01887_),
    .B1(_01875_),
    .B2(_01885_),
    .X(_02141_));
 sky130_fd_sc_hd__a21oi_1 _10444_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__a21o_1 _10445_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02141_),
    .X(_02143_));
 sky130_fd_sc_hd__and3_1 _10446_ (.A(_02138_),
    .B(_02139_),
    .C(_02141_),
    .X(_02145_));
 sky130_fd_sc_hd__nand3_2 _10447_ (.A(_02138_),
    .B(_02139_),
    .C(_02141_),
    .Y(_02146_));
 sky130_fd_sc_hd__a31oi_2 _10448_ (.A1(_02132_),
    .A2(_02134_),
    .A3(_02123_),
    .B1(_02141_),
    .Y(_02147_));
 sky130_fd_sc_hd__a31o_2 _10449_ (.A1(_02132_),
    .A2(_02134_),
    .A3(_02123_),
    .B1(_02141_),
    .X(_02148_));
 sky130_fd_sc_hd__and3_1 _10450_ (.A(_02138_),
    .B(_02139_),
    .C(_02140_),
    .X(_02149_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_02147_),
    .B(_02138_),
    .Y(_02150_));
 sky130_fd_sc_hd__a21oi_1 _10452_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02140_),
    .Y(_02151_));
 sky130_fd_sc_hd__a21o_1 _10453_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02140_),
    .X(_02152_));
 sky130_fd_sc_hd__o2bb2ai_4 _10454_ (.A1_N(_02115_),
    .A2_N(_02116_),
    .B1(_02149_),
    .B2(_02151_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand4_4 _10455_ (.A(_02115_),
    .B(_02116_),
    .C(_02150_),
    .D(_02152_),
    .Y(_02154_));
 sky130_fd_sc_hd__nand4_1 _10456_ (.A(_02115_),
    .B(_02116_),
    .C(_02143_),
    .D(_02146_),
    .Y(_02156_));
 sky130_fd_sc_hd__o2bb2ai_1 _10457_ (.A1_N(_02115_),
    .A2_N(_02116_),
    .B1(_02142_),
    .B2(_02145_),
    .Y(_02157_));
 sky130_fd_sc_hd__a22oi_4 _10458_ (.A1(_01908_),
    .A2(_02107_),
    .B1(_02153_),
    .B2(_02154_),
    .Y(_02158_));
 sky130_fd_sc_hd__o211ai_2 _10459_ (.A1(_01907_),
    .A2(_02106_),
    .B1(_02156_),
    .C1(_02157_),
    .Y(_02159_));
 sky130_fd_sc_hd__a2bb2oi_1 _10460_ (.A1_N(_01905_),
    .A2_N(_02108_),
    .B1(_02156_),
    .B2(_02157_),
    .Y(_02160_));
 sky130_fd_sc_hd__o211ai_4 _10461_ (.A1(_01905_),
    .A2(_02108_),
    .B1(_02153_),
    .C1(_02154_),
    .Y(_02161_));
 sky130_fd_sc_hd__o31a_2 _10462_ (.A1(_02103_),
    .A2(_02104_),
    .A3(_02160_),
    .B1(_02159_),
    .X(_02162_));
 sky130_fd_sc_hd__o211ai_2 _10463_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_02159_),
    .C1(_02161_),
    .Y(_02163_));
 sky130_fd_sc_hd__o21ai_2 _10464_ (.A1(_02158_),
    .A2(_02160_),
    .B1(_02105_),
    .Y(_02164_));
 sky130_fd_sc_hd__o22ai_1 _10465_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_02158_),
    .B2(_02160_),
    .Y(_02165_));
 sky130_fd_sc_hd__nand3_1 _10466_ (.A(_02159_),
    .B(_02161_),
    .C(_02105_),
    .Y(_02167_));
 sky130_fd_sc_hd__nand2_2 _10467_ (.A(_02165_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__a21boi_4 _10468_ (.A1(_01916_),
    .A2(_01924_),
    .B1_N(_01915_),
    .Y(_02169_));
 sky130_fd_sc_hd__nand3_4 _10469_ (.A(_02163_),
    .B(_02164_),
    .C(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__a21o_1 _10470_ (.A1(_02163_),
    .A2(_02164_),
    .B1(_02169_),
    .X(_02171_));
 sky130_fd_sc_hd__a22oi_4 _10471_ (.A1(_01930_),
    .A2(_01934_),
    .B1(_02170_),
    .B2(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__and4_1 _10472_ (.A(_01930_),
    .B(_01934_),
    .C(_02170_),
    .D(_02171_),
    .X(_02173_));
 sky130_fd_sc_hd__nor2_1 _10473_ (.A(_02172_),
    .B(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__o32a_1 _10474_ (.A1(_00288_),
    .A2(_02092_),
    .A3(_02094_),
    .B1(_02172_),
    .B2(_02173_),
    .X(_02175_));
 sky130_fd_sc_hd__xor2_2 _10475_ (.A(_02098_),
    .B(_02174_),
    .X(_02176_));
 sky130_fd_sc_hd__xnor2_4 _10476_ (.A(_02086_),
    .B(_02176_),
    .Y(_02178_));
 sky130_fd_sc_hd__o21a_2 _10477_ (.A1(_01985_),
    .A2(_01983_),
    .B1(_01982_),
    .X(_02179_));
 sky130_fd_sc_hd__o31a_1 _10478_ (.A1(net153),
    .A2(_00361_),
    .A3(_00363_),
    .B1(_01944_),
    .X(_02180_));
 sky130_fd_sc_hd__or4_1 _10479_ (.A(net153),
    .B(_00361_),
    .C(_00363_),
    .D(_01944_),
    .X(_02181_));
 sky130_fd_sc_hd__and2b_1 _10480_ (.A_N(_02180_),
    .B(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__a2111oi_1 _10481_ (.A1(net174),
    .A2(_00530_),
    .B1(_02182_),
    .C1(_06331_),
    .D1(_00527_),
    .Y(_02183_));
 sky130_fd_sc_hd__o21a_1 _10482_ (.A1(_06331_),
    .A2(_00532_),
    .B1(_02182_),
    .X(_02184_));
 sky130_fd_sc_hd__or2_2 _10483_ (.A(_02183_),
    .B(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__a31o_1 _10484_ (.A1(_01731_),
    .A2(_01939_),
    .A3(_01940_),
    .B1(_01956_),
    .X(_02186_));
 sky130_fd_sc_hd__and3_1 _10485_ (.A(_07513_),
    .B(_00189_),
    .C(_00191_),
    .X(_02187_));
 sky130_fd_sc_hd__o32a_1 _10486_ (.A1(_00005_),
    .A2(_00007_),
    .A3(_00071_),
    .B1(_00192_),
    .B2(_07512_),
    .X(_02189_));
 sky130_fd_sc_hd__and3_1 _10487_ (.A(_02187_),
    .B(_00072_),
    .C(_00010_),
    .X(_02190_));
 sky130_fd_sc_hd__or4_1 _10488_ (.A(_07512_),
    .B(_00009_),
    .C(_00071_),
    .D(_00192_),
    .X(_02191_));
 sky130_fd_sc_hd__and4_1 _10489_ (.A(_07200_),
    .B(_00429_),
    .C(_07440_),
    .D(_00275_),
    .X(_02192_));
 sky130_fd_sc_hd__nand4_1 _10490_ (.A(_07200_),
    .B(_00429_),
    .C(_07440_),
    .D(_00275_),
    .Y(_02193_));
 sky130_fd_sc_hd__a32o_1 _10491_ (.A1(_07200_),
    .A2(_00425_),
    .A3(_00427_),
    .B1(_00275_),
    .B2(_07440_),
    .X(_02194_));
 sky130_fd_sc_hd__a221o_1 _10492_ (.A1(_07534_),
    .A2(_07535_),
    .B1(_02193_),
    .B2(_02194_),
    .C1(net143),
    .X(_02195_));
 sky130_fd_sc_hd__o211ai_1 _10493_ (.A1(_07539_),
    .A2(net143),
    .B1(_02193_),
    .C1(_02194_),
    .Y(_02196_));
 sky130_fd_sc_hd__o211a_1 _10494_ (.A1(_02189_),
    .A2(_02190_),
    .B1(_02195_),
    .C1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__a211oi_1 _10495_ (.A1(_02195_),
    .A2(_02196_),
    .B1(_02189_),
    .C1(_02190_),
    .Y(_02198_));
 sky130_fd_sc_hd__a31o_1 _10496_ (.A1(_01949_),
    .A2(_07440_),
    .A3(_00150_),
    .B1(_01946_),
    .X(_02200_));
 sky130_fd_sc_hd__o21ai_1 _10497_ (.A1(_02197_),
    .A2(_02198_),
    .B1(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__or3_1 _10498_ (.A(_02197_),
    .B(_02200_),
    .C(_02198_),
    .X(_02202_));
 sky130_fd_sc_hd__nand2_1 _10499_ (.A(_02201_),
    .B(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__o31ai_2 _10500_ (.A1(_05425_),
    .A2(_00532_),
    .A3(_01965_),
    .B1(_01967_),
    .Y(_02204_));
 sky130_fd_sc_hd__a21boi_2 _10501_ (.A1(_01726_),
    .A2(_01953_),
    .B1_N(_01952_),
    .Y(_02205_));
 sky130_fd_sc_hd__xnor2_1 _10502_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__xnor2_1 _10503_ (.A(_02203_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__a21oi_1 _10504_ (.A1(_01942_),
    .A2(_02186_),
    .B1(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__and3_1 _10505_ (.A(_02207_),
    .B(_02186_),
    .C(_01942_),
    .X(_02209_));
 sky130_fd_sc_hd__o21ai_1 _10506_ (.A1(_02208_),
    .A2(_02209_),
    .B1(_02185_),
    .Y(_02211_));
 sky130_fd_sc_hd__or3_1 _10507_ (.A(_02185_),
    .B(_02208_),
    .C(_02209_),
    .X(_02212_));
 sky130_fd_sc_hd__o21ba_1 _10508_ (.A1(_02185_),
    .A2(_02209_),
    .B1_N(_02208_),
    .X(_02213_));
 sky130_fd_sc_hd__nand2_1 _10509_ (.A(_02211_),
    .B(_02212_),
    .Y(_02214_));
 sky130_fd_sc_hd__or2_1 _10510_ (.A(_01962_),
    .B(_01971_),
    .X(_02215_));
 sky130_fd_sc_hd__and3_1 _10511_ (.A(_02214_),
    .B(_02215_),
    .C(_01961_),
    .X(_02216_));
 sky130_fd_sc_hd__a211o_1 _10512_ (.A1(_01971_),
    .A2(_01961_),
    .B1(_01962_),
    .C1(_02214_),
    .X(_02217_));
 sky130_fd_sc_hd__and2b_1 _10513_ (.A_N(_02216_),
    .B(_02217_),
    .X(_02218_));
 sky130_fd_sc_hd__a21bo_2 _10514_ (.A1(_01976_),
    .A2(_01978_),
    .B1_N(_01975_),
    .X(_02219_));
 sky130_fd_sc_hd__xnor2_4 _10515_ (.A(_02218_),
    .B(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand2_4 _10516_ (.A(_02220_),
    .B(_02179_),
    .Y(_02222_));
 sky130_fd_sc_hd__or2_2 _10517_ (.A(_02179_),
    .B(_02220_),
    .X(_02223_));
 sky130_fd_sc_hd__and2_1 _10518_ (.A(_02222_),
    .B(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__nand2_1 _10519_ (.A(_02222_),
    .B(_02223_),
    .Y(_02225_));
 sky130_fd_sc_hd__o211ai_4 _10520_ (.A1(_01992_),
    .A2(_01986_),
    .B1(_01770_),
    .C1(_01995_),
    .Y(_02226_));
 sky130_fd_sc_hd__o211ai_2 _10521_ (.A1(_01766_),
    .A2(_01768_),
    .B1(_01990_),
    .C1(_01996_),
    .Y(_02227_));
 sky130_fd_sc_hd__o211ai_1 _10522_ (.A1(_01937_),
    .A2(_01988_),
    .B1(_02225_),
    .C1(_02226_),
    .Y(_02228_));
 sky130_fd_sc_hd__o211ai_1 _10523_ (.A1(_01938_),
    .A2(_01989_),
    .B1(_02224_),
    .C1(_02227_),
    .Y(_02229_));
 sky130_fd_sc_hd__o2111ai_1 _10524_ (.A1(_01937_),
    .A2(_01988_),
    .B1(_02222_),
    .C1(_02223_),
    .D1(_02226_),
    .Y(_02230_));
 sky130_fd_sc_hd__o211ai_1 _10525_ (.A1(_01938_),
    .A2(_01989_),
    .B1(_02225_),
    .C1(_02227_),
    .Y(_02231_));
 sky130_fd_sc_hd__nand3_2 _10526_ (.A(_02230_),
    .B(_02231_),
    .C(_02178_),
    .Y(_02233_));
 sky130_fd_sc_hd__nand3b_2 _10527_ (.A_N(_02178_),
    .B(_02228_),
    .C(_02229_),
    .Y(_02234_));
 sky130_fd_sc_hd__nor4_4 _10528_ (.A(net13),
    .B(_02047_),
    .C(net16),
    .D(_01397_),
    .Y(_02235_));
 sky130_fd_sc_hd__o211ai_4 _10529_ (.A1(net16),
    .A2(_02048_),
    .B1(net17),
    .C1(net174),
    .Y(_02236_));
 sky130_fd_sc_hd__o21bai_4 _10530_ (.A1(_00321_),
    .A2(_02235_),
    .B1_N(net17),
    .Y(_02237_));
 sky130_fd_sc_hd__o21ai_4 _10531_ (.A1(_00321_),
    .A2(_02235_),
    .B1(net17),
    .Y(_02238_));
 sky130_fd_sc_hd__or3_4 _10532_ (.A(_00321_),
    .B(net17),
    .C(_02235_),
    .X(_02239_));
 sky130_fd_sc_hd__nand2_8 _10533_ (.A(_02238_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_8 _10534_ (.A(net139),
    .B(_02237_),
    .Y(_02241_));
 sky130_fd_sc_hd__a21o_1 _10535_ (.A1(_02238_),
    .A2(_02239_),
    .B1(_00310_),
    .X(_02242_));
 sky130_fd_sc_hd__and3_1 _10536_ (.A(_05436_),
    .B(_00565_),
    .C(_00566_),
    .X(_02244_));
 sky130_fd_sc_hd__o311ai_2 _10537_ (.A1(_01835_),
    .A2(_01840_),
    .A3(_01836_),
    .B1(_02069_),
    .C1(_02067_),
    .Y(_02245_));
 sky130_fd_sc_hd__o41a_1 _10538_ (.A1(_01819_),
    .A2(_02004_),
    .A3(_02062_),
    .A4(_02063_),
    .B1(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__nand4_4 _10539_ (.A(_02050_),
    .B(_02052_),
    .C(_02055_),
    .D(net33),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_2 _10540_ (.A(_02031_),
    .B(_01798_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand4_4 _10541_ (.A(_02033_),
    .B(_02056_),
    .C(_02247_),
    .D(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__a22oi_2 _10542_ (.A1(_02056_),
    .A2(_02247_),
    .B1(_02248_),
    .B2(_02033_),
    .Y(_02250_));
 sky130_fd_sc_hd__a22o_1 _10543_ (.A1(_02056_),
    .A2(_02247_),
    .B1(_02248_),
    .B2(_02033_),
    .X(_02251_));
 sky130_fd_sc_hd__or4_1 _10544_ (.A(_01576_),
    .B(_01598_),
    .C(_01584_),
    .D(_01586_),
    .X(_02252_));
 sky130_fd_sc_hd__o31ai_4 _10545_ (.A1(_01620_),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_02017_),
    .Y(_02253_));
 sky130_fd_sc_hd__and4_1 _10546_ (.A(net137),
    .B(_01590_),
    .C(_01631_),
    .D(_02133_),
    .X(_02255_));
 sky130_fd_sc_hd__nand4b_4 _10547_ (.A_N(_02015_),
    .B(_01588_),
    .C(_01585_),
    .D(_02133_),
    .Y(_02256_));
 sky130_fd_sc_hd__o31a_1 _10548_ (.A1(_02122_),
    .A2(_02015_),
    .A3(_01589_),
    .B1(_02253_),
    .X(_02257_));
 sky130_fd_sc_hd__o211ai_2 _10549_ (.A1(net168),
    .A2(net163),
    .B1(net145),
    .C1(_01220_),
    .Y(_02258_));
 sky130_fd_sc_hd__a31oi_2 _10550_ (.A1(_01053_),
    .A2(net10),
    .A3(net174),
    .B1(net155),
    .Y(_02259_));
 sky130_fd_sc_hd__nand2_4 _10551_ (.A(_01055_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__a31o_1 _10552_ (.A1(_01053_),
    .A2(net10),
    .A3(net174),
    .B1(net158),
    .X(_02261_));
 sky130_fd_sc_hd__o32a_1 _10553_ (.A1(net158),
    .A2(_01054_),
    .A3(_01056_),
    .B1(net155),
    .B2(_00903_),
    .X(_02262_));
 sky130_fd_sc_hd__o21ai_2 _10554_ (.A1(_01054_),
    .A2(_02261_),
    .B1(_02022_),
    .Y(_02263_));
 sky130_fd_sc_hd__o211ai_2 _10555_ (.A1(_01054_),
    .A2(_02261_),
    .B1(_04726_),
    .C1(_00904_),
    .Y(_02264_));
 sky130_fd_sc_hd__nand4_1 _10556_ (.A(net156),
    .B(_01055_),
    .C(_01057_),
    .D(_02022_),
    .Y(_02266_));
 sky130_fd_sc_hd__nand3_2 _10557_ (.A(_02258_),
    .B(_02264_),
    .C(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__o2111ai_4 _10558_ (.A1(_01797_),
    .A2(_02260_),
    .B1(_02263_),
    .C1(_01222_),
    .D1(_02866_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand4_1 _10559_ (.A(_02866_),
    .B(_01222_),
    .C(_02264_),
    .D(_02266_),
    .Y(_02269_));
 sky130_fd_sc_hd__o221ai_1 _10560_ (.A1(_01797_),
    .A2(_02260_),
    .B1(net159),
    .B2(_01221_),
    .C1(_02263_),
    .Y(_02270_));
 sky130_fd_sc_hd__nand2_1 _10561_ (.A(_02269_),
    .B(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hd__nand4_4 _10562_ (.A(_02253_),
    .B(_02256_),
    .C(_02267_),
    .D(_02268_),
    .Y(_02272_));
 sky130_fd_sc_hd__a22oi_2 _10563_ (.A1(_02253_),
    .A2(_02256_),
    .B1(_02267_),
    .B2(_02268_),
    .Y(_02273_));
 sky130_fd_sc_hd__a22o_1 _10564_ (.A1(_02253_),
    .A2(_02256_),
    .B1(_02267_),
    .B2(_02268_),
    .X(_02274_));
 sky130_fd_sc_hd__and3_1 _10565_ (.A(_02866_),
    .B(net141),
    .C(_02021_),
    .X(_02275_));
 sky130_fd_sc_hd__a31oi_4 _10566_ (.A1(_02866_),
    .A2(net141),
    .A3(_02021_),
    .B1(_02023_),
    .Y(_02277_));
 sky130_fd_sc_hd__and3_1 _10567_ (.A(_02272_),
    .B(_02274_),
    .C(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__nand3_1 _10568_ (.A(_02272_),
    .B(_02274_),
    .C(_02277_),
    .Y(_02279_));
 sky130_fd_sc_hd__o2bb2a_1 _10569_ (.A1_N(_02272_),
    .A2_N(_02274_),
    .B1(_02275_),
    .B2(_02023_),
    .X(_02280_));
 sky130_fd_sc_hd__a21o_1 _10570_ (.A1(_02272_),
    .A2(_02274_),
    .B1(_02277_),
    .X(_02281_));
 sky130_fd_sc_hd__o211a_1 _10571_ (.A1(_02023_),
    .A2(_02275_),
    .B1(_02274_),
    .C1(_02272_),
    .X(_02282_));
 sky130_fd_sc_hd__a211oi_1 _10572_ (.A1(_02272_),
    .A2(_02274_),
    .B1(_02275_),
    .C1(_02023_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _10573_ (.A(_02279_),
    .B(_02281_),
    .Y(_02284_));
 sky130_fd_sc_hd__o211ai_1 _10574_ (.A1(_02278_),
    .A2(_02280_),
    .B1(_02249_),
    .C1(_02251_),
    .Y(_02285_));
 sky130_fd_sc_hd__o2bb2ai_1 _10575_ (.A1_N(_02249_),
    .A2_N(_02251_),
    .B1(_02282_),
    .B2(_02283_),
    .Y(_02286_));
 sky130_fd_sc_hd__o2bb2ai_1 _10576_ (.A1_N(_02249_),
    .A2_N(_02251_),
    .B1(_02278_),
    .B2(_02280_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand4_1 _10577_ (.A(_02249_),
    .B(_02251_),
    .C(_02279_),
    .D(_02281_),
    .Y(_02289_));
 sky130_fd_sc_hd__a31o_1 _10578_ (.A1(_02010_),
    .A2(_02034_),
    .A3(_02036_),
    .B1(_02011_),
    .X(_02290_));
 sky130_fd_sc_hd__a31o_1 _10579_ (.A1(_02012_),
    .A2(_02037_),
    .A3(_02038_),
    .B1(_02009_),
    .X(_02291_));
 sky130_fd_sc_hd__nand3_2 _10580_ (.A(_02288_),
    .B(_02289_),
    .C(_02290_),
    .Y(_02292_));
 sky130_fd_sc_hd__inv_2 _10581_ (.A(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__nand3_2 _10582_ (.A(_02285_),
    .B(_02286_),
    .C(_02291_),
    .Y(_02294_));
 sky130_fd_sc_hd__o32a_1 _10583_ (.A1(_02122_),
    .A2(_01406_),
    .A3(_01791_),
    .B1(_01822_),
    .B2(_01292_),
    .X(_02295_));
 sky130_fd_sc_hd__o21ai_1 _10584_ (.A1(_01292_),
    .A2(_01822_),
    .B1(_02018_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor4_4 _10585_ (.A(_01292_),
    .B(_01791_),
    .C(_02017_),
    .D(_01822_),
    .Y(_02297_));
 sky130_fd_sc_hd__or2_1 _10586_ (.A(_02295_),
    .B(_02297_),
    .X(_02299_));
 sky130_fd_sc_hd__o32a_2 _10587_ (.A1(_00900_),
    .A2(_02049_),
    .A3(_02051_),
    .B1(_02295_),
    .B2(_02297_),
    .X(_02300_));
 sky130_fd_sc_hd__and4b_2 _10588_ (.A_N(_02299_),
    .B(_02052_),
    .C(_02050_),
    .D(_00911_),
    .X(_02301_));
 sky130_fd_sc_hd__o221a_1 _10589_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_02295_),
    .B2(_02297_),
    .C1(_02054_),
    .X(_02302_));
 sky130_fd_sc_hd__a21oi_1 _10590_ (.A1(_00911_),
    .A2(_02054_),
    .B1(_02299_),
    .Y(_02303_));
 sky130_fd_sc_hd__o2bb2ai_1 _10591_ (.A1_N(_02292_),
    .A2_N(_02294_),
    .B1(_02302_),
    .B2(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__o21ai_1 _10592_ (.A1(_02300_),
    .A2(_02301_),
    .B1(_02294_),
    .Y(_02305_));
 sky130_fd_sc_hd__o211ai_1 _10593_ (.A1(_02300_),
    .A2(_02301_),
    .B1(_02292_),
    .C1(_02294_),
    .Y(_02306_));
 sky130_fd_sc_hd__a21boi_1 _10594_ (.A1(_02044_),
    .A2(_02060_),
    .B1_N(_02043_),
    .Y(_02307_));
 sky130_fd_sc_hd__a21o_1 _10595_ (.A1(_02304_),
    .A2(_02306_),
    .B1(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__o211ai_2 _10596_ (.A1(_02305_),
    .A2(_02293_),
    .B1(_02304_),
    .C1(_02307_),
    .Y(_02310_));
 sky130_fd_sc_hd__o211ai_2 _10597_ (.A1(_02064_),
    .A2(_02062_),
    .B1(_02310_),
    .C1(_02245_),
    .Y(_02311_));
 sky130_fd_sc_hd__and3_1 _10598_ (.A(_02246_),
    .B(_02308_),
    .C(_02310_),
    .X(_02312_));
 sky130_fd_sc_hd__a21o_1 _10599_ (.A1(_02308_),
    .A2(_02310_),
    .B1(_02246_),
    .X(_02313_));
 sky130_fd_sc_hd__and2b_1 _10600_ (.A_N(_02312_),
    .B(_02313_),
    .X(_02314_));
 sky130_fd_sc_hd__a21oi_1 _10601_ (.A1(_05436_),
    .A2(_00569_),
    .B1(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__a31o_1 _10602_ (.A1(_05392_),
    .A2(_05414_),
    .A3(_00569_),
    .B1(_02314_),
    .X(_02316_));
 sky130_fd_sc_hd__and3_1 _10603_ (.A(_02314_),
    .B(_05436_),
    .C(_00569_),
    .X(_02317_));
 sky130_fd_sc_hd__a41o_1 _10604_ (.A1(_05436_),
    .A2(net147),
    .A3(net146),
    .A4(_02314_),
    .B1(_02315_),
    .X(_02318_));
 sky130_fd_sc_hd__a21oi_1 _10605_ (.A1(net33),
    .A2(_02240_),
    .B1(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__and3_1 _10606_ (.A(_02318_),
    .B(_02240_),
    .C(net33),
    .X(_02321_));
 sky130_fd_sc_hd__and4b_1 _10607_ (.A_N(_02317_),
    .B(_02240_),
    .C(net33),
    .D(_02316_),
    .X(_02322_));
 sky130_fd_sc_hd__o21a_1 _10608_ (.A1(_00310_),
    .A2(_02241_),
    .B1(_02318_),
    .X(_02323_));
 sky130_fd_sc_hd__nor2_1 _10609_ (.A(_02322_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__o211ai_1 _10610_ (.A1(_02319_),
    .A2(_02321_),
    .B1(_02233_),
    .C1(_02234_),
    .Y(_02325_));
 sky130_fd_sc_hd__a21o_1 _10611_ (.A1(_02233_),
    .A2(_02234_),
    .B1(_02324_),
    .X(_02326_));
 sky130_fd_sc_hd__o2bb2ai_1 _10612_ (.A1_N(_02233_),
    .A2_N(_02234_),
    .B1(_02319_),
    .B2(_02321_),
    .Y(_02327_));
 sky130_fd_sc_hd__o211ai_1 _10613_ (.A1(_02322_),
    .A2(_02323_),
    .B1(_02233_),
    .C1(_02234_),
    .Y(_02328_));
 sky130_fd_sc_hd__nand2_1 _10614_ (.A(_02327_),
    .B(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _10615_ (.A(_02325_),
    .B(_02326_),
    .Y(_02330_));
 sky130_fd_sc_hd__and2_1 _10616_ (.A(_02001_),
    .B(_02075_),
    .X(_02332_));
 sky130_fd_sc_hd__nand2_1 _10617_ (.A(_02001_),
    .B(_02075_),
    .Y(_02333_));
 sky130_fd_sc_hd__a22o_1 _10618_ (.A1(_02001_),
    .A2(_02075_),
    .B1(_02327_),
    .B2(_02328_),
    .X(_02334_));
 sky130_fd_sc_hd__a21o_1 _10619_ (.A1(_02325_),
    .A2(_02326_),
    .B1(_02333_),
    .X(_02335_));
 sky130_fd_sc_hd__o211ai_2 _10620_ (.A1(_01646_),
    .A2(_01853_),
    .B1(_02080_),
    .C1(_02081_),
    .Y(_02336_));
 sky130_fd_sc_hd__nand4_1 _10621_ (.A(_02078_),
    .B(_02334_),
    .C(_02335_),
    .D(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__a22o_1 _10622_ (.A1(_02334_),
    .A2(_02335_),
    .B1(_02336_),
    .B2(_02078_),
    .X(_02338_));
 sky130_fd_sc_hd__nand2_1 _10623_ (.A(_02337_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__a311o_1 _10624_ (.A1(_01645_),
    .A2(_01861_),
    .A3(_02084_),
    .B1(_02339_),
    .C1(_00834_),
    .X(_02340_));
 sky130_fd_sc_hd__a2bb2o_1 _10625_ (.A1_N(_00834_),
    .A2_N(_02085_),
    .B1(_02337_),
    .B2(_02338_),
    .X(_02341_));
 sky130_fd_sc_hd__and2_1 _10626_ (.A(_02340_),
    .B(_02341_),
    .X(net81));
 sky130_fd_sc_hd__and4_1 _10627_ (.A(_01645_),
    .B(_01861_),
    .C(_02339_),
    .D(_02084_),
    .X(_02343_));
 sky130_fd_sc_hd__a21bo_1 _10628_ (.A1(_02233_),
    .A2(_02324_),
    .B1_N(_02234_),
    .X(_02344_));
 sky130_fd_sc_hd__a32o_1 _10629_ (.A1(_02314_),
    .A2(_05436_),
    .A3(_00569_),
    .B1(_02240_),
    .B2(net33),
    .X(_02345_));
 sky130_fd_sc_hd__a31o_1 _10630_ (.A1(_02316_),
    .A2(_02240_),
    .A3(net33),
    .B1(_02317_),
    .X(_02346_));
 sky130_fd_sc_hd__nor2_4 _10631_ (.A(net16),
    .B(net17),
    .Y(_02347_));
 sky130_fd_sc_hd__or2_1 _10632_ (.A(net16),
    .B(net17),
    .X(_02348_));
 sky130_fd_sc_hd__nand4_4 _10633_ (.A(_01581_),
    .B(_02347_),
    .C(_00693_),
    .D(_00715_),
    .Y(_02349_));
 sky130_fd_sc_hd__a311oi_4 _10634_ (.A1(_01581_),
    .A2(_02045_),
    .A3(_02347_),
    .B1(net18),
    .C1(_00321_),
    .Y(_02350_));
 sky130_fd_sc_hd__a21boi_4 _10635_ (.A1(_02349_),
    .A2(net174),
    .B1_N(net18),
    .Y(_02351_));
 sky130_fd_sc_hd__o311a_4 _10636_ (.A1(_01582_),
    .A2(_02047_),
    .A3(_02348_),
    .B1(net18),
    .C1(net174),
    .X(_02353_));
 sky130_fd_sc_hd__a21oi_4 _10637_ (.A1(_02349_),
    .A2(net174),
    .B1(net18),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_8 _10638_ (.A(_02350_),
    .B(_02351_),
    .Y(_02355_));
 sky130_fd_sc_hd__nor2_8 _10639_ (.A(_02353_),
    .B(_02354_),
    .Y(_02356_));
 sky130_fd_sc_hd__or4_4 _10640_ (.A(_00310_),
    .B(_00900_),
    .C(_02241_),
    .D(_02355_),
    .X(_02357_));
 sky130_fd_sc_hd__a32o_1 _10641_ (.A1(_00911_),
    .A2(net139),
    .A3(_02237_),
    .B1(_02356_),
    .B2(net33),
    .X(_02358_));
 sky130_fd_sc_hd__o31a_2 _10642_ (.A1(_00900_),
    .A2(_02355_),
    .A3(_02242_),
    .B1(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__o32a_1 _10643_ (.A1(_05425_),
    .A2(_00898_),
    .A3(_00901_),
    .B1(_06331_),
    .B2(_00570_),
    .X(_02360_));
 sky130_fd_sc_hd__and3_1 _10644_ (.A(_02244_),
    .B(_00904_),
    .C(_06341_),
    .X(_02361_));
 sky130_fd_sc_hd__or4_2 _10645_ (.A(_05425_),
    .B(_06331_),
    .C(_00570_),
    .D(_00903_),
    .X(_02362_));
 sky130_fd_sc_hd__a31o_1 _10646_ (.A1(_06341_),
    .A2(_00904_),
    .A3(_02244_),
    .B1(_02360_),
    .X(_02364_));
 sky130_fd_sc_hd__o31ai_4 _10647_ (.A1(_02293_),
    .A2(_02300_),
    .A3(_02301_),
    .B1(_02294_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _10648_ (.A(_02292_),
    .B(_02305_),
    .Y(_02366_));
 sky130_fd_sc_hd__or3_4 _10649_ (.A(_01292_),
    .B(_02049_),
    .C(_02051_),
    .X(_02367_));
 sky130_fd_sc_hd__or4_2 _10650_ (.A(_02210_),
    .B(_01584_),
    .C(_01586_),
    .D(_01822_),
    .X(_02368_));
 sky130_fd_sc_hd__o32a_2 _10651_ (.A1(_02122_),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(_01620_),
    .X(_02369_));
 sky130_fd_sc_hd__a31o_1 _10652_ (.A1(_02199_),
    .A2(_01590_),
    .A3(_01823_),
    .B1(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__xnor2_4 _10653_ (.A(_02367_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__o21ai_1 _10654_ (.A1(_02282_),
    .A2(_02283_),
    .B1(_02251_),
    .Y(_02372_));
 sky130_fd_sc_hd__o211a_1 _10655_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_02054_),
    .C1(_02296_),
    .X(_02373_));
 sky130_fd_sc_hd__a31oi_2 _10656_ (.A1(_00911_),
    .A2(_02054_),
    .A3(_02296_),
    .B1(_02297_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand2_1 _10657_ (.A(_02272_),
    .B(_02277_),
    .Y(_02376_));
 sky130_fd_sc_hd__o211ai_4 _10658_ (.A1(_02273_),
    .A2(_02277_),
    .B1(_02375_),
    .C1(_02272_),
    .Y(_02377_));
 sky130_fd_sc_hd__o221a_1 _10659_ (.A1(_02257_),
    .A2(_02271_),
    .B1(_02297_),
    .B2(_02373_),
    .C1(_02376_),
    .X(_02378_));
 sky130_fd_sc_hd__o221ai_4 _10660_ (.A1(_02257_),
    .A2(_02271_),
    .B1(_02297_),
    .B2(_02373_),
    .C1(_02376_),
    .Y(_02379_));
 sky130_fd_sc_hd__o32a_1 _10661_ (.A1(net158),
    .A2(_02022_),
    .A3(_01058_),
    .B1(net159),
    .B2(_01221_),
    .X(_02380_));
 sky130_fd_sc_hd__o32ai_1 _10662_ (.A1(net158),
    .A2(_00903_),
    .A3(_02260_),
    .B1(_02258_),
    .B2(_02262_),
    .Y(_02381_));
 sky130_fd_sc_hd__o221a_1 _10663_ (.A1(net168),
    .A2(net163),
    .B1(_01396_),
    .B2(_01403_),
    .C1(_01400_),
    .X(_02382_));
 sky130_fd_sc_hd__o31ai_4 _10664_ (.A1(net158),
    .A2(_01217_),
    .A3(_01219_),
    .B1(_02260_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand3b_1 _10665_ (.A_N(_02260_),
    .B(_01222_),
    .C(net156),
    .Y(_02384_));
 sky130_fd_sc_hd__a31o_1 _10666_ (.A1(net156),
    .A2(net145),
    .A3(_01220_),
    .B1(_02260_),
    .X(_02386_));
 sky130_fd_sc_hd__nand4_2 _10667_ (.A(net156),
    .B(net145),
    .C(_01220_),
    .D(_02260_),
    .Y(_02387_));
 sky130_fd_sc_hd__o211ai_1 _10668_ (.A1(net136),
    .A2(net159),
    .B1(_02387_),
    .C1(_02386_),
    .Y(_02388_));
 sky130_fd_sc_hd__o2111ai_1 _10669_ (.A1(net168),
    .A2(net163),
    .B1(net137),
    .C1(_02383_),
    .D1(_02384_),
    .Y(_02389_));
 sky130_fd_sc_hd__o2111ai_4 _10670_ (.A1(net168),
    .A2(net163),
    .B1(_02387_),
    .C1(net137),
    .D1(_02386_),
    .Y(_02390_));
 sky130_fd_sc_hd__o211ai_2 _10671_ (.A1(net159),
    .A2(net136),
    .B1(_02383_),
    .C1(_02384_),
    .Y(_02391_));
 sky130_fd_sc_hd__o211ai_4 _10672_ (.A1(_02262_),
    .A2(_02380_),
    .B1(_02390_),
    .C1(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__nand3_2 _10673_ (.A(_02381_),
    .B(_02388_),
    .C(_02389_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand3_2 _10674_ (.A(_02392_),
    .B(_02393_),
    .C(_02255_),
    .Y(_02394_));
 sky130_fd_sc_hd__o2bb2ai_2 _10675_ (.A1_N(_02392_),
    .A2_N(_02393_),
    .B1(_02017_),
    .B2(_02252_),
    .Y(_02395_));
 sky130_fd_sc_hd__a22o_1 _10676_ (.A1(_02377_),
    .A2(_02379_),
    .B1(_02394_),
    .B2(_02395_),
    .X(_02397_));
 sky130_fd_sc_hd__nand4_4 _10677_ (.A(_02377_),
    .B(_02379_),
    .C(_02394_),
    .D(_02395_),
    .Y(_02398_));
 sky130_fd_sc_hd__a22oi_4 _10678_ (.A1(_02249_),
    .A2(_02372_),
    .B1(_02397_),
    .B2(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__o2111a_2 _10679_ (.A1(_02284_),
    .A2(_02250_),
    .B1(_02249_),
    .C1(_02398_),
    .D1(_02397_),
    .X(_02400_));
 sky130_fd_sc_hd__o2111ai_2 _10680_ (.A1(_02284_),
    .A2(_02250_),
    .B1(_02249_),
    .C1(_02398_),
    .D1(_02397_),
    .Y(_02401_));
 sky130_fd_sc_hd__o21ai_2 _10681_ (.A1(_02399_),
    .A2(_02400_),
    .B1(_02371_),
    .Y(_02402_));
 sky130_fd_sc_hd__a21oi_1 _10682_ (.A1(_02371_),
    .A2(_02401_),
    .B1(_02399_),
    .Y(_02403_));
 sky130_fd_sc_hd__o31a_1 _10683_ (.A1(_02371_),
    .A2(_02399_),
    .A3(_02400_),
    .B1(_02402_),
    .X(_02404_));
 sky130_fd_sc_hd__o31ai_2 _10684_ (.A1(_02371_),
    .A2(_02399_),
    .A3(_02400_),
    .B1(_02402_),
    .Y(_02405_));
 sky130_fd_sc_hd__o311ai_2 _10685_ (.A1(_02371_),
    .A2(_02399_),
    .A3(_02400_),
    .B1(_02402_),
    .C1(_02365_),
    .Y(_02406_));
 sky130_fd_sc_hd__nand2_1 _10686_ (.A(_02366_),
    .B(_02405_),
    .Y(_02408_));
 sky130_fd_sc_hd__nand4_1 _10687_ (.A(_02308_),
    .B(_02311_),
    .C(_02406_),
    .D(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__a22o_1 _10688_ (.A1(_02308_),
    .A2(_02311_),
    .B1(_02406_),
    .B2(_02408_),
    .X(_02410_));
 sky130_fd_sc_hd__o211a_1 _10689_ (.A1(_02360_),
    .A2(_02361_),
    .B1(_02409_),
    .C1(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__a21oi_2 _10690_ (.A1(_02409_),
    .A2(_02410_),
    .B1(_02364_),
    .Y(_02412_));
 sky130_fd_sc_hd__nor2_1 _10691_ (.A(_02411_),
    .B(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__o21bai_2 _10692_ (.A1(_02411_),
    .A2(_02412_),
    .B1_N(_02359_),
    .Y(_02414_));
 sky130_fd_sc_hd__nand2_1 _10693_ (.A(_02359_),
    .B(_02413_),
    .Y(_02415_));
 sky130_fd_sc_hd__and3_1 _10694_ (.A(_02346_),
    .B(_02414_),
    .C(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__nand4_1 _10695_ (.A(_02316_),
    .B(_02345_),
    .C(_02414_),
    .D(_02415_),
    .Y(_02417_));
 sky130_fd_sc_hd__a21oi_1 _10696_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_02346_),
    .Y(_02419_));
 sky130_fd_sc_hd__a41o_1 _10697_ (.A1(_02316_),
    .A2(_02345_),
    .A3(_02414_),
    .A4(_02415_),
    .B1(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__inv_2 _10698_ (.A(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__o32ai_4 _10699_ (.A1(_02098_),
    .A2(_02172_),
    .A3(_02173_),
    .B1(_02086_),
    .B2(_02175_),
    .Y(_02422_));
 sky130_fd_sc_hd__o32a_1 _10700_ (.A1(_07146_),
    .A2(_07168_),
    .A3(_00580_),
    .B1(_00744_),
    .B2(_05327_),
    .X(_02423_));
 sky130_fd_sc_hd__and4_1 _10701_ (.A(_07200_),
    .B(_00743_),
    .C(_00581_),
    .D(_05316_),
    .X(_02424_));
 sky130_fd_sc_hd__nor2_1 _10702_ (.A(_02423_),
    .B(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__nor4_1 _10703_ (.A(net46),
    .B(_02088_),
    .C(net49),
    .D(_01535_),
    .Y(_02426_));
 sky130_fd_sc_hd__o211ai_4 _10704_ (.A1(net49),
    .A2(_02091_),
    .B1(net50),
    .C1(net173),
    .Y(_02427_));
 sky130_fd_sc_hd__o21bai_4 _10705_ (.A1(_00299_),
    .A2(net138),
    .B1_N(net50),
    .Y(_02428_));
 sky130_fd_sc_hd__o21ai_4 _10706_ (.A1(_00299_),
    .A2(net138),
    .B1(net50),
    .Y(_02430_));
 sky130_fd_sc_hd__or3_4 _10707_ (.A(_00299_),
    .B(net50),
    .C(net138),
    .X(_02431_));
 sky130_fd_sc_hd__nand2_8 _10708_ (.A(_02430_),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_8 _10709_ (.A(_02427_),
    .B(_02428_),
    .Y(_02433_));
 sky130_fd_sc_hd__and4_1 _10710_ (.A(_00998_),
    .B(_02432_),
    .C(_02097_),
    .D(net1),
    .X(_02434_));
 sky130_fd_sc_hd__or4_4 _10711_ (.A(_00288_),
    .B(_00987_),
    .C(_02433_),
    .D(_02096_),
    .X(_02435_));
 sky130_fd_sc_hd__o32a_1 _10712_ (.A1(_00987_),
    .A2(_02092_),
    .A3(_02094_),
    .B1(_02433_),
    .B2(_00288_),
    .X(_02436_));
 sky130_fd_sc_hd__nor2_1 _10713_ (.A(_02434_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__a31o_2 _10714_ (.A1(_04255_),
    .A2(_02102_),
    .A3(_00743_),
    .B1(_02099_),
    .X(_02438_));
 sky130_fd_sc_hd__nand3_4 _10715_ (.A(_02138_),
    .B(_02148_),
    .C(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__a21oi_2 _10716_ (.A1(_02138_),
    .A2(_02148_),
    .B1(_02438_),
    .Y(_02441_));
 sky130_fd_sc_hd__o21bai_4 _10717_ (.A1(_02137_),
    .A2(_02147_),
    .B1_N(_02438_),
    .Y(_02442_));
 sky130_fd_sc_hd__a21oi_1 _10718_ (.A1(_01886_),
    .A2(_02125_),
    .B1(_02131_),
    .Y(_02443_));
 sky130_fd_sc_hd__o21ai_1 _10719_ (.A1(_01667_),
    .A2(_02127_),
    .B1(_02131_),
    .Y(_02444_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_02126_),
    .B(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__a31o_1 _10721_ (.A1(_01535_),
    .A2(net46),
    .A3(net173),
    .B1(_01958_),
    .X(_02446_));
 sky130_fd_sc_hd__and3_1 _10722_ (.A(_01969_),
    .B(_01539_),
    .C(_01541_),
    .X(_02447_));
 sky130_fd_sc_hd__a221o_1 _10723_ (.A1(_01903_),
    .A2(_01925_),
    .B1(_01535_),
    .B2(_01537_),
    .C1(_01540_),
    .X(_02448_));
 sky130_fd_sc_hd__o211ai_2 _10724_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_01659_),
    .C1(net140),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_4 _10725_ (.A(_02127_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__o221a_1 _10726_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01423_),
    .B2(_01445_),
    .C1(_01172_),
    .X(_02452_));
 sky130_fd_sc_hd__o2111ai_4 _10727_ (.A1(_01095_),
    .A2(_01117_),
    .B1(_01499_),
    .C1(_01659_),
    .D1(net140),
    .Y(_02453_));
 sky130_fd_sc_hd__nand4_1 _10728_ (.A(_01664_),
    .B(net135),
    .C(_01880_),
    .D(_02452_),
    .Y(_02454_));
 sky130_fd_sc_hd__o2111ai_4 _10729_ (.A1(_02453_),
    .A2(_01882_),
    .B1(_01544_),
    .C1(_01969_),
    .D1(_02450_),
    .Y(_02455_));
 sky130_fd_sc_hd__o2bb2ai_2 _10730_ (.A1_N(_02450_),
    .A2_N(_02454_),
    .B1(_01540_),
    .B2(_02446_),
    .Y(_02456_));
 sky130_fd_sc_hd__a21o_1 _10731_ (.A1(_02450_),
    .A2(_02454_),
    .B1(_02448_),
    .X(_02457_));
 sky130_fd_sc_hd__o221ai_4 _10732_ (.A1(_01958_),
    .A2(_01542_),
    .B1(_01882_),
    .B2(_02453_),
    .C1(_02450_),
    .Y(_02458_));
 sky130_fd_sc_hd__o211ai_4 _10733_ (.A1(_02128_),
    .A2(_02443_),
    .B1(_02455_),
    .C1(_02456_),
    .Y(_02459_));
 sky130_fd_sc_hd__a22oi_2 _10734_ (.A1(_02126_),
    .A2(_02444_),
    .B1(_02455_),
    .B2(_02456_),
    .Y(_02460_));
 sky130_fd_sc_hd__nand3_4 _10735_ (.A(_02457_),
    .B(_02458_),
    .C(_02445_),
    .Y(_02461_));
 sky130_fd_sc_hd__nand4_2 _10736_ (.A(_02461_),
    .B(_01871_),
    .C(_02459_),
    .D(_02118_),
    .Y(_02463_));
 sky130_fd_sc_hd__o2bb2ai_1 _10737_ (.A1_N(_02459_),
    .A2_N(_02461_),
    .B1(_01872_),
    .B2(_02117_),
    .Y(_02464_));
 sky130_fd_sc_hd__a21oi_1 _10738_ (.A1(_02459_),
    .A2(_02461_),
    .B1(_02120_),
    .Y(_02465_));
 sky130_fd_sc_hd__a21o_1 _10739_ (.A1(_02459_),
    .A2(_02461_),
    .B1(_02120_),
    .X(_02466_));
 sky130_fd_sc_hd__and3_1 _10740_ (.A(_02120_),
    .B(_02459_),
    .C(_02461_),
    .X(_02467_));
 sky130_fd_sc_hd__o211ai_4 _10741_ (.A1(_01872_),
    .A2(_02117_),
    .B1(_02459_),
    .C1(_02461_),
    .Y(_02468_));
 sky130_fd_sc_hd__o2bb2ai_4 _10742_ (.A1_N(_02439_),
    .A2_N(_02442_),
    .B1(_02465_),
    .B2(_02467_),
    .Y(_02469_));
 sky130_fd_sc_hd__nand4_4 _10743_ (.A(_02439_),
    .B(_02442_),
    .C(_02466_),
    .D(_02468_),
    .Y(_02470_));
 sky130_fd_sc_hd__a31oi_4 _10744_ (.A1(_02116_),
    .A2(_02143_),
    .A3(_02146_),
    .B1(_02114_),
    .Y(_02471_));
 sky130_fd_sc_hd__a21oi_2 _10745_ (.A1(_02469_),
    .A2(_02470_),
    .B1(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__a21o_1 _10746_ (.A1(_02469_),
    .A2(_02470_),
    .B1(_02471_),
    .X(_02474_));
 sky130_fd_sc_hd__o32a_2 _10747_ (.A1(_03906_),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_01272_),
    .B2(_02636_),
    .X(_02475_));
 sky130_fd_sc_hd__a31o_1 _10748_ (.A1(_03917_),
    .A2(_01273_),
    .A3(_02118_),
    .B1(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__and3_1 _10749_ (.A(_04255_),
    .B(_01038_),
    .C(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__a21oi_2 _10750_ (.A1(_04255_),
    .A2(_01038_),
    .B1(_02476_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_1 _10751_ (.A(_02477_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__inv_2 _10752_ (.A(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__nand3_4 _10753_ (.A(_02471_),
    .B(_02470_),
    .C(_02469_),
    .Y(_02481_));
 sky130_fd_sc_hd__a21oi_4 _10754_ (.A1(_02481_),
    .A2(_02480_),
    .B1(_02472_),
    .Y(_02482_));
 sky130_fd_sc_hd__o211ai_4 _10755_ (.A1(_02477_),
    .A2(_02478_),
    .B1(_02481_),
    .C1(_02474_),
    .Y(_02483_));
 sky130_fd_sc_hd__a21o_1 _10756_ (.A1(_02474_),
    .A2(_02481_),
    .B1(_02480_),
    .X(_02485_));
 sky130_fd_sc_hd__a311o_1 _10757_ (.A1(_02469_),
    .A2(_02471_),
    .A3(_02470_),
    .B1(_02480_),
    .C1(_02472_),
    .X(_02486_));
 sky130_fd_sc_hd__a21oi_4 _10758_ (.A1(_02474_),
    .A2(_02481_),
    .B1(_02479_),
    .Y(_02487_));
 sky130_fd_sc_hd__nand2_2 _10759_ (.A(_02483_),
    .B(_02485_),
    .Y(_02488_));
 sky130_fd_sc_hd__o2111ai_4 _10760_ (.A1(_02105_),
    .A2(_02158_),
    .B1(_02161_),
    .C1(_02483_),
    .D1(_02485_),
    .Y(_02489_));
 sky130_fd_sc_hd__nand2_4 _10761_ (.A(_02486_),
    .B(_02162_),
    .Y(_02490_));
 sky130_fd_sc_hd__nand3b_1 _10762_ (.A_N(_02487_),
    .B(_02162_),
    .C(_02486_),
    .Y(_02491_));
 sky130_fd_sc_hd__o211ai_4 _10763_ (.A1(_02168_),
    .A2(_02169_),
    .B1(_01931_),
    .C1(_01933_),
    .Y(_02492_));
 sky130_fd_sc_hd__nand3_1 _10764_ (.A(_01930_),
    .B(_01934_),
    .C(_02170_),
    .Y(_02493_));
 sky130_fd_sc_hd__a22oi_1 _10765_ (.A1(_02489_),
    .A2(_02491_),
    .B1(_02492_),
    .B2(_02170_),
    .Y(_02494_));
 sky130_fd_sc_hd__a22o_1 _10766_ (.A1(_02489_),
    .A2(_02491_),
    .B1(_02492_),
    .B2(_02170_),
    .X(_02496_));
 sky130_fd_sc_hd__o2111a_1 _10767_ (.A1(_02490_),
    .A2(_02487_),
    .B1(_02170_),
    .C1(_02489_),
    .D1(_02492_),
    .X(_02497_));
 sky130_fd_sc_hd__o2111ai_1 _10768_ (.A1(_02490_),
    .A2(_02487_),
    .B1(_02170_),
    .C1(_02489_),
    .D1(_02492_),
    .Y(_02498_));
 sky130_fd_sc_hd__nand3_1 _10769_ (.A(_02496_),
    .B(_02498_),
    .C(_02437_),
    .Y(_02499_));
 sky130_fd_sc_hd__o22ai_2 _10770_ (.A1(_02434_),
    .A2(_02436_),
    .B1(_02494_),
    .B2(_02497_),
    .Y(_02500_));
 sky130_fd_sc_hd__nand2_1 _10771_ (.A(_02499_),
    .B(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__a2bb2o_1 _10772_ (.A1_N(_02423_),
    .A2_N(_02424_),
    .B1(_02499_),
    .B2(_02500_),
    .X(_02502_));
 sky130_fd_sc_hd__nand3_1 _10773_ (.A(_02500_),
    .B(_02425_),
    .C(_02499_),
    .Y(_02503_));
 sky130_fd_sc_hd__o211a_2 _10774_ (.A1(_02423_),
    .A2(_02424_),
    .B1(_02499_),
    .C1(_02500_),
    .X(_02504_));
 sky130_fd_sc_hd__nand3_4 _10775_ (.A(_02422_),
    .B(_02502_),
    .C(_02503_),
    .Y(_02505_));
 sky130_fd_sc_hd__a21o_2 _10776_ (.A1(_02501_),
    .A2(_02425_),
    .B1(_02422_),
    .X(_02507_));
 sky130_fd_sc_hd__o21a_1 _10777_ (.A1(_02504_),
    .A2(_02507_),
    .B1(_02505_),
    .X(_02508_));
 sky130_fd_sc_hd__o211ai_4 _10778_ (.A1(_01937_),
    .A2(_01988_),
    .B1(_02223_),
    .C1(_02226_),
    .Y(_02509_));
 sky130_fd_sc_hd__o211ai_2 _10779_ (.A1(_01938_),
    .A2(_01989_),
    .B1(_02222_),
    .C1(_02227_),
    .Y(_02510_));
 sky130_fd_sc_hd__o21ai_2 _10780_ (.A1(_02179_),
    .A2(_02220_),
    .B1(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__a21o_1 _10781_ (.A1(_02204_),
    .A2(_02205_),
    .B1(_02203_),
    .X(_02512_));
 sky130_fd_sc_hd__o21a_1 _10782_ (.A1(_02204_),
    .A2(_02205_),
    .B1(_02512_),
    .X(_02513_));
 sky130_fd_sc_hd__or3_1 _10783_ (.A(_06331_),
    .B(_00532_),
    .C(_02180_),
    .X(_02514_));
 sky130_fd_sc_hd__nor2_1 _10784_ (.A(_02200_),
    .B(_02198_),
    .Y(_02515_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(_02197_),
    .B(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__a21oi_1 _10786_ (.A1(_02181_),
    .A2(_02514_),
    .B1(_02516_),
    .Y(_02518_));
 sky130_fd_sc_hd__o311a_1 _10787_ (.A1(_06331_),
    .A2(_00532_),
    .A3(_02180_),
    .B1(_02181_),
    .C1(_02516_),
    .X(_02519_));
 sky130_fd_sc_hd__a31o_1 _10788_ (.A1(_07540_),
    .A2(_00150_),
    .A3(_02194_),
    .B1(_02192_),
    .X(_02520_));
 sky130_fd_sc_hd__or4_1 _10789_ (.A(_00067_),
    .B(_00069_),
    .C(_00145_),
    .D(_00147_),
    .X(_02521_));
 sky130_fd_sc_hd__o32a_1 _10790_ (.A1(_07539_),
    .A2(_00270_),
    .A3(_00272_),
    .B1(_07441_),
    .B2(_00428_),
    .X(_02522_));
 sky130_fd_sc_hd__o211a_1 _10791_ (.A1(_00266_),
    .A2(_00268_),
    .B1(_00429_),
    .C1(_07540_),
    .X(_02523_));
 sky130_fd_sc_hd__a21oi_1 _10792_ (.A1(_07440_),
    .A2(_02523_),
    .B1(_02522_),
    .Y(_02524_));
 sky130_fd_sc_hd__xnor2_1 _10793_ (.A(_02521_),
    .B(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__nor2_1 _10794_ (.A(_02520_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__nand2_1 _10795_ (.A(_02525_),
    .B(_02520_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2b_1 _10796_ (.A_N(_02526_),
    .B(_02527_),
    .Y(_02529_));
 sky130_fd_sc_hd__xor2_1 _10797_ (.A(_02190_),
    .B(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__o21a_1 _10798_ (.A1(_02518_),
    .A2(_02519_),
    .B1(_02530_),
    .X(_02531_));
 sky130_fd_sc_hd__nor3_1 _10799_ (.A(_02518_),
    .B(_02519_),
    .C(_02530_),
    .Y(_02532_));
 sky130_fd_sc_hd__nor2_1 _10800_ (.A(_02531_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__o211a_1 _10801_ (.A1(_02204_),
    .A2(_02205_),
    .B1(_02512_),
    .C1(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__or2_1 _10802_ (.A(_02513_),
    .B(_02533_),
    .X(_02535_));
 sky130_fd_sc_hd__xnor2_1 _10803_ (.A(_02513_),
    .B(_02533_),
    .Y(_02536_));
 sky130_fd_sc_hd__and3_1 _10804_ (.A(_02187_),
    .B(_00367_),
    .C(_00010_),
    .X(_02537_));
 sky130_fd_sc_hd__or4_1 _10805_ (.A(_07512_),
    .B(_00009_),
    .C(_00192_),
    .D(_00366_),
    .X(_02538_));
 sky130_fd_sc_hd__o32a_1 _10806_ (.A1(_07512_),
    .A2(_00361_),
    .A3(_00363_),
    .B1(_00009_),
    .B2(_00192_),
    .X(_02539_));
 sky130_fd_sc_hd__o22a_1 _10807_ (.A1(net153),
    .A2(_00532_),
    .B1(_02537_),
    .B2(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__or4_1 _10808_ (.A(net153),
    .B(_00532_),
    .C(_02537_),
    .D(_02539_),
    .X(_02541_));
 sky130_fd_sc_hd__and2b_1 _10809_ (.A_N(_02540_),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__xnor2_2 _10810_ (.A(_02536_),
    .B(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__xnor2_1 _10811_ (.A(_02213_),
    .B(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__a21o_1 _10812_ (.A1(_02217_),
    .A2(_02219_),
    .B1(_02216_),
    .X(_02545_));
 sky130_fd_sc_hd__and2_2 _10813_ (.A(_02544_),
    .B(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__nor2_2 _10814_ (.A(_02545_),
    .B(_02544_),
    .Y(_02547_));
 sky130_fd_sc_hd__or2_2 _10815_ (.A(_02546_),
    .B(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__inv_2 _10816_ (.A(_02548_),
    .Y(_02550_));
 sky130_fd_sc_hd__o211ai_2 _10817_ (.A1(_02179_),
    .A2(_02220_),
    .B1(_02550_),
    .C1(_02510_),
    .Y(_02551_));
 sky130_fd_sc_hd__o211ai_2 _10818_ (.A1(_02546_),
    .A2(_02547_),
    .B1(_02222_),
    .C1(_02509_),
    .Y(_02552_));
 sky130_fd_sc_hd__o2111a_1 _10819_ (.A1(_02507_),
    .A2(_02504_),
    .B1(_02505_),
    .C1(_02551_),
    .D1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__o2111ai_2 _10820_ (.A1(_02507_),
    .A2(_02504_),
    .B1(_02505_),
    .C1(_02551_),
    .D1(_02552_),
    .Y(_02554_));
 sky130_fd_sc_hd__a21oi_1 _10821_ (.A1(_02551_),
    .A2(_02552_),
    .B1(_02508_),
    .Y(_02555_));
 sky130_fd_sc_hd__a21o_1 _10822_ (.A1(_02551_),
    .A2(_02552_),
    .B1(_02508_),
    .X(_02556_));
 sky130_fd_sc_hd__o21ai_1 _10823_ (.A1(_02553_),
    .A2(_02555_),
    .B1(_02421_),
    .Y(_02557_));
 sky130_fd_sc_hd__o211ai_1 _10824_ (.A1(_02416_),
    .A2(_02419_),
    .B1(_02554_),
    .C1(_02556_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand3_1 _10825_ (.A(_02556_),
    .B(_02421_),
    .C(_02554_),
    .Y(_02559_));
 sky130_fd_sc_hd__o22ai_1 _10826_ (.A1(_02416_),
    .A2(_02419_),
    .B1(_02553_),
    .B2(_02555_),
    .Y(_02561_));
 sky130_fd_sc_hd__nand2_1 _10827_ (.A(_02557_),
    .B(_02558_),
    .Y(_02562_));
 sky130_fd_sc_hd__a21o_1 _10828_ (.A1(_02559_),
    .A2(_02561_),
    .B1(_02344_),
    .X(_02563_));
 sky130_fd_sc_hd__nand3_1 _10829_ (.A(_02561_),
    .B(_02344_),
    .C(_02559_),
    .Y(_02564_));
 sky130_fd_sc_hd__o211ai_2 _10830_ (.A1(_02333_),
    .A2(_02329_),
    .B1(_02078_),
    .C1(_02336_),
    .Y(_02565_));
 sky130_fd_sc_hd__and4_1 _10831_ (.A(_02334_),
    .B(_02563_),
    .C(_02564_),
    .D(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__a22oi_1 _10832_ (.A1(_02563_),
    .A2(_02564_),
    .B1(_02565_),
    .B2(_02334_),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_1 _10833_ (.A(_02566_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__or3_1 _10834_ (.A(_00834_),
    .B(_02568_),
    .C(_02343_),
    .X(_02569_));
 sky130_fd_sc_hd__o21ai_1 _10835_ (.A1(_00834_),
    .A2(_02343_),
    .B1(_02568_),
    .Y(_02570_));
 sky130_fd_sc_hd__and2_1 _10836_ (.A(_02569_),
    .B(_02570_),
    .X(net82));
 sky130_fd_sc_hd__a31o_1 _10837_ (.A1(_02085_),
    .A2(_02339_),
    .A3(_02568_),
    .B1(_00834_),
    .X(_02572_));
 sky130_fd_sc_hd__o21ai_2 _10838_ (.A1(_02421_),
    .A2(_02553_),
    .B1(_02556_),
    .Y(_02573_));
 sky130_fd_sc_hd__a31o_1 _10839_ (.A1(_02377_),
    .A2(_02394_),
    .A3(_02395_),
    .B1(_02378_),
    .X(_02574_));
 sky130_fd_sc_hd__or4_2 _10840_ (.A(_03479_),
    .B(_03522_),
    .C(_01399_),
    .D(_01404_),
    .X(_02575_));
 sky130_fd_sc_hd__and3_1 _10841_ (.A(_04726_),
    .B(net145),
    .C(_01220_),
    .X(_02576_));
 sky130_fd_sc_hd__o2bb2ai_1 _10842_ (.A1_N(_02382_),
    .A2_N(_02383_),
    .B1(net158),
    .B2(_01058_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_1 _10843_ (.A(_02577_),
    .B(_02576_),
    .Y(_02578_));
 sky130_fd_sc_hd__a21oi_2 _10844_ (.A1(_02383_),
    .A2(_02382_),
    .B1(_02576_),
    .Y(_02579_));
 sky130_fd_sc_hd__o31a_1 _10845_ (.A1(net158),
    .A2(_01399_),
    .A3(_01404_),
    .B1(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__o2bb2ai_2 _10846_ (.A1_N(_02576_),
    .A2_N(_02577_),
    .B1(_02579_),
    .B2(_02575_),
    .Y(_02582_));
 sky130_fd_sc_hd__o32a_1 _10847_ (.A1(net158),
    .A2(net136),
    .A3(_02578_),
    .B1(_02580_),
    .B2(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__o22ai_1 _10848_ (.A1(_02575_),
    .A2(_02578_),
    .B1(_02580_),
    .B2(_02582_),
    .Y(_02584_));
 sky130_fd_sc_hd__o21ai_1 _10849_ (.A1(_02367_),
    .A2(_02369_),
    .B1(_02368_),
    .Y(_02585_));
 sky130_fd_sc_hd__o21ai_1 _10850_ (.A1(_02017_),
    .A2(_02252_),
    .B1(_02393_),
    .Y(_02586_));
 sky130_fd_sc_hd__nand2_1 _10851_ (.A(_02392_),
    .B(_02255_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand3_2 _10852_ (.A(_02585_),
    .B(_02586_),
    .C(_02392_),
    .Y(_02588_));
 sky130_fd_sc_hd__o2111ai_4 _10853_ (.A1(_02369_),
    .A2(_02367_),
    .B1(_02368_),
    .C1(_02393_),
    .D1(_02587_),
    .Y(_02589_));
 sky130_fd_sc_hd__a21o_1 _10854_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02584_),
    .X(_02590_));
 sky130_fd_sc_hd__nand3_1 _10855_ (.A(_02584_),
    .B(_02588_),
    .C(_02589_),
    .Y(_02591_));
 sky130_fd_sc_hd__a21o_1 _10856_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02583_),
    .X(_02593_));
 sky130_fd_sc_hd__nand3_1 _10857_ (.A(_02589_),
    .B(_02583_),
    .C(_02588_),
    .Y(_02594_));
 sky130_fd_sc_hd__and3_1 _10858_ (.A(_02590_),
    .B(_02591_),
    .C(_02574_),
    .X(_02595_));
 sky130_fd_sc_hd__nand3_1 _10859_ (.A(_02590_),
    .B(_02591_),
    .C(_02574_),
    .Y(_02596_));
 sky130_fd_sc_hd__nand3b_2 _10860_ (.A_N(_02574_),
    .B(_02593_),
    .C(_02594_),
    .Y(_02597_));
 sky130_fd_sc_hd__and3_1 _10861_ (.A(_01631_),
    .B(_02050_),
    .C(_02052_),
    .X(_02598_));
 sky130_fd_sc_hd__and4_1 _10862_ (.A(_01590_),
    .B(_01820_),
    .C(_01821_),
    .D(_02899_),
    .X(_02599_));
 sky130_fd_sc_hd__o32a_1 _10863_ (.A1(net159),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(_02122_),
    .X(_02600_));
 sky130_fd_sc_hd__o22ai_2 _10864_ (.A1(net159),
    .A2(_01589_),
    .B1(_01822_),
    .B2(_02122_),
    .Y(_02601_));
 sky130_fd_sc_hd__o32a_1 _10865_ (.A1(_01620_),
    .A2(_02049_),
    .A3(_02051_),
    .B1(_02599_),
    .B2(_02600_),
    .X(_02602_));
 sky130_fd_sc_hd__o311a_1 _10866_ (.A1(_02910_),
    .A2(_01589_),
    .A3(_01822_),
    .B1(_02598_),
    .C1(_02601_),
    .X(_02604_));
 sky130_fd_sc_hd__nor2_1 _10867_ (.A(_02602_),
    .B(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__a21bo_1 _10868_ (.A1(_02596_),
    .A2(_02597_),
    .B1_N(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__o211ai_1 _10869_ (.A1(_02602_),
    .A2(_02604_),
    .B1(_02596_),
    .C1(_02597_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand3b_1 _10870_ (.A_N(_02403_),
    .B(_02606_),
    .C(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__a221o_1 _10871_ (.A1(_02371_),
    .A2(_02401_),
    .B1(_02606_),
    .B2(_02607_),
    .C1(_02399_),
    .X(_02609_));
 sky130_fd_sc_hd__nand2_1 _10872_ (.A(_02608_),
    .B(_02609_),
    .Y(_02610_));
 sky130_fd_sc_hd__o211ai_2 _10873_ (.A1(_02366_),
    .A2(_02405_),
    .B1(_02308_),
    .C1(_02311_),
    .Y(_02611_));
 sky130_fd_sc_hd__o211ai_2 _10874_ (.A1(_02365_),
    .A2(_02404_),
    .B1(_02608_),
    .C1(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__o211ai_2 _10875_ (.A1(_02365_),
    .A2(_02404_),
    .B1(_02610_),
    .C1(_02611_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21o_1 _10876_ (.A1(_02408_),
    .A2(_02611_),
    .B1(_02610_),
    .X(_02615_));
 sky130_fd_sc_hd__a32o_1 _10877_ (.A1(_06341_),
    .A2(_00899_),
    .A3(_00902_),
    .B1(_00569_),
    .B2(net151),
    .X(_02616_));
 sky130_fd_sc_hd__or4_1 _10878_ (.A(_06331_),
    .B(net152),
    .C(_00570_),
    .D(_00903_),
    .X(_02617_));
 sky130_fd_sc_hd__a22oi_1 _10879_ (.A1(_05436_),
    .A2(net141),
    .B1(_02616_),
    .B2(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__and4_1 _10880_ (.A(_05436_),
    .B(net141),
    .C(_02616_),
    .D(_02617_),
    .X(_02619_));
 sky130_fd_sc_hd__nor2_1 _10881_ (.A(_02618_),
    .B(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__xor2_2 _10882_ (.A(_02362_),
    .B(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__and3_1 _10883_ (.A(_02613_),
    .B(_02615_),
    .C(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__a21oi_1 _10884_ (.A1(_02613_),
    .A2(_02615_),
    .B1(_02621_),
    .Y(_02623_));
 sky130_fd_sc_hd__a21o_1 _10885_ (.A1(_02613_),
    .A2(_02615_),
    .B1(_02621_),
    .X(_02624_));
 sky130_fd_sc_hd__nor2_2 _10886_ (.A(net17),
    .B(net18),
    .Y(_02626_));
 sky130_fd_sc_hd__nand4b_4 _10887_ (.A_N(net18),
    .B(_01581_),
    .C(_02045_),
    .D(_02347_),
    .Y(_02627_));
 sky130_fd_sc_hd__a21oi_4 _10888_ (.A1(_02627_),
    .A2(net174),
    .B1(net19),
    .Y(_02628_));
 sky130_fd_sc_hd__a21o_4 _10889_ (.A1(_02627_),
    .A2(net174),
    .B1(net19),
    .X(_02629_));
 sky130_fd_sc_hd__o311a_4 _10890_ (.A1(_02348_),
    .A2(net18),
    .A3(_02048_),
    .B1(net19),
    .C1(net174),
    .X(_02630_));
 sky130_fd_sc_hd__o211ai_4 _10891_ (.A1(net18),
    .A2(_02349_),
    .B1(net19),
    .C1(net174),
    .Y(_02631_));
 sky130_fd_sc_hd__nand2_8 _10892_ (.A(_02629_),
    .B(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__nor2_8 _10893_ (.A(_02628_),
    .B(_02630_),
    .Y(_02633_));
 sky130_fd_sc_hd__o32a_1 _10894_ (.A1(_00900_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_01292_),
    .B2(_02241_),
    .X(_02634_));
 sky130_fd_sc_hd__and4_1 _10895_ (.A(_02240_),
    .B(_02356_),
    .C(_00911_),
    .D(_01303_),
    .X(_02635_));
 sky130_fd_sc_hd__or4_1 _10896_ (.A(_00900_),
    .B(_01292_),
    .C(_02241_),
    .D(_02355_),
    .X(_02637_));
 sky130_fd_sc_hd__o32a_1 _10897_ (.A1(_00310_),
    .A2(_02628_),
    .A3(_02630_),
    .B1(_02634_),
    .B2(_02635_),
    .X(_02638_));
 sky130_fd_sc_hd__or4_2 _10898_ (.A(_00310_),
    .B(_02632_),
    .C(_02634_),
    .D(_02635_),
    .X(_02639_));
 sky130_fd_sc_hd__nand2b_2 _10899_ (.A_N(_02638_),
    .B(_02639_),
    .Y(_02640_));
 sky130_fd_sc_hd__xnor2_4 _10900_ (.A(_02357_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__o21bai_2 _10901_ (.A1(_02622_),
    .A2(_02623_),
    .B1_N(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__nand3b_2 _10902_ (.A_N(_02622_),
    .B(_02624_),
    .C(_02641_),
    .Y(_02643_));
 sky130_fd_sc_hd__o21bai_2 _10903_ (.A1(_02359_),
    .A2(_02412_),
    .B1_N(_02411_),
    .Y(_02644_));
 sky130_fd_sc_hd__and3_1 _10904_ (.A(_02642_),
    .B(_02643_),
    .C(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__a21oi_2 _10905_ (.A1(_02642_),
    .A2(_02643_),
    .B1(_02644_),
    .Y(_02646_));
 sky130_fd_sc_hd__or2_1 _10906_ (.A(_02645_),
    .B(_02646_),
    .X(_02648_));
 sky130_fd_sc_hd__and4_1 _10907_ (.A(_02346_),
    .B(_02414_),
    .C(_02415_),
    .D(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__nor2_1 _10908_ (.A(_02416_),
    .B(_02648_),
    .Y(_02650_));
 sky130_fd_sc_hd__o21ai_1 _10909_ (.A1(_02534_),
    .A2(_02542_),
    .B1(_02535_),
    .Y(_02651_));
 sky130_fd_sc_hd__o21ba_1 _10910_ (.A1(_02519_),
    .A2(_02530_),
    .B1_N(_02518_),
    .X(_02652_));
 sky130_fd_sc_hd__o31a_1 _10911_ (.A1(net153),
    .A2(_00532_),
    .A3(_02539_),
    .B1(_02538_),
    .X(_02653_));
 sky130_fd_sc_hd__o21a_1 _10912_ (.A1(_02191_),
    .A2(_02526_),
    .B1(_02527_),
    .X(_02654_));
 sky130_fd_sc_hd__xnor2_1 _10913_ (.A(_02653_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__or4_1 _10914_ (.A(_00067_),
    .B(_00069_),
    .C(_00270_),
    .D(_00272_),
    .X(_02656_));
 sky130_fd_sc_hd__o32a_1 _10915_ (.A1(_07441_),
    .A2(_00270_),
    .A3(_00272_),
    .B1(_02521_),
    .B2(_02522_),
    .X(_02657_));
 sky130_fd_sc_hd__or3_1 _10916_ (.A(_07539_),
    .B(_00428_),
    .C(_02657_),
    .X(_02659_));
 sky130_fd_sc_hd__o32a_1 _10917_ (.A1(_00071_),
    .A2(net143),
    .A3(_02522_),
    .B1(_00428_),
    .B2(_07539_),
    .X(_02660_));
 sky130_fd_sc_hd__or4_1 _10918_ (.A(_00071_),
    .B(_00270_),
    .C(_00272_),
    .D(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__o32a_1 _10919_ (.A1(_07539_),
    .A2(_00428_),
    .A3(_02657_),
    .B1(_02656_),
    .B2(_02660_),
    .X(_02662_));
 sky130_fd_sc_hd__o21ai_1 _10920_ (.A1(_00071_),
    .A2(_00274_),
    .B1(_02660_),
    .Y(_02663_));
 sky130_fd_sc_hd__o2bb2a_1 _10921_ (.A1_N(_02663_),
    .A2_N(_02662_),
    .B1(_02659_),
    .B2(_02656_),
    .X(_02664_));
 sky130_fd_sc_hd__xnor2_1 _10922_ (.A(_02655_),
    .B(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _10923_ (.A(_02665_),
    .B(_02652_),
    .Y(_02666_));
 sky130_fd_sc_hd__or2_1 _10924_ (.A(_02652_),
    .B(_02665_),
    .X(_02667_));
 sky130_fd_sc_hd__o32a_1 _10925_ (.A1(_00005_),
    .A2(_00007_),
    .A3(_00366_),
    .B1(_00192_),
    .B2(net143),
    .X(_02668_));
 sky130_fd_sc_hd__or4_1 _10926_ (.A(_00145_),
    .B(_00147_),
    .C(_00361_),
    .D(_00363_),
    .X(_02670_));
 sky130_fd_sc_hd__and4_1 _10927_ (.A(_00010_),
    .B(_00150_),
    .C(_00193_),
    .D(_00367_),
    .X(_02671_));
 sky130_fd_sc_hd__o22ai_1 _10928_ (.A1(_07512_),
    .A2(_00532_),
    .B1(_02668_),
    .B2(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__or4_1 _10929_ (.A(_07512_),
    .B(_00532_),
    .C(_02668_),
    .D(_02671_),
    .X(_02673_));
 sky130_fd_sc_hd__nand2_1 _10930_ (.A(_02672_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__nand3_1 _10931_ (.A(_02666_),
    .B(_02667_),
    .C(_02674_),
    .Y(_02675_));
 sky130_fd_sc_hd__a21o_1 _10932_ (.A1(_02666_),
    .A2(_02667_),
    .B1(_02674_),
    .X(_02676_));
 sky130_fd_sc_hd__and3_1 _10933_ (.A(_02676_),
    .B(_02651_),
    .C(_02675_),
    .X(_02677_));
 sky130_fd_sc_hd__a21o_1 _10934_ (.A1(_02675_),
    .A2(_02676_),
    .B1(_02651_),
    .X(_02678_));
 sky130_fd_sc_hd__nand2b_2 _10935_ (.A_N(_02677_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__a22o_1 _10936_ (.A1(_02213_),
    .A2(_02543_),
    .B1(_02219_),
    .B2(_02217_),
    .X(_02681_));
 sky130_fd_sc_hd__o22ai_4 _10937_ (.A1(_02213_),
    .A2(_02543_),
    .B1(_02216_),
    .B2(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__xor2_4 _10938_ (.A(_02679_),
    .B(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__a31o_1 _10939_ (.A1(_02222_),
    .A2(_02509_),
    .A3(_02548_),
    .B1(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__o2111a_1 _10940_ (.A1(_02546_),
    .A2(_02547_),
    .B1(_02222_),
    .C1(_02683_),
    .D1(_02509_),
    .X(_02685_));
 sky130_fd_sc_hd__o2111ai_4 _10941_ (.A1(_02546_),
    .A2(_02547_),
    .B1(_02222_),
    .C1(_02683_),
    .D1(_02509_),
    .Y(_02686_));
 sky130_fd_sc_hd__a32o_1 _10942_ (.A1(_02437_),
    .A2(_02496_),
    .A3(_02498_),
    .B1(_02500_),
    .B2(_02425_),
    .X(_02687_));
 sky130_fd_sc_hd__nor2_4 _10943_ (.A(net49),
    .B(net50),
    .Y(_02688_));
 sky130_fd_sc_hd__or2_1 _10944_ (.A(net49),
    .B(net50),
    .X(_02689_));
 sky130_fd_sc_hd__nand4b_4 _10945_ (.A_N(_01535_),
    .B(_02087_),
    .C(_02688_),
    .D(_00682_),
    .Y(_02690_));
 sky130_fd_sc_hd__a21oi_4 _10946_ (.A1(_02690_),
    .A2(net173),
    .B1(net51),
    .Y(_02692_));
 sky130_fd_sc_hd__a21o_4 _10947_ (.A1(_02690_),
    .A2(net173),
    .B1(net51),
    .X(_02693_));
 sky130_fd_sc_hd__o311a_4 _10948_ (.A1(net49),
    .A2(net50),
    .A3(_02091_),
    .B1(net51),
    .C1(net173),
    .X(_02694_));
 sky130_fd_sc_hd__a211o_4 _10949_ (.A1(_02090_),
    .A2(_02688_),
    .B1(_00299_),
    .C1(_00736_),
    .X(_02695_));
 sky130_fd_sc_hd__nand2_8 _10950_ (.A(_02693_),
    .B(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__nor2_8 _10951_ (.A(_02692_),
    .B(_02694_),
    .Y(_02697_));
 sky130_fd_sc_hd__a31o_1 _10952_ (.A1(_02690_),
    .A2(net51),
    .A3(net173),
    .B1(_00987_),
    .X(_02698_));
 sky130_fd_sc_hd__nor2_1 _10953_ (.A(_02692_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__and3_1 _10954_ (.A(net1),
    .B(_02432_),
    .C(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__a32o_1 _10955_ (.A1(_00998_),
    .A2(_02427_),
    .A3(_02428_),
    .B1(_02697_),
    .B2(net1),
    .X(_02701_));
 sky130_fd_sc_hd__o41ai_2 _10956_ (.A1(_00288_),
    .A2(_02433_),
    .A3(_02692_),
    .A4(_02698_),
    .B1(_02701_),
    .Y(_02703_));
 sky130_fd_sc_hd__o31a_1 _10957_ (.A1(net166),
    .A2(_02092_),
    .A3(_02094_),
    .B1(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__or3_1 _10958_ (.A(net166),
    .B(_02096_),
    .C(_02703_),
    .X(_02705_));
 sky130_fd_sc_hd__nand2b_2 _10959_ (.A_N(_02704_),
    .B(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__xor2_4 _10960_ (.A(_02435_),
    .B(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__o211ai_4 _10961_ (.A1(_02168_),
    .A2(_02169_),
    .B1(_02489_),
    .C1(_02493_),
    .Y(_02708_));
 sky130_fd_sc_hd__o211ai_4 _10962_ (.A1(_02490_),
    .A2(_02487_),
    .B1(_02170_),
    .C1(_02492_),
    .Y(_02709_));
 sky130_fd_sc_hd__a32oi_4 _10963_ (.A1(_02138_),
    .A2(_02438_),
    .A3(_02148_),
    .B1(_02464_),
    .B2(_02463_),
    .Y(_02710_));
 sky130_fd_sc_hd__a31oi_2 _10964_ (.A1(_02439_),
    .A2(_02466_),
    .A3(_02468_),
    .B1(_02441_),
    .Y(_02711_));
 sky130_fd_sc_hd__o32a_1 _10965_ (.A1(_03906_),
    .A2(_01188_),
    .A3(_02117_),
    .B1(_04244_),
    .B2(_01037_),
    .X(_02712_));
 sky130_fd_sc_hd__nor2_1 _10966_ (.A(_02475_),
    .B(_02712_),
    .Y(_02714_));
 sky130_fd_sc_hd__o21ai_1 _10967_ (.A1(_01872_),
    .A2(_02117_),
    .B1(_02459_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand3_4 _10968_ (.A(_02461_),
    .B(_02714_),
    .C(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__o221ai_4 _10969_ (.A1(_02475_),
    .A2(_02712_),
    .B1(_02120_),
    .B2(_02460_),
    .C1(_02459_),
    .Y(_02717_));
 sky130_fd_sc_hd__or3_2 _10970_ (.A(_01958_),
    .B(_01658_),
    .C(_01660_),
    .X(_02718_));
 sky130_fd_sc_hd__a21oi_1 _10971_ (.A1(_02127_),
    .A2(_02449_),
    .B1(_02448_),
    .Y(_02719_));
 sky130_fd_sc_hd__and3_1 _10972_ (.A(_01499_),
    .B(net135),
    .C(_01880_),
    .X(_02720_));
 sky130_fd_sc_hd__o21ai_4 _10973_ (.A1(_02124_),
    .A2(_02719_),
    .B1(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__a21oi_1 _10974_ (.A1(_02450_),
    .A2(_02447_),
    .B1(_02720_),
    .Y(_02722_));
 sky130_fd_sc_hd__a31o_1 _10975_ (.A1(_01969_),
    .A2(_01544_),
    .A3(_02450_),
    .B1(_02720_),
    .X(_02723_));
 sky130_fd_sc_hd__a22oi_2 _10976_ (.A1(_01969_),
    .A2(_01664_),
    .B1(_02721_),
    .B2(_02723_),
    .Y(_02725_));
 sky130_fd_sc_hd__and4_1 _10977_ (.A(_01969_),
    .B(_01664_),
    .C(_02721_),
    .D(_02723_),
    .X(_02726_));
 sky130_fd_sc_hd__a21oi_2 _10978_ (.A1(_02721_),
    .A2(_02723_),
    .B1(_02718_),
    .Y(_02727_));
 sky130_fd_sc_hd__o311a_1 _10979_ (.A1(_01958_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_02721_),
    .C1(_02723_),
    .X(_02728_));
 sky130_fd_sc_hd__o211ai_2 _10980_ (.A1(_02725_),
    .A2(_02726_),
    .B1(_02716_),
    .C1(_02717_),
    .Y(_02729_));
 sky130_fd_sc_hd__o2bb2ai_2 _10981_ (.A1_N(_02716_),
    .A2_N(_02717_),
    .B1(_02727_),
    .B2(_02728_),
    .Y(_02730_));
 sky130_fd_sc_hd__o2bb2ai_1 _10982_ (.A1_N(_02716_),
    .A2_N(_02717_),
    .B1(_02725_),
    .B2(_02726_),
    .Y(_02731_));
 sky130_fd_sc_hd__o211ai_2 _10983_ (.A1(_02727_),
    .A2(_02728_),
    .B1(_02716_),
    .C1(_02717_),
    .Y(_02732_));
 sky130_fd_sc_hd__nand2_1 _10984_ (.A(_02729_),
    .B(_02730_),
    .Y(_02733_));
 sky130_fd_sc_hd__nand3_2 _10985_ (.A(_02711_),
    .B(_02731_),
    .C(_02732_),
    .Y(_02734_));
 sky130_fd_sc_hd__and3_1 _10986_ (.A(_03917_),
    .B(_01539_),
    .C(_01541_),
    .X(_02736_));
 sky130_fd_sc_hd__and3_1 _10987_ (.A(_02736_),
    .B(_01273_),
    .C(_02647_),
    .X(_02737_));
 sky130_fd_sc_hd__o32a_2 _10988_ (.A1(_02636_),
    .A2(_01538_),
    .A3(_01540_),
    .B1(_03906_),
    .B2(_01272_),
    .X(_02738_));
 sky130_fd_sc_hd__o32a_1 _10989_ (.A1(_04244_),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_02737_),
    .B2(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__nor4_2 _10990_ (.A(_04244_),
    .B(_01188_),
    .C(_02737_),
    .D(_02738_),
    .Y(_02740_));
 sky130_fd_sc_hd__nor2_1 _10991_ (.A(_02739_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__inv_2 _10992_ (.A(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__o211a_1 _10993_ (.A1(_02441_),
    .A2(_02710_),
    .B1(_02729_),
    .C1(_02730_),
    .X(_02743_));
 sky130_fd_sc_hd__o211ai_2 _10994_ (.A1(_02441_),
    .A2(_02710_),
    .B1(_02729_),
    .C1(_02730_),
    .Y(_02744_));
 sky130_fd_sc_hd__a31o_1 _10995_ (.A1(_02711_),
    .A2(_02731_),
    .A3(_02732_),
    .B1(_02741_),
    .X(_02745_));
 sky130_fd_sc_hd__o31a_2 _10996_ (.A1(_02739_),
    .A2(_02740_),
    .A3(_02743_),
    .B1(_02734_),
    .X(_02747_));
 sky130_fd_sc_hd__inv_2 _10997_ (.A(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__o211a_1 _10998_ (.A1(_02739_),
    .A2(_02740_),
    .B1(_02744_),
    .C1(_02734_),
    .X(_02749_));
 sky130_fd_sc_hd__a21oi_1 _10999_ (.A1(_02734_),
    .A2(_02744_),
    .B1(_02742_),
    .Y(_02750_));
 sky130_fd_sc_hd__a21o_1 _11000_ (.A1(_02734_),
    .A2(_02744_),
    .B1(_02742_),
    .X(_02751_));
 sky130_fd_sc_hd__o21a_2 _11001_ (.A1(_02743_),
    .A2(_02745_),
    .B1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o211ai_4 _11002_ (.A1(_02745_),
    .A2(_02743_),
    .B1(_02482_),
    .C1(_02751_),
    .Y(_02753_));
 sky130_fd_sc_hd__o21bai_2 _11003_ (.A1(_02749_),
    .A2(_02750_),
    .B1_N(_02482_),
    .Y(_02754_));
 sky130_fd_sc_hd__and2_1 _11004_ (.A(_02753_),
    .B(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__nand2_1 _11005_ (.A(_02753_),
    .B(_02754_),
    .Y(_02756_));
 sky130_fd_sc_hd__o211ai_1 _11006_ (.A1(_02490_),
    .A2(_02487_),
    .B1(_02756_),
    .C1(_02708_),
    .Y(_02758_));
 sky130_fd_sc_hd__o211ai_1 _11007_ (.A1(_02162_),
    .A2(_02488_),
    .B1(_02755_),
    .C1(_02709_),
    .Y(_02759_));
 sky130_fd_sc_hd__o211ai_2 _11008_ (.A1(_02162_),
    .A2(_02488_),
    .B1(_02709_),
    .C1(_02756_),
    .Y(_02760_));
 sky130_fd_sc_hd__o211ai_2 _11009_ (.A1(_02487_),
    .A2(_02490_),
    .B1(_02708_),
    .C1(_02755_),
    .Y(_02761_));
 sky130_fd_sc_hd__nand3_1 _11010_ (.A(_02760_),
    .B(_02761_),
    .C(_02707_),
    .Y(_02762_));
 sky130_fd_sc_hd__nand3b_2 _11011_ (.A_N(_02707_),
    .B(_02758_),
    .C(_02759_),
    .Y(_02763_));
 sky130_fd_sc_hd__and4_1 _11012_ (.A(_05316_),
    .B(_00743_),
    .C(_01038_),
    .D(_07200_),
    .X(_02764_));
 sky130_fd_sc_hd__o32a_1 _11013_ (.A1(_05327_),
    .A2(_01033_),
    .A3(_01035_),
    .B1(_07189_),
    .B2(_00744_),
    .X(_02765_));
 sky130_fd_sc_hd__o32a_1 _11014_ (.A1(_07441_),
    .A2(_00576_),
    .A3(_00578_),
    .B1(_02764_),
    .B2(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__or4_1 _11015_ (.A(_07441_),
    .B(_00580_),
    .C(_02764_),
    .D(_02765_),
    .X(_02767_));
 sky130_fd_sc_hd__nand2b_1 _11016_ (.A_N(_02766_),
    .B(_02767_),
    .Y(_02769_));
 sky130_fd_sc_hd__o31a_1 _11017_ (.A1(_07189_),
    .A2(_00744_),
    .A3(_02086_),
    .B1(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__nor4_1 _11018_ (.A(_07189_),
    .B(_00744_),
    .C(_02086_),
    .D(_02769_),
    .Y(_02771_));
 sky130_fd_sc_hd__nor2_1 _11019_ (.A(_02770_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__nand3_1 _11020_ (.A(_02762_),
    .B(_02763_),
    .C(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__o2bb2ai_1 _11021_ (.A1_N(_02762_),
    .A2_N(_02763_),
    .B1(_02770_),
    .B2(_02771_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand3_2 _11022_ (.A(_02687_),
    .B(_02773_),
    .C(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__a21oi_1 _11023_ (.A1(_02773_),
    .A2(_02774_),
    .B1(_02687_),
    .Y(_02776_));
 sky130_fd_sc_hd__a21o_1 _11024_ (.A1(_02773_),
    .A2(_02774_),
    .B1(_02687_),
    .X(_02777_));
 sky130_fd_sc_hd__a21oi_1 _11025_ (.A1(_02775_),
    .A2(_02777_),
    .B1(_02505_),
    .Y(_02778_));
 sky130_fd_sc_hd__and3_1 _11026_ (.A(_02505_),
    .B(_02775_),
    .C(_02777_),
    .X(_02780_));
 sky130_fd_sc_hd__or2_4 _11027_ (.A(_02778_),
    .B(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__a21oi_2 _11028_ (.A1(_02684_),
    .A2(_02686_),
    .B1(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__and3_1 _11029_ (.A(_02684_),
    .B(_02686_),
    .C(_02781_),
    .X(_02783_));
 sky130_fd_sc_hd__a311o_1 _11030_ (.A1(_02684_),
    .A2(_02686_),
    .A3(_02781_),
    .B1(_02650_),
    .C1(_02649_),
    .X(_02784_));
 sky130_fd_sc_hd__o22ai_2 _11031_ (.A1(_02649_),
    .A2(_02650_),
    .B1(_02782_),
    .B2(_02783_),
    .Y(_02785_));
 sky130_fd_sc_hd__o21a_1 _11032_ (.A1(_02782_),
    .A2(_02784_),
    .B1(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__o211ai_2 _11033_ (.A1(_02782_),
    .A2(_02784_),
    .B1(_02573_),
    .C1(_02785_),
    .Y(_02787_));
 sky130_fd_sc_hd__a211o_1 _11034_ (.A1(_02420_),
    .A2(_02554_),
    .B1(_02555_),
    .C1(_02786_),
    .X(_02788_));
 sky130_fd_sc_hd__o211ai_2 _11035_ (.A1(_02330_),
    .A2(_02332_),
    .B1(_02564_),
    .C1(_02565_),
    .Y(_02789_));
 sky130_fd_sc_hd__o2111ai_1 _11036_ (.A1(_02344_),
    .A2(_02562_),
    .B1(_02787_),
    .C1(_02788_),
    .D1(_02789_),
    .Y(_02791_));
 sky130_fd_sc_hd__a22o_1 _11037_ (.A1(_02787_),
    .A2(_02788_),
    .B1(_02789_),
    .B2(_02563_),
    .X(_02792_));
 sky130_fd_sc_hd__nand2_1 _11038_ (.A(_02791_),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__xor2_1 _11039_ (.A(_02572_),
    .B(_02793_),
    .X(net83));
 sky130_fd_sc_hd__nand4_1 _11040_ (.A(_02793_),
    .B(_02339_),
    .C(_02085_),
    .D(_02568_),
    .Y(_02794_));
 sky130_fd_sc_hd__and2b_1 _11041_ (.A_N(_02782_),
    .B(_02784_),
    .X(_02795_));
 sky130_fd_sc_hd__a31o_1 _11042_ (.A1(_02613_),
    .A2(_02615_),
    .A3(_02621_),
    .B1(_02641_),
    .X(_02796_));
 sky130_fd_sc_hd__a32o_1 _11043_ (.A1(net151),
    .A2(_00899_),
    .A3(_00902_),
    .B1(_00569_),
    .B2(_07513_),
    .X(_02797_));
 sky130_fd_sc_hd__or4_1 _11044_ (.A(_07508_),
    .B(_07510_),
    .C(_00898_),
    .D(_00901_),
    .X(_02798_));
 sky130_fd_sc_hd__nand4_2 _11045_ (.A(_00569_),
    .B(_00904_),
    .C(net151),
    .D(_07513_),
    .Y(_02799_));
 sky130_fd_sc_hd__a32o_1 _11046_ (.A1(_06341_),
    .A2(_01055_),
    .A3(_01057_),
    .B1(_02797_),
    .B2(_02799_),
    .X(_02801_));
 sky130_fd_sc_hd__and4_1 _11047_ (.A(_06341_),
    .B(net141),
    .C(_02797_),
    .D(_02799_),
    .X(_02802_));
 sky130_fd_sc_hd__nand4_1 _11048_ (.A(_06341_),
    .B(net141),
    .C(_02797_),
    .D(_02799_),
    .Y(_02803_));
 sky130_fd_sc_hd__a32o_1 _11049_ (.A1(_05392_),
    .A2(_05414_),
    .A3(_01222_),
    .B1(_02801_),
    .B2(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__o2111ai_1 _11050_ (.A1(_05359_),
    .A2(_05370_),
    .B1(_01222_),
    .C1(_02801_),
    .D1(_02803_),
    .Y(_02805_));
 sky130_fd_sc_hd__nand2_1 _11051_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__o41a_1 _11052_ (.A1(_06331_),
    .A2(net152),
    .A3(_00570_),
    .A4(_00903_),
    .B1(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__or2_1 _11053_ (.A(_02617_),
    .B(_02806_),
    .X(_02808_));
 sky130_fd_sc_hd__nand2b_1 _11054_ (.A_N(_02807_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__o21ba_1 _11055_ (.A1(_02362_),
    .A2(_02618_),
    .B1_N(_02619_),
    .X(_02810_));
 sky130_fd_sc_hd__xor2_1 _11056_ (.A(_02809_),
    .B(_02810_),
    .X(_02812_));
 sky130_fd_sc_hd__inv_2 _11057_ (.A(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__a32o_1 _11058_ (.A1(_02899_),
    .A2(_01590_),
    .A3(_01823_),
    .B1(_02601_),
    .B2(_02598_),
    .X(_02814_));
 sky130_fd_sc_hd__a21oi_1 _11059_ (.A1(_02598_),
    .A2(_02601_),
    .B1(_02599_),
    .Y(_02815_));
 sky130_fd_sc_hd__o211ai_4 _11060_ (.A1(_02579_),
    .A2(_02575_),
    .B1(_02578_),
    .C1(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__nand2_1 _11061_ (.A(_02582_),
    .B(_02814_),
    .Y(_02817_));
 sky130_fd_sc_hd__nand4_1 _11062_ (.A(_01405_),
    .B(_01590_),
    .C(net156),
    .D(_04726_),
    .Y(_02818_));
 sky130_fd_sc_hd__o32a_1 _11063_ (.A1(net158),
    .A2(_01584_),
    .A3(_01586_),
    .B1(net155),
    .B2(net136),
    .X(_02819_));
 sky130_fd_sc_hd__a32o_1 _11064_ (.A1(net156),
    .A2(_01585_),
    .A3(_01588_),
    .B1(_01405_),
    .B2(_04726_),
    .X(_02820_));
 sky130_fd_sc_hd__a22oi_2 _11065_ (.A1(_02866_),
    .A2(_01823_),
    .B1(_02818_),
    .B2(_02820_),
    .Y(_02821_));
 sky130_fd_sc_hd__and4_1 _11066_ (.A(_02866_),
    .B(_01823_),
    .C(_02818_),
    .D(_02820_),
    .X(_02823_));
 sky130_fd_sc_hd__nor2_1 _11067_ (.A(_02821_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__a2bb2o_1 _11068_ (.A1_N(_02821_),
    .A2_N(_02823_),
    .B1(_02582_),
    .B2(_02814_),
    .X(_02825_));
 sky130_fd_sc_hd__nand3_2 _11069_ (.A(_02824_),
    .B(_02817_),
    .C(_02816_),
    .Y(_02826_));
 sky130_fd_sc_hd__o2bb2ai_2 _11070_ (.A1_N(_02816_),
    .A2_N(_02817_),
    .B1(_02821_),
    .B2(_02823_),
    .Y(_02827_));
 sky130_fd_sc_hd__nand2_1 _11071_ (.A(_02583_),
    .B(_02588_),
    .Y(_02828_));
 sky130_fd_sc_hd__a22oi_4 _11072_ (.A1(_02826_),
    .A2(_02827_),
    .B1(_02828_),
    .B2(_02589_),
    .Y(_02829_));
 sky130_fd_sc_hd__and4_1 _11073_ (.A(_02589_),
    .B(_02826_),
    .C(_02827_),
    .D(_02828_),
    .X(_02830_));
 sky130_fd_sc_hd__nand4_1 _11074_ (.A(_02589_),
    .B(_02826_),
    .C(_02827_),
    .D(_02828_),
    .Y(_02831_));
 sky130_fd_sc_hd__a2111o_1 _11075_ (.A1(_02046_),
    .A2(_02068_),
    .B1(_02053_),
    .C1(_02829_),
    .D1(_02830_),
    .X(_02832_));
 sky130_fd_sc_hd__o22ai_4 _11076_ (.A1(_02122_),
    .A2(_02053_),
    .B1(_02829_),
    .B2(_02830_),
    .Y(_02834_));
 sky130_fd_sc_hd__and2_1 _11077_ (.A(_02832_),
    .B(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__o21a_1 _11078_ (.A1(_02602_),
    .A2(_02604_),
    .B1(_02596_),
    .X(_02836_));
 sky130_fd_sc_hd__o21a_1 _11079_ (.A1(_02595_),
    .A2(_02605_),
    .B1(_02597_),
    .X(_02837_));
 sky130_fd_sc_hd__a21oi_2 _11080_ (.A1(_02832_),
    .A2(_02834_),
    .B1(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21o_1 _11081_ (.A1(_02832_),
    .A2(_02834_),
    .B1(_02837_),
    .X(_02839_));
 sky130_fd_sc_hd__nand2_1 _11082_ (.A(_02835_),
    .B(_02597_),
    .Y(_02840_));
 sky130_fd_sc_hd__and3_1 _11083_ (.A(_02832_),
    .B(_02834_),
    .C(_02837_),
    .X(_02841_));
 sky130_fd_sc_hd__nand2_1 _11084_ (.A(_02609_),
    .B(_02612_),
    .Y(_02842_));
 sky130_fd_sc_hd__o21ai_1 _11085_ (.A1(_02838_),
    .A2(_02841_),
    .B1(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__o211ai_4 _11086_ (.A1(_02836_),
    .A2(_02840_),
    .B1(_02609_),
    .C1(_02612_),
    .Y(_02845_));
 sky130_fd_sc_hd__o21ai_1 _11087_ (.A1(_02838_),
    .A2(_02845_),
    .B1(_02843_),
    .Y(_02846_));
 sky130_fd_sc_hd__o211a_1 _11088_ (.A1(_02845_),
    .A2(_02838_),
    .B1(_02813_),
    .C1(_02843_),
    .X(_02847_));
 sky130_fd_sc_hd__o211ai_2 _11089_ (.A1(_02845_),
    .A2(_02838_),
    .B1(_02813_),
    .C1(_02843_),
    .Y(_02848_));
 sky130_fd_sc_hd__nand2_1 _11090_ (.A(_02812_),
    .B(_02846_),
    .Y(_02849_));
 sky130_fd_sc_hd__nor2_1 _11091_ (.A(net18),
    .B(net19),
    .Y(_02850_));
 sky130_fd_sc_hd__nand4_4 _11092_ (.A(_01581_),
    .B(_02045_),
    .C(_02347_),
    .D(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__o211ai_4 _11093_ (.A1(net19),
    .A2(_02627_),
    .B1(_00747_),
    .C1(net25),
    .Y(_02852_));
 sky130_fd_sc_hd__a21o_4 _11094_ (.A1(_02851_),
    .A2(net25),
    .B1(_00747_),
    .X(_02853_));
 sky130_fd_sc_hd__o211ai_4 _11095_ (.A1(net19),
    .A2(_02627_),
    .B1(net20),
    .C1(net25),
    .Y(_02854_));
 sky130_fd_sc_hd__a21o_4 _11096_ (.A1(_02851_),
    .A2(net25),
    .B1(net20),
    .X(_02856_));
 sky130_fd_sc_hd__nand2_8 _11097_ (.A(_02854_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__nand2_8 _11098_ (.A(_02852_),
    .B(_02853_),
    .Y(_02858_));
 sky130_fd_sc_hd__a32o_1 _11099_ (.A1(_01631_),
    .A2(net139),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_01303_),
    .X(_02859_));
 sky130_fd_sc_hd__nand4_2 _11100_ (.A(_02240_),
    .B(_02356_),
    .C(_01303_),
    .D(_01631_),
    .Y(_02860_));
 sky130_fd_sc_hd__a32o_1 _11101_ (.A1(_00911_),
    .A2(_02629_),
    .A3(_02631_),
    .B1(_02859_),
    .B2(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__and4_1 _11102_ (.A(_00911_),
    .B(_02633_),
    .C(_02859_),
    .D(_02860_),
    .X(_02862_));
 sky130_fd_sc_hd__o2111ai_1 _11103_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_02633_),
    .C1(_02859_),
    .D1(_02860_),
    .Y(_02863_));
 sky130_fd_sc_hd__o2bb2a_1 _11104_ (.A1_N(_02861_),
    .A2_N(_02863_),
    .B1(_00310_),
    .B2(_02857_),
    .X(_02864_));
 sky130_fd_sc_hd__and4_1 _11105_ (.A(_02861_),
    .B(net33),
    .C(_02858_),
    .D(_02863_),
    .X(_02865_));
 sky130_fd_sc_hd__or3_1 _11106_ (.A(_02865_),
    .B(_02637_),
    .C(_02864_),
    .X(_02867_));
 sky130_fd_sc_hd__o21ai_1 _11107_ (.A1(_02864_),
    .A2(_02865_),
    .B1(_02637_),
    .Y(_02868_));
 sky130_fd_sc_hd__o21ai_2 _11108_ (.A1(_02357_),
    .A2(_02638_),
    .B1(_02639_),
    .Y(_02869_));
 sky130_fd_sc_hd__a21o_1 _11109_ (.A1(_02867_),
    .A2(_02868_),
    .B1(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__nand3_1 _11110_ (.A(_02867_),
    .B(_02868_),
    .C(_02869_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_1 _11111_ (.A(_02870_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__nand3_2 _11112_ (.A(_02848_),
    .B(_02849_),
    .C(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__a21o_1 _11113_ (.A1(_02848_),
    .A2(_02849_),
    .B1(_02872_),
    .X(_02874_));
 sky130_fd_sc_hd__a22o_1 _11114_ (.A1(_02624_),
    .A2(_02796_),
    .B1(_02873_),
    .B2(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__o2111ai_4 _11115_ (.A1(_02641_),
    .A2(_02622_),
    .B1(_02624_),
    .C1(_02873_),
    .D1(_02874_),
    .Y(_02876_));
 sky130_fd_sc_hd__a31oi_2 _11116_ (.A1(_02642_),
    .A2(_02643_),
    .A3(_02644_),
    .B1(_02417_),
    .Y(_02878_));
 sky130_fd_sc_hd__a211oi_2 _11117_ (.A1(_02875_),
    .A2(_02876_),
    .B1(_02878_),
    .C1(_02646_),
    .Y(_02879_));
 sky130_fd_sc_hd__o21ai_1 _11118_ (.A1(_02646_),
    .A2(_02878_),
    .B1(_02876_),
    .Y(_02880_));
 sky130_fd_sc_hd__o211a_1 _11119_ (.A1(_02646_),
    .A2(_02878_),
    .B1(_02876_),
    .C1(_02875_),
    .X(_02881_));
 sky130_fd_sc_hd__or2_1 _11120_ (.A(_02879_),
    .B(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__a21o_1 _11121_ (.A1(_02665_),
    .A2(_02652_),
    .B1(_02674_),
    .X(_02883_));
 sky130_fd_sc_hd__a21o_1 _11122_ (.A1(_02653_),
    .A2(_02654_),
    .B1(_02664_),
    .X(_02884_));
 sky130_fd_sc_hd__o21a_1 _11123_ (.A1(_02653_),
    .A2(_02654_),
    .B1(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__a32o_1 _11124_ (.A1(_00072_),
    .A2(_00425_),
    .A3(_00427_),
    .B1(_00193_),
    .B2(_00275_),
    .X(_02886_));
 sky130_fd_sc_hd__and4_1 _11125_ (.A(_00072_),
    .B(_00193_),
    .C(_00275_),
    .D(_00429_),
    .X(_02887_));
 sky130_fd_sc_hd__o31a_1 _11126_ (.A1(_00192_),
    .A2(_00428_),
    .A3(_02656_),
    .B1(_02886_),
    .X(_02889_));
 sky130_fd_sc_hd__xnor2_1 _11127_ (.A(_02670_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__o32a_1 _11128_ (.A1(_00009_),
    .A2(_00192_),
    .A3(_02670_),
    .B1(_00532_),
    .B2(_07512_),
    .X(_02891_));
 sky130_fd_sc_hd__a211oi_1 _11129_ (.A1(_02659_),
    .A2(_02661_),
    .B1(_02668_),
    .C1(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__o211a_1 _11130_ (.A1(_02668_),
    .A2(_02891_),
    .B1(_02659_),
    .C1(_02661_),
    .X(_02893_));
 sky130_fd_sc_hd__o21ba_1 _11131_ (.A1(_02890_),
    .A2(_02892_),
    .B1_N(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__o21ai_1 _11132_ (.A1(_02892_),
    .A2(_02893_),
    .B1(_02890_),
    .Y(_02895_));
 sky130_fd_sc_hd__or3_1 _11133_ (.A(_02890_),
    .B(_02892_),
    .C(_02893_),
    .X(_02896_));
 sky130_fd_sc_hd__and2_1 _11134_ (.A(_02895_),
    .B(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__xnor2_1 _11135_ (.A(_02885_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__o21ai_1 _11136_ (.A1(_00009_),
    .A2(_00532_),
    .B1(_02898_),
    .Y(_02900_));
 sky130_fd_sc_hd__or4_1 _11137_ (.A(_00005_),
    .B(_00007_),
    .C(_00532_),
    .D(_02898_),
    .X(_02901_));
 sky130_fd_sc_hd__nand2_1 _11138_ (.A(_02900_),
    .B(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__and3_1 _11139_ (.A(_02667_),
    .B(_02883_),
    .C(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__a21o_1 _11140_ (.A1(_02667_),
    .A2(_02883_),
    .B1(_02902_),
    .X(_02904_));
 sky130_fd_sc_hd__nand2b_1 _11141_ (.A_N(_02903_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__inv_2 _11142_ (.A(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__o21a_1 _11143_ (.A1(_02677_),
    .A2(_02682_),
    .B1(_02678_),
    .X(_02907_));
 sky130_fd_sc_hd__nor2_2 _11144_ (.A(_02906_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__o211a_2 _11145_ (.A1(_02677_),
    .A2(_02682_),
    .B1(_02906_),
    .C1(_02678_),
    .X(_02909_));
 sky130_fd_sc_hd__or2_1 _11146_ (.A(_02908_),
    .B(_02909_),
    .X(_02911_));
 sky130_fd_sc_hd__a41o_1 _11147_ (.A1(_02509_),
    .A2(_02683_),
    .A3(_02548_),
    .A4(_02222_),
    .B1(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__o2111ai_4 _11148_ (.A1(_02908_),
    .A2(_02909_),
    .B1(_02548_),
    .C1(_02683_),
    .D1(_02511_),
    .Y(_02913_));
 sky130_fd_sc_hd__nand2_1 _11149_ (.A(_02912_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__a32oi_4 _11150_ (.A1(_02707_),
    .A2(_02760_),
    .A3(_02761_),
    .B1(_02763_),
    .B2(_02772_),
    .Y(_02915_));
 sky130_fd_sc_hd__and3_1 _11151_ (.A(net164),
    .B(_02427_),
    .C(_02428_),
    .X(_02916_));
 sky130_fd_sc_hd__nor2_2 _11152_ (.A(net50),
    .B(net51),
    .Y(_02917_));
 sky130_fd_sc_hd__nor3_1 _11153_ (.A(_02689_),
    .B(net51),
    .C(_02091_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand4b_2 _11154_ (.A_N(_01656_),
    .B(_02087_),
    .C(_02688_),
    .D(_00736_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21oi_4 _11155_ (.A1(_02919_),
    .A2(net173),
    .B1(net52),
    .Y(_02920_));
 sky130_fd_sc_hd__a21o_4 _11156_ (.A1(_02919_),
    .A2(net173),
    .B1(net52),
    .X(_02922_));
 sky130_fd_sc_hd__o311a_4 _11157_ (.A1(_02689_),
    .A2(net51),
    .A3(_02091_),
    .B1(net52),
    .C1(net173),
    .X(_02923_));
 sky130_fd_sc_hd__o211ai_4 _11158_ (.A1(net51),
    .A2(_02690_),
    .B1(net52),
    .C1(net173),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_8 _11159_ (.A(_02922_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__nor2_8 _11160_ (.A(_02920_),
    .B(_02923_),
    .Y(_02926_));
 sky130_fd_sc_hd__and3_1 _11161_ (.A(_02926_),
    .B(_02699_),
    .C(net1),
    .X(_02927_));
 sky130_fd_sc_hd__nand4_1 _11162_ (.A(net1),
    .B(_02699_),
    .C(_02922_),
    .D(_02924_),
    .Y(_02928_));
 sky130_fd_sc_hd__a31o_1 _11163_ (.A1(net1),
    .A2(_02922_),
    .A3(_02924_),
    .B1(_02699_),
    .X(_02929_));
 sky130_fd_sc_hd__and3_1 _11164_ (.A(_02928_),
    .B(_02929_),
    .C(_02916_),
    .X(_02930_));
 sky130_fd_sc_hd__nand4_1 _11165_ (.A(net164),
    .B(_02928_),
    .C(_02929_),
    .D(_02432_),
    .Y(_02931_));
 sky130_fd_sc_hd__a32o_1 _11166_ (.A1(net164),
    .A2(_02427_),
    .A3(_02428_),
    .B1(_02928_),
    .B2(_02929_),
    .X(_02933_));
 sky130_fd_sc_hd__a32o_1 _11167_ (.A1(_01499_),
    .A2(_02093_),
    .A3(_02095_),
    .B1(_02931_),
    .B2(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__o2111ai_1 _11168_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_02097_),
    .C1(_02931_),
    .D1(_02933_),
    .Y(_02935_));
 sky130_fd_sc_hd__a31o_1 _11169_ (.A1(_01499_),
    .A2(_02093_),
    .A3(_02095_),
    .B1(_02930_),
    .X(_02936_));
 sky130_fd_sc_hd__a21oi_1 _11170_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02700_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand3_1 _11171_ (.A(_02934_),
    .B(_02935_),
    .C(_02700_),
    .Y(_02938_));
 sky130_fd_sc_hd__nand2b_1 _11172_ (.A_N(_02937_),
    .B(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__o41a_1 _11173_ (.A1(_00987_),
    .A2(_02098_),
    .A3(_02433_),
    .A4(_02704_),
    .B1(_02705_),
    .X(_02940_));
 sky130_fd_sc_hd__o211a_1 _11174_ (.A1(_02704_),
    .A2(_02435_),
    .B1(_02938_),
    .C1(_02705_),
    .X(_02941_));
 sky130_fd_sc_hd__xnor2_2 _11175_ (.A(_02939_),
    .B(_02940_),
    .Y(_02942_));
 sky130_fd_sc_hd__o211ai_4 _11176_ (.A1(_02490_),
    .A2(_02487_),
    .B1(_02753_),
    .C1(_02708_),
    .Y(_02944_));
 sky130_fd_sc_hd__o221ai_4 _11177_ (.A1(_02162_),
    .A2(_02488_),
    .B1(_02752_),
    .B2(_02482_),
    .C1(_02709_),
    .Y(_02945_));
 sky130_fd_sc_hd__a22o_1 _11178_ (.A1(_04201_),
    .A2(_04212_),
    .B1(_01266_),
    .B2(_01267_),
    .X(_02946_));
 sky130_fd_sc_hd__o21ai_1 _11179_ (.A1(_02727_),
    .A2(_02728_),
    .B1(_02717_),
    .Y(_02947_));
 sky130_fd_sc_hd__o21ai_1 _11180_ (.A1(_02718_),
    .A2(_02722_),
    .B1(_02721_),
    .Y(_02948_));
 sky130_fd_sc_hd__a2111oi_1 _11181_ (.A1(_04201_),
    .A2(_04212_),
    .B1(_01184_),
    .C1(_01186_),
    .D1(_02738_),
    .Y(_02949_));
 sky130_fd_sc_hd__o32a_1 _11182_ (.A1(_03906_),
    .A2(_01542_),
    .A3(_02117_),
    .B1(_04244_),
    .B2(_01188_),
    .X(_02950_));
 sky130_fd_sc_hd__o21ai_1 _11183_ (.A1(_02737_),
    .A2(_02949_),
    .B1(_02948_),
    .Y(_02951_));
 sky130_fd_sc_hd__o221a_1 _11184_ (.A1(_02738_),
    .A2(_02950_),
    .B1(_02718_),
    .B2(_02722_),
    .C1(_02721_),
    .X(_02952_));
 sky130_fd_sc_hd__o221ai_2 _11185_ (.A1(_02738_),
    .A2(_02950_),
    .B1(_02718_),
    .B2(_02722_),
    .C1(_02721_),
    .Y(_02953_));
 sky130_fd_sc_hd__or3_1 _11186_ (.A(_02636_),
    .B(_01658_),
    .C(_01660_),
    .X(_02955_));
 sky130_fd_sc_hd__o32a_1 _11187_ (.A1(_02636_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_01882_),
    .B2(_01958_),
    .X(_02956_));
 sky130_fd_sc_hd__a32o_1 _11188_ (.A1(_01969_),
    .A2(net135),
    .A3(_01880_),
    .B1(_02647_),
    .B2(_01664_),
    .X(_02957_));
 sky130_fd_sc_hd__and4_1 _11189_ (.A(_01969_),
    .B(_02647_),
    .C(_01664_),
    .D(_01883_),
    .X(_02958_));
 sky130_fd_sc_hd__o32a_1 _11190_ (.A1(_03906_),
    .A2(_01538_),
    .A3(_01540_),
    .B1(_02956_),
    .B2(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__o311a_1 _11191_ (.A1(_02636_),
    .A2(_01882_),
    .A3(_02718_),
    .B1(_02736_),
    .C1(_02957_),
    .X(_02960_));
 sky130_fd_sc_hd__o211ai_2 _11192_ (.A1(_02959_),
    .A2(_02960_),
    .B1(_02951_),
    .C1(_02953_),
    .Y(_02961_));
 sky130_fd_sc_hd__a211o_1 _11193_ (.A1(_02951_),
    .A2(_02953_),
    .B1(_02959_),
    .C1(_02960_),
    .X(_02962_));
 sky130_fd_sc_hd__and4_1 _11194_ (.A(_02716_),
    .B(_02947_),
    .C(_02961_),
    .D(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__nand4_1 _11195_ (.A(_02716_),
    .B(_02947_),
    .C(_02961_),
    .D(_02962_),
    .Y(_02964_));
 sky130_fd_sc_hd__a22o_1 _11196_ (.A1(_02716_),
    .A2(_02947_),
    .B1(_02961_),
    .B2(_02962_),
    .X(_02966_));
 sky130_fd_sc_hd__a21oi_1 _11197_ (.A1(_02964_),
    .A2(_02966_),
    .B1(_02946_),
    .Y(_02967_));
 sky130_fd_sc_hd__and3_1 _11198_ (.A(_02946_),
    .B(_02964_),
    .C(_02966_),
    .X(_02968_));
 sky130_fd_sc_hd__nor2_2 _11199_ (.A(_02967_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__inv_2 _11200_ (.A(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__o221a_1 _11201_ (.A1(_02711_),
    .A2(_02733_),
    .B1(_02967_),
    .B2(_02968_),
    .C1(_02745_),
    .X(_02971_));
 sky130_fd_sc_hd__o311a_1 _11202_ (.A1(_02739_),
    .A2(_02740_),
    .A3(_02743_),
    .B1(_02969_),
    .C1(_02734_),
    .X(_02972_));
 sky130_fd_sc_hd__or3_1 _11203_ (.A(_02748_),
    .B(_02967_),
    .C(_02968_),
    .X(_02973_));
 sky130_fd_sc_hd__nor2_1 _11204_ (.A(_02971_),
    .B(_02972_),
    .Y(_02974_));
 sky130_fd_sc_hd__o211ai_2 _11205_ (.A1(_02971_),
    .A2(_02972_),
    .B1(_02753_),
    .C1(_02945_),
    .Y(_02975_));
 sky130_fd_sc_hd__o211ai_2 _11206_ (.A1(_02482_),
    .A2(_02752_),
    .B1(_02944_),
    .C1(_02974_),
    .Y(_02977_));
 sky130_fd_sc_hd__o221ai_2 _11207_ (.A1(_02482_),
    .A2(_02752_),
    .B1(_02971_),
    .B2(_02972_),
    .C1(_02944_),
    .Y(_02978_));
 sky130_fd_sc_hd__nand3_1 _11208_ (.A(_02974_),
    .B(_02945_),
    .C(_02753_),
    .Y(_02979_));
 sky130_fd_sc_hd__nand3_1 _11209_ (.A(_02977_),
    .B(_02942_),
    .C(_02975_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand3b_2 _11210_ (.A_N(_02942_),
    .B(_02978_),
    .C(_02979_),
    .Y(_02981_));
 sky130_fd_sc_hd__a32o_1 _11211_ (.A1(_05316_),
    .A2(_01185_),
    .A3(_01187_),
    .B1(_07200_),
    .B2(_01038_),
    .X(_02982_));
 sky130_fd_sc_hd__or4_2 _11212_ (.A(_05327_),
    .B(_07189_),
    .C(_01037_),
    .D(_01188_),
    .X(_02983_));
 sky130_fd_sc_hd__nand4_1 _11213_ (.A(_02983_),
    .B(_00743_),
    .C(_07440_),
    .D(_02982_),
    .Y(_02984_));
 sky130_fd_sc_hd__a32o_1 _11214_ (.A1(net162),
    .A2(_00743_),
    .A3(_07437_),
    .B1(_02983_),
    .B2(_02982_),
    .X(_02985_));
 sky130_fd_sc_hd__a32o_1 _11215_ (.A1(_07540_),
    .A2(_00577_),
    .A3(_00579_),
    .B1(_02984_),
    .B2(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__nand4_1 _11216_ (.A(_07540_),
    .B(_00581_),
    .C(_02984_),
    .D(_02985_),
    .Y(_02988_));
 sky130_fd_sc_hd__nand2_1 _11217_ (.A(_02986_),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__o41a_1 _11218_ (.A1(_05327_),
    .A2(_07189_),
    .A3(_00744_),
    .A4(_01037_),
    .B1(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__and3_1 _11219_ (.A(_02986_),
    .B(_02988_),
    .C(_02764_),
    .X(_02991_));
 sky130_fd_sc_hd__a31o_1 _11220_ (.A1(_02764_),
    .A2(_02986_),
    .A3(_02988_),
    .B1(_02990_),
    .X(_02992_));
 sky130_fd_sc_hd__o41a_2 _11221_ (.A1(_07189_),
    .A2(_00744_),
    .A3(_02086_),
    .A4(_02766_),
    .B1(_02767_),
    .X(_02993_));
 sky130_fd_sc_hd__xnor2_4 _11222_ (.A(_02992_),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__nand3_1 _11223_ (.A(_02980_),
    .B(_02981_),
    .C(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__a21o_1 _11224_ (.A1(_02980_),
    .A2(_02981_),
    .B1(_02994_),
    .X(_02996_));
 sky130_fd_sc_hd__nand3_2 _11225_ (.A(_02996_),
    .B(_02915_),
    .C(_02995_),
    .Y(_02997_));
 sky130_fd_sc_hd__a21oi_1 _11226_ (.A1(_02995_),
    .A2(_02996_),
    .B1(_02915_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21o_1 _11227_ (.A1(_02995_),
    .A2(_02996_),
    .B1(_02915_),
    .X(_03000_));
 sky130_fd_sc_hd__nand2_4 _11228_ (.A(_02997_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__o21ai_4 _11229_ (.A1(_02505_),
    .A2(_02776_),
    .B1(_02775_),
    .Y(_03002_));
 sky130_fd_sc_hd__xnor2_4 _11230_ (.A(_03001_),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__xor2_4 _11231_ (.A(_03001_),
    .B(_03002_),
    .X(_03004_));
 sky130_fd_sc_hd__a21oi_1 _11232_ (.A1(_02912_),
    .A2(_02913_),
    .B1(_03003_),
    .Y(_03005_));
 sky130_fd_sc_hd__a21o_1 _11233_ (.A1(_02912_),
    .A2(_02913_),
    .B1(_03003_),
    .X(_03006_));
 sky130_fd_sc_hd__nand3_1 _11234_ (.A(_02912_),
    .B(_02913_),
    .C(_03003_),
    .Y(_03007_));
 sky130_fd_sc_hd__o22a_1 _11235_ (.A1(_02879_),
    .A2(_02881_),
    .B1(_02914_),
    .B2(_03004_),
    .X(_03008_));
 sky130_fd_sc_hd__o221a_1 _11236_ (.A1(_02879_),
    .A2(_02881_),
    .B1(_02914_),
    .B2(_03004_),
    .C1(_03006_),
    .X(_03010_));
 sky130_fd_sc_hd__a21oi_1 _11237_ (.A1(_03006_),
    .A2(_03007_),
    .B1(_02882_),
    .Y(_03011_));
 sky130_fd_sc_hd__a21o_1 _11238_ (.A1(_03006_),
    .A2(_03008_),
    .B1(_03011_),
    .X(_03012_));
 sky130_fd_sc_hd__nor2_1 _11239_ (.A(_02795_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__o21ai_1 _11240_ (.A1(_03010_),
    .A2(_03011_),
    .B1(_02795_),
    .Y(_03014_));
 sky130_fd_sc_hd__and2b_1 _11241_ (.A_N(_03013_),
    .B(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__o211ai_2 _11242_ (.A1(_02344_),
    .A2(_02562_),
    .B1(_02787_),
    .C1(_02789_),
    .Y(_03016_));
 sky130_fd_sc_hd__o21a_1 _11243_ (.A1(_02573_),
    .A2(_02786_),
    .B1(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__xnor2_1 _11244_ (.A(_03015_),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__xor2_1 _11245_ (.A(_03015_),
    .B(_03017_),
    .X(_03019_));
 sky130_fd_sc_hd__a21o_1 _11246_ (.A1(_00845_),
    .A2(_02794_),
    .B1(_03018_),
    .X(_03021_));
 sky130_fd_sc_hd__a311o_1 _11247_ (.A1(_02343_),
    .A2(_02568_),
    .A3(_02793_),
    .B1(_00834_),
    .C1(_03019_),
    .X(_03022_));
 sky130_fd_sc_hd__and2_1 _11248_ (.A(_03021_),
    .B(_03022_),
    .X(net84));
 sky130_fd_sc_hd__and4_1 _11249_ (.A(_02568_),
    .B(_02793_),
    .C(_03019_),
    .D(_02343_),
    .X(_03023_));
 sky130_fd_sc_hd__o22a_1 _11250_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_02794_),
    .B2(_03018_),
    .X(_03024_));
 sky130_fd_sc_hd__a31o_1 _11251_ (.A1(_00150_),
    .A2(_00367_),
    .A3(_02886_),
    .B1(_02887_),
    .X(_03025_));
 sky130_fd_sc_hd__or3_1 _11252_ (.A(_00145_),
    .B(_00147_),
    .C(_00532_),
    .X(_03026_));
 sky130_fd_sc_hd__o32a_1 _11253_ (.A1(_00270_),
    .A2(_00272_),
    .A3(_00366_),
    .B1(_00428_),
    .B2(_00192_),
    .X(_03027_));
 sky130_fd_sc_hd__and4_1 _11254_ (.A(_00193_),
    .B(_00275_),
    .C(_00367_),
    .D(_00429_),
    .X(_03028_));
 sky130_fd_sc_hd__or2_1 _11255_ (.A(_03027_),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__xnor2_1 _11256_ (.A(_03026_),
    .B(_03029_),
    .Y(_03031_));
 sky130_fd_sc_hd__nand2b_1 _11257_ (.A_N(_03031_),
    .B(_02894_),
    .Y(_03032_));
 sky130_fd_sc_hd__nand2b_1 _11258_ (.A_N(_02894_),
    .B(_03031_),
    .Y(_03033_));
 sky130_fd_sc_hd__and3_1 _11259_ (.A(_03025_),
    .B(_03032_),
    .C(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__a21oi_1 _11260_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_03025_),
    .Y(_03035_));
 sky130_fd_sc_hd__or2_1 _11261_ (.A(_03034_),
    .B(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__o32a_1 _11262_ (.A1(_00005_),
    .A2(_00007_),
    .A3(_00532_),
    .B1(_02885_),
    .B2(_02897_),
    .X(_03037_));
 sky130_fd_sc_hd__a21o_1 _11263_ (.A1(_02885_),
    .A2(_02897_),
    .B1(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__nand2_1 _11264_ (.A(_03036_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__nor2_1 _11265_ (.A(_03038_),
    .B(_03036_),
    .Y(_03040_));
 sky130_fd_sc_hd__a211o_1 _11266_ (.A1(_02885_),
    .A2(_02897_),
    .B1(_03036_),
    .C1(_03037_),
    .X(_03042_));
 sky130_fd_sc_hd__nand2_2 _11267_ (.A(_03039_),
    .B(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__o21ai_4 _11268_ (.A1(_02903_),
    .A2(_02907_),
    .B1(_02904_),
    .Y(_03044_));
 sky130_fd_sc_hd__xnor2_4 _11269_ (.A(_03043_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__o211ai_2 _11270_ (.A1(_02908_),
    .A2(_02909_),
    .B1(_03045_),
    .C1(_02685_),
    .Y(_03046_));
 sky130_fd_sc_hd__a41o_1 _11271_ (.A1(_02511_),
    .A2(_02548_),
    .A3(_02683_),
    .A4(_02911_),
    .B1(_03045_),
    .X(_03047_));
 sky130_fd_sc_hd__a32oi_4 _11272_ (.A1(_02942_),
    .A2(_02975_),
    .A3(_02977_),
    .B1(_02981_),
    .B2(_02994_),
    .Y(_03048_));
 sky130_fd_sc_hd__nand4_2 _11273_ (.A(_07200_),
    .B(_01189_),
    .C(_01273_),
    .D(_05316_),
    .Y(_03049_));
 sky130_fd_sc_hd__a31oi_2 _11274_ (.A1(_01265_),
    .A2(net45),
    .A3(net173),
    .B1(_05327_),
    .Y(_03050_));
 sky130_fd_sc_hd__a32o_1 _11275_ (.A1(_07200_),
    .A2(_01185_),
    .A3(_01187_),
    .B1(_01269_),
    .B2(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__a211o_1 _11276_ (.A1(_01269_),
    .A2(_03050_),
    .B1(_07189_),
    .C1(_01188_),
    .X(_03053_));
 sky130_fd_sc_hd__o211ai_2 _11277_ (.A1(_07189_),
    .A2(_01188_),
    .B1(_01273_),
    .C1(_05316_),
    .Y(_03054_));
 sky130_fd_sc_hd__o311a_1 _11278_ (.A1(_07441_),
    .A2(_01033_),
    .A3(_01035_),
    .B1(_03053_),
    .C1(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__o211ai_2 _11279_ (.A1(_01037_),
    .A2(_07441_),
    .B1(_03054_),
    .C1(_03053_),
    .Y(_03056_));
 sky130_fd_sc_hd__nand4_2 _11280_ (.A(_01038_),
    .B(_03049_),
    .C(_03051_),
    .D(_07440_),
    .Y(_03057_));
 sky130_fd_sc_hd__a211o_1 _11281_ (.A1(_03056_),
    .A2(_03057_),
    .B1(net149),
    .C1(_00744_),
    .X(_03058_));
 sky130_fd_sc_hd__o211ai_2 _11282_ (.A1(_00744_),
    .A2(net149),
    .B1(_03057_),
    .C1(_03056_),
    .Y(_03059_));
 sky130_fd_sc_hd__and3_1 _11283_ (.A(_02983_),
    .B(_03058_),
    .C(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__nand3_1 _11284_ (.A(_02983_),
    .B(_03058_),
    .C(_03059_),
    .Y(_03061_));
 sky130_fd_sc_hd__a21o_1 _11285_ (.A1(_03058_),
    .A2(_03059_),
    .B1(_02983_),
    .X(_03062_));
 sky130_fd_sc_hd__a22oi_1 _11286_ (.A1(_00072_),
    .A2(_00581_),
    .B1(_03061_),
    .B2(_03062_),
    .Y(_03064_));
 sky130_fd_sc_hd__nand4_1 _11287_ (.A(_00072_),
    .B(_00581_),
    .C(_03061_),
    .D(_03062_),
    .Y(_03065_));
 sky130_fd_sc_hd__and2b_1 _11288_ (.A_N(_03064_),
    .B(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__and3_1 _11289_ (.A(_07540_),
    .B(_00581_),
    .C(_02985_),
    .X(_03067_));
 sky130_fd_sc_hd__a41o_1 _11290_ (.A1(_07440_),
    .A2(_00743_),
    .A3(_02982_),
    .A4(_02983_),
    .B1(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__nand2_1 _11291_ (.A(_03066_),
    .B(_03068_),
    .Y(_03069_));
 sky130_fd_sc_hd__nor2_1 _11292_ (.A(_03066_),
    .B(_03068_),
    .Y(_03070_));
 sky130_fd_sc_hd__or2_1 _11293_ (.A(_03066_),
    .B(_03068_),
    .X(_03071_));
 sky130_fd_sc_hd__o21ba_1 _11294_ (.A1(_02993_),
    .A2(_02990_),
    .B1_N(_02991_),
    .X(_03072_));
 sky130_fd_sc_hd__a21oi_1 _11295_ (.A1(_03069_),
    .A2(_03071_),
    .B1(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__nand3_1 _11296_ (.A(_03069_),
    .B(_03071_),
    .C(_03072_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2b_2 _11297_ (.A_N(_03073_),
    .B(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__and3_1 _11298_ (.A(_01499_),
    .B(_02427_),
    .C(_02428_),
    .X(_03077_));
 sky130_fd_sc_hd__nor2_4 _11299_ (.A(net51),
    .B(net52),
    .Y(_03078_));
 sky130_fd_sc_hd__nand4b_4 _11300_ (.A_N(_01656_),
    .B(_02087_),
    .C(_02688_),
    .D(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_1 _11301_ (.A(_03079_),
    .B(net173),
    .Y(_03080_));
 sky130_fd_sc_hd__a311oi_4 _11302_ (.A1(_02090_),
    .A2(_02688_),
    .A3(_03078_),
    .B1(_00758_),
    .C1(_00299_),
    .Y(_03081_));
 sky130_fd_sc_hd__a311o_4 _11303_ (.A1(_02090_),
    .A2(_02688_),
    .A3(_03078_),
    .B1(_00758_),
    .C1(_00299_),
    .X(_03082_));
 sky130_fd_sc_hd__a21oi_4 _11304_ (.A1(_03079_),
    .A2(net173),
    .B1(net53),
    .Y(_03083_));
 sky130_fd_sc_hd__a21o_4 _11305_ (.A1(_03079_),
    .A2(net173),
    .B1(net53),
    .X(_03084_));
 sky130_fd_sc_hd__nand2_8 _11306_ (.A(_03082_),
    .B(_03084_),
    .Y(_03086_));
 sky130_fd_sc_hd__nor2_8 _11307_ (.A(net132),
    .B(net130),
    .Y(_03087_));
 sky130_fd_sc_hd__a21oi_1 _11308_ (.A1(_00758_),
    .A2(_03080_),
    .B1(_00288_),
    .Y(_03088_));
 sky130_fd_sc_hd__o32ai_4 _11309_ (.A1(_00288_),
    .A2(_03081_),
    .A3(_03083_),
    .B1(_00987_),
    .B2(_02925_),
    .Y(_03089_));
 sky130_fd_sc_hd__o2111ai_4 _11310_ (.A1(_00921_),
    .A2(_00943_),
    .B1(net1),
    .C1(_03082_),
    .D1(_03084_),
    .Y(_03090_));
 sky130_fd_sc_hd__and4_1 _11311_ (.A(_02926_),
    .B(_03088_),
    .C(_03082_),
    .D(_00998_),
    .X(_03091_));
 sky130_fd_sc_hd__nand4_1 _11312_ (.A(_02926_),
    .B(_03088_),
    .C(_03082_),
    .D(_00998_),
    .Y(_03092_));
 sky130_fd_sc_hd__o2111a_1 _11313_ (.A1(_03090_),
    .A2(_02925_),
    .B1(_02697_),
    .C1(net164),
    .D1(_03089_),
    .X(_03093_));
 sky130_fd_sc_hd__o2111ai_4 _11314_ (.A1(_03090_),
    .A2(_02925_),
    .B1(_02697_),
    .C1(net164),
    .D1(_03089_),
    .Y(_03094_));
 sky130_fd_sc_hd__a22oi_1 _11315_ (.A1(net164),
    .A2(_02697_),
    .B1(_03089_),
    .B2(_03092_),
    .Y(_03095_));
 sky130_fd_sc_hd__a22o_1 _11316_ (.A1(net164),
    .A2(_02697_),
    .B1(_03089_),
    .B2(_03092_),
    .X(_03097_));
 sky130_fd_sc_hd__o22ai_2 _11317_ (.A1(_02433_),
    .A2(_01488_),
    .B1(_03095_),
    .B2(_03093_),
    .Y(_03098_));
 sky130_fd_sc_hd__o2111ai_4 _11318_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_02432_),
    .C1(_03094_),
    .D1(_03097_),
    .Y(_03099_));
 sky130_fd_sc_hd__a21oi_1 _11319_ (.A1(_03098_),
    .A2(_03099_),
    .B1(_02927_),
    .Y(_03100_));
 sky130_fd_sc_hd__a32o_1 _11320_ (.A1(net1),
    .A2(_02926_),
    .A3(_02699_),
    .B1(_03099_),
    .B2(_03098_),
    .X(_03101_));
 sky130_fd_sc_hd__nand3_2 _11321_ (.A(_03098_),
    .B(_03099_),
    .C(_02927_),
    .Y(_03102_));
 sky130_fd_sc_hd__a22o_1 _11322_ (.A1(_01969_),
    .A2(_02097_),
    .B1(_03101_),
    .B2(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__o2111ai_4 _11323_ (.A1(_01892_),
    .A2(_01914_),
    .B1(_02097_),
    .C1(_03101_),
    .D1(_03102_),
    .Y(_03104_));
 sky130_fd_sc_hd__a31o_1 _11324_ (.A1(_01499_),
    .A2(_02097_),
    .A3(_02933_),
    .B1(_02930_),
    .X(_03105_));
 sky130_fd_sc_hd__nand4_1 _11325_ (.A(_02933_),
    .B(_02936_),
    .C(_03103_),
    .D(_03104_),
    .Y(_03106_));
 sky130_fd_sc_hd__a21oi_1 _11326_ (.A1(_03103_),
    .A2(_03104_),
    .B1(_03105_),
    .Y(_03108_));
 sky130_fd_sc_hd__a22o_1 _11327_ (.A1(_02933_),
    .A2(_02936_),
    .B1(_03103_),
    .B2(_03104_),
    .X(_03109_));
 sky130_fd_sc_hd__a21oi_1 _11328_ (.A1(_02938_),
    .A2(_02940_),
    .B1(_02937_),
    .Y(_03110_));
 sky130_fd_sc_hd__a2bb2o_1 _11329_ (.A1_N(_02937_),
    .A2_N(_02941_),
    .B1(_03106_),
    .B2(_03109_),
    .X(_03111_));
 sky130_fd_sc_hd__or4bb_1 _11330_ (.A(_02937_),
    .B(_02941_),
    .C_N(_03106_),
    .D_N(_03109_),
    .X(_03112_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(_03111_),
    .B(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__nand2_1 _11332_ (.A(_03111_),
    .B(_03112_),
    .Y(_03114_));
 sky130_fd_sc_hd__and3_1 _11333_ (.A(_04255_),
    .B(_01539_),
    .C(_01541_),
    .X(_03115_));
 sky130_fd_sc_hd__o32a_1 _11334_ (.A1(_03906_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_01882_),
    .B2(_02636_),
    .X(_03116_));
 sky130_fd_sc_hd__and4_1 _11335_ (.A(_02647_),
    .B(_03917_),
    .C(_01664_),
    .D(_01883_),
    .X(_03117_));
 sky130_fd_sc_hd__nor2_1 _11336_ (.A(_03116_),
    .B(_03117_),
    .Y(_03119_));
 sky130_fd_sc_hd__xnor2_2 _11337_ (.A(_03115_),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__o31a_2 _11338_ (.A1(_02952_),
    .A2(_02959_),
    .A3(_02960_),
    .B1(_02951_),
    .X(_03121_));
 sky130_fd_sc_hd__xnor2_1 _11339_ (.A(_03120_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__a31o_1 _11340_ (.A1(_03917_),
    .A2(_01544_),
    .A3(_02957_),
    .B1(_02958_),
    .X(_03123_));
 sky130_fd_sc_hd__and2b_1 _11341_ (.A_N(_03123_),
    .B(_03122_),
    .X(_03124_));
 sky130_fd_sc_hd__and2b_1 _11342_ (.A_N(_03122_),
    .B(_03123_),
    .X(_03125_));
 sky130_fd_sc_hd__nor2_1 _11343_ (.A(_03124_),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__o21ai_2 _11344_ (.A1(_02946_),
    .A2(_02963_),
    .B1(_02966_),
    .Y(_03127_));
 sky130_fd_sc_hd__nand2_4 _11345_ (.A(_03126_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__o21bai_4 _11346_ (.A1(_03124_),
    .A2(_03125_),
    .B1_N(_03127_),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(_03128_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__o211ai_2 _11348_ (.A1(_02747_),
    .A2(_02969_),
    .B1(_02944_),
    .C1(_02754_),
    .Y(_03132_));
 sky130_fd_sc_hd__o211ai_4 _11349_ (.A1(_02748_),
    .A2(_02970_),
    .B1(_02945_),
    .C1(_02753_),
    .Y(_03133_));
 sky130_fd_sc_hd__o211ai_1 _11350_ (.A1(_02747_),
    .A2(_02969_),
    .B1(_03131_),
    .C1(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__o211ai_2 _11351_ (.A1(_02748_),
    .A2(_02970_),
    .B1(_03130_),
    .C1(_03132_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand3b_1 _11352_ (.A_N(_03131_),
    .B(_03132_),
    .C(_02973_),
    .Y(_03136_));
 sky130_fd_sc_hd__o2111ai_2 _11353_ (.A1(_02747_),
    .A2(_02969_),
    .B1(_03128_),
    .C1(_03130_),
    .D1(_03133_),
    .Y(_03137_));
 sky130_fd_sc_hd__o211ai_2 _11354_ (.A1(_02748_),
    .A2(_02970_),
    .B1(_03131_),
    .C1(_03132_),
    .Y(_03138_));
 sky130_fd_sc_hd__nand3_2 _11355_ (.A(_03114_),
    .B(_03137_),
    .C(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__nand3_1 _11356_ (.A(_03134_),
    .B(_03136_),
    .C(_03113_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand3_1 _11357_ (.A(_03076_),
    .B(_03139_),
    .C(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__a21o_1 _11358_ (.A1(_03139_),
    .A2(_03141_),
    .B1(_03076_),
    .X(_03143_));
 sky130_fd_sc_hd__and4b_2 _11359_ (.A_N(_03076_),
    .B(_03114_),
    .C(_03137_),
    .D(_03138_),
    .X(_03144_));
 sky130_fd_sc_hd__a21boi_2 _11360_ (.A1(_03076_),
    .A2(_03139_),
    .B1_N(_03141_),
    .Y(_03145_));
 sky130_fd_sc_hd__inv_2 _11361_ (.A(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__and4_1 _11362_ (.A(_03076_),
    .B(_03134_),
    .C(_03136_),
    .D(_03113_),
    .X(_03147_));
 sky130_fd_sc_hd__o21ai_2 _11363_ (.A1(_03147_),
    .A2(_03145_),
    .B1(_03048_),
    .Y(_03148_));
 sky130_fd_sc_hd__o221a_1 _11364_ (.A1(_03076_),
    .A2(_03139_),
    .B1(_03147_),
    .B2(_03145_),
    .C1(_03048_),
    .X(_03149_));
 sky130_fd_sc_hd__a21oi_4 _11365_ (.A1(_03142_),
    .A2(_03143_),
    .B1(_03048_),
    .Y(_03150_));
 sky130_fd_sc_hd__a21oi_4 _11366_ (.A1(_03002_),
    .A2(_02997_),
    .B1(_02999_),
    .Y(_03152_));
 sky130_fd_sc_hd__or3_1 _11367_ (.A(_03152_),
    .B(_03150_),
    .C(_03149_),
    .X(_03153_));
 sky130_fd_sc_hd__o21ai_1 _11368_ (.A1(_03149_),
    .A2(_03150_),
    .B1(_03152_),
    .Y(_03154_));
 sky130_fd_sc_hd__and2_2 _11369_ (.A(_03153_),
    .B(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__a21oi_1 _11370_ (.A1(_03046_),
    .A2(_03047_),
    .B1(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__a21o_1 _11371_ (.A1(_03046_),
    .A2(_03047_),
    .B1(_03155_),
    .X(_03157_));
 sky130_fd_sc_hd__nand3_1 _11372_ (.A(_03046_),
    .B(_03047_),
    .C(_03155_),
    .Y(_03158_));
 sky130_fd_sc_hd__o21a_1 _11373_ (.A1(_02847_),
    .A2(_02872_),
    .B1(_02849_),
    .X(_03159_));
 sky130_fd_sc_hd__a31o_1 _11374_ (.A1(_02861_),
    .A2(net33),
    .A3(_02858_),
    .B1(_02862_),
    .X(_03160_));
 sky130_fd_sc_hd__a32o_1 _11375_ (.A1(_02133_),
    .A2(net139),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_01631_),
    .X(_03161_));
 sky130_fd_sc_hd__nand4_4 _11376_ (.A(_02240_),
    .B(_02356_),
    .C(_01631_),
    .D(_02133_),
    .Y(_03163_));
 sky130_fd_sc_hd__o2111ai_2 _11377_ (.A1(_01238_),
    .A2(_01249_),
    .B1(_02633_),
    .C1(_03161_),
    .D1(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__a22oi_1 _11378_ (.A1(_01303_),
    .A2(_02633_),
    .B1(_03161_),
    .B2(_03163_),
    .Y(_03165_));
 sky130_fd_sc_hd__a32o_1 _11379_ (.A1(_01303_),
    .A2(_02629_),
    .A3(_02631_),
    .B1(_03161_),
    .B2(_03163_),
    .X(_03166_));
 sky130_fd_sc_hd__a32o_1 _11380_ (.A1(_00911_),
    .A2(_02854_),
    .A3(_02856_),
    .B1(_03164_),
    .B2(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__o2111ai_1 _11381_ (.A1(_00856_),
    .A2(_00878_),
    .B1(_02858_),
    .C1(_03164_),
    .D1(_03166_),
    .Y(_03168_));
 sky130_fd_sc_hd__a21bo_1 _11382_ (.A1(_03167_),
    .A2(_03168_),
    .B1_N(_02860_),
    .X(_03169_));
 sky130_fd_sc_hd__nand3b_1 _11383_ (.A_N(_02860_),
    .B(_03167_),
    .C(_03168_),
    .Y(_03170_));
 sky130_fd_sc_hd__inv_2 _11384_ (.A(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__nor2_2 _11385_ (.A(net19),
    .B(net20),
    .Y(_03172_));
 sky130_fd_sc_hd__nand3_4 _11386_ (.A(_02235_),
    .B(_02626_),
    .C(_03172_),
    .Y(_03174_));
 sky130_fd_sc_hd__a21oi_4 _11387_ (.A1(_03174_),
    .A2(net25),
    .B1(net21),
    .Y(_03175_));
 sky130_fd_sc_hd__a21o_4 _11388_ (.A1(_03174_),
    .A2(net25),
    .B1(net21),
    .X(_03176_));
 sky130_fd_sc_hd__o311a_4 _11389_ (.A1(net19),
    .A2(net20),
    .A3(_02627_),
    .B1(net21),
    .C1(net25),
    .X(_03177_));
 sky130_fd_sc_hd__o211ai_4 _11390_ (.A1(net20),
    .A2(_02851_),
    .B1(net21),
    .C1(net25),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_8 _11391_ (.A(_03176_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__nor2_8 _11392_ (.A(_03175_),
    .B(_03177_),
    .Y(_03180_));
 sky130_fd_sc_hd__a32o_1 _11393_ (.A1(net33),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_03169_),
    .B2(_03170_),
    .X(_03181_));
 sky130_fd_sc_hd__nand4_1 _11394_ (.A(_03169_),
    .B(_03170_),
    .C(_03180_),
    .D(net33),
    .Y(_03182_));
 sky130_fd_sc_hd__a21oi_1 _11395_ (.A1(_03181_),
    .A2(_03182_),
    .B1(_03160_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand3_1 _11396_ (.A(_03181_),
    .B(_03182_),
    .C(_03160_),
    .Y(_03185_));
 sky130_fd_sc_hd__and2b_1 _11397_ (.A_N(_03183_),
    .B(_03185_),
    .X(_03186_));
 sky130_fd_sc_hd__a21boi_2 _11398_ (.A1(_02868_),
    .A2(_02869_),
    .B1_N(_02867_),
    .Y(_03187_));
 sky130_fd_sc_hd__xnor2_2 _11399_ (.A(_03186_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__a31o_1 _11400_ (.A1(_05436_),
    .A2(_01222_),
    .A3(_02801_),
    .B1(_02802_),
    .X(_03189_));
 sky130_fd_sc_hd__o221a_1 _11401_ (.A1(_05359_),
    .A2(_05370_),
    .B1(_01396_),
    .B2(_01403_),
    .C1(_01400_),
    .X(_03190_));
 sky130_fd_sc_hd__o211ai_4 _11402_ (.A1(_00003_),
    .A2(_00004_),
    .B1(net147),
    .C1(net146),
    .Y(_03191_));
 sky130_fd_sc_hd__o21ai_1 _11403_ (.A1(_07512_),
    .A2(_00903_),
    .B1(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__and4_1 _11404_ (.A(_00569_),
    .B(_00904_),
    .C(_07513_),
    .D(_00010_),
    .X(_03193_));
 sky130_fd_sc_hd__nand4_1 _11405_ (.A(_00569_),
    .B(_00904_),
    .C(_07513_),
    .D(_00010_),
    .Y(_03194_));
 sky130_fd_sc_hd__a22o_1 _11406_ (.A1(net151),
    .A2(net141),
    .B1(_03192_),
    .B2(_03194_),
    .X(_03196_));
 sky130_fd_sc_hd__nand4_1 _11407_ (.A(net151),
    .B(net141),
    .C(_03192_),
    .D(_03194_),
    .Y(_03197_));
 sky130_fd_sc_hd__a32o_1 _11408_ (.A1(_06309_),
    .A2(_06320_),
    .A3(_01222_),
    .B1(_03196_),
    .B2(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__o2111ai_1 _11409_ (.A1(_06265_),
    .A2(_06287_),
    .B1(_01222_),
    .C1(_03196_),
    .D1(_03197_),
    .Y(_03199_));
 sky130_fd_sc_hd__nand2_1 _11410_ (.A(_03198_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__a21boi_1 _11411_ (.A1(_03198_),
    .A2(_03199_),
    .B1_N(_02799_),
    .Y(_03201_));
 sky130_fd_sc_hd__nand2_1 _11412_ (.A(_02799_),
    .B(_03200_),
    .Y(_03202_));
 sky130_fd_sc_hd__nor2_1 _11413_ (.A(_02799_),
    .B(_03200_),
    .Y(_03203_));
 sky130_fd_sc_hd__a311o_1 _11414_ (.A1(_05392_),
    .A2(_05414_),
    .A3(_01405_),
    .B1(_03201_),
    .C1(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__o21ai_1 _11415_ (.A1(_03201_),
    .A2(_03203_),
    .B1(_03190_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_1 _11416_ (.A(_03204_),
    .B(_03205_),
    .Y(_03207_));
 sky130_fd_sc_hd__nand2_1 _11417_ (.A(_03189_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__nor2_1 _11418_ (.A(_03189_),
    .B(_03207_),
    .Y(_03209_));
 sky130_fd_sc_hd__a311o_1 _11419_ (.A1(_05436_),
    .A2(_01222_),
    .A3(_02801_),
    .B1(_02802_),
    .C1(_03207_),
    .X(_03210_));
 sky130_fd_sc_hd__o21a_1 _11420_ (.A1(_02807_),
    .A2(_02810_),
    .B1(_02808_),
    .X(_03211_));
 sky130_fd_sc_hd__and3b_1 _11421_ (.A_N(_03211_),
    .B(_03210_),
    .C(_03208_),
    .X(_03212_));
 sky130_fd_sc_hd__a21boi_1 _11422_ (.A1(_03208_),
    .A2(_03210_),
    .B1_N(_03211_),
    .Y(_03213_));
 sky130_fd_sc_hd__or2_1 _11423_ (.A(_03212_),
    .B(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__o32a_1 _11424_ (.A1(net155),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(net158),
    .X(_03215_));
 sky130_fd_sc_hd__a311o_1 _11425_ (.A1(net156),
    .A2(_01820_),
    .A3(_01821_),
    .B1(net155),
    .C1(_01589_),
    .X(_03216_));
 sky130_fd_sc_hd__a311o_1 _11426_ (.A1(_04726_),
    .A2(_01585_),
    .A3(_01588_),
    .B1(_01822_),
    .C1(net158),
    .X(_03218_));
 sky130_fd_sc_hd__a22oi_1 _11427_ (.A1(_02866_),
    .A2(_02054_),
    .B1(_03216_),
    .B2(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__nand4_1 _11428_ (.A(_02866_),
    .B(_02054_),
    .C(_03216_),
    .D(_03218_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2b_1 _11429_ (.A_N(_03219_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__a21oi_1 _11430_ (.A1(_02816_),
    .A2(_02825_),
    .B1(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__o211ai_2 _11431_ (.A1(_02582_),
    .A2(_02814_),
    .B1(_02825_),
    .C1(_03221_),
    .Y(_03223_));
 sky130_fd_sc_hd__nand2b_1 _11432_ (.A_N(_03222_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__o31a_1 _11433_ (.A1(net159),
    .A2(_01822_),
    .A3(_02819_),
    .B1(_02818_),
    .X(_03225_));
 sky130_fd_sc_hd__xnor2_1 _11434_ (.A(_03224_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__o31a_1 _11435_ (.A1(_02122_),
    .A2(_02053_),
    .A3(_02829_),
    .B1(_02831_),
    .X(_03227_));
 sky130_fd_sc_hd__nor2_2 _11436_ (.A(_03226_),
    .B(_03227_),
    .Y(_03229_));
 sky130_fd_sc_hd__and2_1 _11437_ (.A(_03226_),
    .B(_03227_),
    .X(_03230_));
 sky130_fd_sc_hd__nor2_1 _11438_ (.A(_03229_),
    .B(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__o211ai_1 _11439_ (.A1(_02841_),
    .A2(_02842_),
    .B1(_02839_),
    .C1(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__a21o_1 _11440_ (.A1(_02839_),
    .A2(_02845_),
    .B1(_03231_),
    .X(_03233_));
 sky130_fd_sc_hd__a211o_1 _11441_ (.A1(_02839_),
    .A2(_02845_),
    .B1(_03229_),
    .C1(_03230_),
    .X(_03234_));
 sky130_fd_sc_hd__o221a_1 _11442_ (.A1(_02835_),
    .A2(_02837_),
    .B1(_03229_),
    .B2(_03230_),
    .C1(_02845_),
    .X(_03235_));
 sky130_fd_sc_hd__nand3b_1 _11443_ (.A_N(_03214_),
    .B(_03232_),
    .C(_03233_),
    .Y(_03236_));
 sky130_fd_sc_hd__nand3b_1 _11444_ (.A_N(_03235_),
    .B(_03214_),
    .C(_03234_),
    .Y(_03237_));
 sky130_fd_sc_hd__a21bo_1 _11445_ (.A1(_03236_),
    .A2(_03237_),
    .B1_N(_03188_),
    .X(_03238_));
 sky130_fd_sc_hd__nand3b_1 _11446_ (.A_N(_03188_),
    .B(_03236_),
    .C(_03237_),
    .Y(_03240_));
 sky130_fd_sc_hd__a21boi_2 _11447_ (.A1(_03237_),
    .A2(_03188_),
    .B1_N(_03236_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand3_1 _11448_ (.A(_03159_),
    .B(_03238_),
    .C(_03240_),
    .Y(_03242_));
 sky130_fd_sc_hd__a21o_1 _11449_ (.A1(_03238_),
    .A2(_03240_),
    .B1(_03159_),
    .X(_03243_));
 sky130_fd_sc_hd__nand2_1 _11450_ (.A(_03242_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand2_1 _11451_ (.A(_02875_),
    .B(_02880_),
    .Y(_03245_));
 sky130_fd_sc_hd__xor2_2 _11452_ (.A(_03244_),
    .B(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__nand3_1 _11453_ (.A(_03157_),
    .B(_03158_),
    .C(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__a21o_1 _11454_ (.A1(_03157_),
    .A2(_03158_),
    .B1(_03246_),
    .X(_03248_));
 sky130_fd_sc_hd__or3_1 _11455_ (.A(_02879_),
    .B(_02881_),
    .C(_03005_),
    .X(_03249_));
 sky130_fd_sc_hd__o211ai_2 _11456_ (.A1(_03005_),
    .A2(_03008_),
    .B1(_03247_),
    .C1(_03248_),
    .Y(_03250_));
 sky130_fd_sc_hd__a22o_1 _11457_ (.A1(_03247_),
    .A2(_03248_),
    .B1(_03249_),
    .B2(_03007_),
    .X(_03251_));
 sky130_fd_sc_hd__nand2_1 _11458_ (.A(_03250_),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__o211ai_2 _11459_ (.A1(_02573_),
    .A2(_02786_),
    .B1(_03014_),
    .C1(_03016_),
    .Y(_03253_));
 sky130_fd_sc_hd__a31o_1 _11460_ (.A1(_02788_),
    .A2(_03014_),
    .A3(_03016_),
    .B1(_03013_),
    .X(_03254_));
 sky130_fd_sc_hd__xnor2_2 _11461_ (.A(_03252_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__xnor2_1 _11462_ (.A(_03024_),
    .B(_03255_),
    .Y(net85));
 sky130_fd_sc_hd__a2bb2o_1 _11463_ (.A1_N(_00812_),
    .A2_N(_00823_),
    .B1(_03023_),
    .B2(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__o211ai_4 _11464_ (.A1(_02795_),
    .A2(_03012_),
    .B1(_03250_),
    .C1(_03253_),
    .Y(_03257_));
 sky130_fd_sc_hd__o21ai_1 _11465_ (.A1(_03246_),
    .A2(_03156_),
    .B1(_03158_),
    .Y(_03258_));
 sky130_fd_sc_hd__inv_2 _11466_ (.A(_03258_),
    .Y(_03260_));
 sky130_fd_sc_hd__o32a_1 _11467_ (.A1(net143),
    .A2(_00532_),
    .A3(_03027_),
    .B1(_00192_),
    .B2(_00274_),
    .X(_03261_));
 sky130_fd_sc_hd__or4_1 _11468_ (.A(_00361_),
    .B(_00363_),
    .C(_00428_),
    .D(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__o32a_1 _11469_ (.A1(net143),
    .A2(_00532_),
    .A3(_03027_),
    .B1(_00366_),
    .B2(_00428_),
    .X(_03263_));
 sky130_fd_sc_hd__o31a_1 _11470_ (.A1(_00274_),
    .A2(_00532_),
    .A3(_03263_),
    .B1(_03262_),
    .X(_03264_));
 sky130_fd_sc_hd__o21ai_1 _11471_ (.A1(_00274_),
    .A2(_00532_),
    .B1(_03263_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _11472_ (.A(_03264_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__o31a_1 _11473_ (.A1(_00274_),
    .A2(_00532_),
    .A3(_03262_),
    .B1(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__a21boi_2 _11474_ (.A1(_03025_),
    .A2(_03033_),
    .B1_N(_03032_),
    .Y(_03268_));
 sky130_fd_sc_hd__a21oi_2 _11475_ (.A1(_03044_),
    .A2(_03039_),
    .B1(_03040_),
    .Y(_03269_));
 sky130_fd_sc_hd__a21o_1 _11476_ (.A1(_03267_),
    .A2(_03268_),
    .B1(_03269_),
    .X(_03271_));
 sky130_fd_sc_hd__xor2_1 _11477_ (.A(_03267_),
    .B(_03268_),
    .X(_03272_));
 sky130_fd_sc_hd__xnor2_2 _11478_ (.A(_03269_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__o2111ai_4 _11479_ (.A1(_02908_),
    .A2(_02909_),
    .B1(_03045_),
    .C1(_03273_),
    .D1(_02685_),
    .Y(_03274_));
 sky130_fd_sc_hd__a31o_1 _11480_ (.A1(_02685_),
    .A2(_02911_),
    .A3(_03045_),
    .B1(_03273_),
    .X(_03275_));
 sky130_fd_sc_hd__o21a_1 _11481_ (.A1(_03072_),
    .A2(_03070_),
    .B1(_03069_),
    .X(_03276_));
 sky130_fd_sc_hd__or4_1 _11482_ (.A(_00188_),
    .B(_00190_),
    .C(_00576_),
    .D(_00578_),
    .X(_03277_));
 sky130_fd_sc_hd__o31a_1 _11483_ (.A1(net149),
    .A2(_00744_),
    .A3(_03055_),
    .B1(_03057_),
    .X(_03278_));
 sky130_fd_sc_hd__a32o_1 _11484_ (.A1(_07540_),
    .A2(_01034_),
    .A3(_01036_),
    .B1(_00743_),
    .B2(_00072_),
    .X(_03279_));
 sky130_fd_sc_hd__nand4_1 _11485_ (.A(_00743_),
    .B(_01038_),
    .C(_07540_),
    .D(_00072_),
    .Y(_03280_));
 sky130_fd_sc_hd__nand2_1 _11486_ (.A(_03279_),
    .B(_03280_),
    .Y(_03282_));
 sky130_fd_sc_hd__o2111ai_1 _11487_ (.A1(_07125_),
    .A2(_07135_),
    .B1(_05316_),
    .C1(_01269_),
    .D1(_01271_),
    .Y(_03283_));
 sky130_fd_sc_hd__nor2_1 _11488_ (.A(_03283_),
    .B(_01542_),
    .Y(_03284_));
 sky130_fd_sc_hd__nand4_2 _11489_ (.A(_03050_),
    .B(_01544_),
    .C(_01269_),
    .D(_07200_),
    .Y(_03285_));
 sky130_fd_sc_hd__a221o_1 _11490_ (.A1(_05294_),
    .A2(_05305_),
    .B1(_01535_),
    .B2(_01537_),
    .C1(_01540_),
    .X(_03286_));
 sky130_fd_sc_hd__o32a_1 _11491_ (.A1(_05327_),
    .A2(_01538_),
    .A3(_01540_),
    .B1(_07189_),
    .B2(_01272_),
    .X(_03287_));
 sky130_fd_sc_hd__a32o_1 _11492_ (.A1(_05316_),
    .A2(_01539_),
    .A3(_01541_),
    .B1(_07200_),
    .B2(_01273_),
    .X(_03288_));
 sky130_fd_sc_hd__o221ai_4 _11493_ (.A1(_01181_),
    .A2(_01182_),
    .B1(_03284_),
    .B2(_03287_),
    .C1(_07440_),
    .Y(_03289_));
 sky130_fd_sc_hd__o211ai_2 _11494_ (.A1(_07441_),
    .A2(_01188_),
    .B1(_03285_),
    .C1(_03288_),
    .Y(_03290_));
 sky130_fd_sc_hd__nand3_2 _11495_ (.A(_03282_),
    .B(_03289_),
    .C(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__a21o_1 _11496_ (.A1(_03289_),
    .A2(_03290_),
    .B1(_03282_),
    .X(_03293_));
 sky130_fd_sc_hd__nand2_1 _11497_ (.A(_03049_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__nand3_1 _11498_ (.A(_03049_),
    .B(_03291_),
    .C(_03293_),
    .Y(_03295_));
 sky130_fd_sc_hd__a21o_1 _11499_ (.A1(_03291_),
    .A2(_03293_),
    .B1(_03049_),
    .X(_03296_));
 sky130_fd_sc_hd__nand3_1 _11500_ (.A(_03278_),
    .B(_03295_),
    .C(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__a21o_1 _11501_ (.A1(_03295_),
    .A2(_03296_),
    .B1(_03278_),
    .X(_03298_));
 sky130_fd_sc_hd__a32o_1 _11502_ (.A1(_00189_),
    .A2(_00191_),
    .A3(_00581_),
    .B1(_03297_),
    .B2(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__o2111ai_1 _11503_ (.A1(_00186_),
    .A2(_00187_),
    .B1(_00581_),
    .C1(_03297_),
    .D1(_03298_),
    .Y(_03300_));
 sky130_fd_sc_hd__nand2_1 _11504_ (.A(_03299_),
    .B(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__o31a_1 _11505_ (.A1(_00067_),
    .A2(_00069_),
    .A3(_00580_),
    .B1(_03062_),
    .X(_03302_));
 sky130_fd_sc_hd__a311o_1 _11506_ (.A1(_02983_),
    .A2(_03058_),
    .A3(_03059_),
    .B1(_03302_),
    .C1(_03301_),
    .X(_03304_));
 sky130_fd_sc_hd__o311a_1 _11507_ (.A1(net148),
    .A2(_00580_),
    .A3(_03060_),
    .B1(_03062_),
    .C1(_03301_),
    .X(_03305_));
 sky130_fd_sc_hd__o21ai_2 _11508_ (.A1(_03276_),
    .A2(_03305_),
    .B1(_03304_),
    .Y(_03306_));
 sky130_fd_sc_hd__a21o_1 _11509_ (.A1(_03276_),
    .A2(_03305_),
    .B1(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__o41a_1 _11510_ (.A1(_03060_),
    .A2(_03276_),
    .A3(_03301_),
    .A4(_03302_),
    .B1(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__and3_1 _11511_ (.A(_02614_),
    .B(_02625_),
    .C(_02097_),
    .X(_03309_));
 sky130_fd_sc_hd__a31o_1 _11512_ (.A1(_01499_),
    .A2(_03097_),
    .A3(_02432_),
    .B1(_03093_),
    .X(_03310_));
 sky130_fd_sc_hd__nor2_2 _11513_ (.A(net52),
    .B(net53),
    .Y(_03311_));
 sky130_fd_sc_hd__nand4_4 _11514_ (.A(_02090_),
    .B(_02688_),
    .C(_03078_),
    .D(_00758_),
    .Y(_03312_));
 sky130_fd_sc_hd__a31oi_4 _11515_ (.A1(net138),
    .A2(_02917_),
    .A3(_03311_),
    .B1(_00299_),
    .Y(_03313_));
 sky130_fd_sc_hd__nor2_4 _11516_ (.A(_00299_),
    .B(_00780_),
    .Y(_03315_));
 sky130_fd_sc_hd__o21ai_4 _11517_ (.A1(net53),
    .A2(_03079_),
    .B1(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__a21oi_4 _11518_ (.A1(_03312_),
    .A2(net173),
    .B1(net54),
    .Y(_03317_));
 sky130_fd_sc_hd__a21o_4 _11519_ (.A1(_03312_),
    .A2(net173),
    .B1(net54),
    .X(_03318_));
 sky130_fd_sc_hd__a21o_4 _11520_ (.A1(_03312_),
    .A2(_03315_),
    .B1(_03317_),
    .X(_03319_));
 sky130_fd_sc_hd__a21oi_4 _11521_ (.A1(_03312_),
    .A2(_03315_),
    .B1(_03317_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand3_4 _11522_ (.A(_03318_),
    .B(net1),
    .C(_03316_),
    .Y(_03321_));
 sky130_fd_sc_hd__o31ai_4 _11523_ (.A1(_00987_),
    .A2(_03081_),
    .A3(_03083_),
    .B1(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__o21ai_1 _11524_ (.A1(_03090_),
    .A2(_03319_),
    .B1(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__o21ai_1 _11525_ (.A1(net166),
    .A2(_02925_),
    .B1(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__o2111ai_1 _11526_ (.A1(_03090_),
    .A2(_03319_),
    .B1(_03322_),
    .C1(_02926_),
    .D1(net164),
    .Y(_03326_));
 sky130_fd_sc_hd__and3_1 _11527_ (.A(net164),
    .B(_02926_),
    .C(_03323_),
    .X(_03327_));
 sky130_fd_sc_hd__o211ai_1 _11528_ (.A1(_01095_),
    .A2(_01117_),
    .B1(_02926_),
    .C1(_03323_),
    .Y(_03328_));
 sky130_fd_sc_hd__o221ai_2 _11529_ (.A1(net166),
    .A2(_02925_),
    .B1(_03090_),
    .B2(_03319_),
    .C1(_03322_),
    .Y(_03329_));
 sky130_fd_sc_hd__o32a_1 _11530_ (.A1(_01488_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_01958_),
    .B2(_02433_),
    .X(_03330_));
 sky130_fd_sc_hd__and3_1 _11531_ (.A(_01969_),
    .B(_02693_),
    .C(_02695_),
    .X(_03331_));
 sky130_fd_sc_hd__and3_1 _11532_ (.A(_03077_),
    .B(_02697_),
    .C(_01969_),
    .X(_03332_));
 sky130_fd_sc_hd__a21oi_1 _11533_ (.A1(_03077_),
    .A2(_03331_),
    .B1(_03330_),
    .Y(_03333_));
 sky130_fd_sc_hd__a31o_1 _11534_ (.A1(_01969_),
    .A2(_02697_),
    .A3(_03077_),
    .B1(_03330_),
    .X(_03334_));
 sky130_fd_sc_hd__nand3_1 _11535_ (.A(_03324_),
    .B(_03326_),
    .C(_03333_),
    .Y(_03335_));
 sky130_fd_sc_hd__o21ai_1 _11536_ (.A1(_03330_),
    .A2(_03332_),
    .B1(_03329_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand3_1 _11537_ (.A(_03328_),
    .B(_03329_),
    .C(_03334_),
    .Y(_03338_));
 sky130_fd_sc_hd__a21oi_1 _11538_ (.A1(_03335_),
    .A2(_03338_),
    .B1(_03091_),
    .Y(_03339_));
 sky130_fd_sc_hd__and3_1 _11539_ (.A(_03338_),
    .B(_03091_),
    .C(_03335_),
    .X(_03340_));
 sky130_fd_sc_hd__o211ai_1 _11540_ (.A1(_03337_),
    .A2(_03327_),
    .B1(_03091_),
    .C1(_03335_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand3b_2 _11541_ (.A_N(_03339_),
    .B(_03341_),
    .C(_03310_),
    .Y(_03342_));
 sky130_fd_sc_hd__o21bai_2 _11542_ (.A1(_03339_),
    .A2(_03340_),
    .B1_N(_03310_),
    .Y(_03343_));
 sky130_fd_sc_hd__a21oi_1 _11543_ (.A1(_03342_),
    .A2(_03343_),
    .B1(_03309_),
    .Y(_03344_));
 sky130_fd_sc_hd__a32o_1 _11544_ (.A1(_02614_),
    .A2(_02625_),
    .A3(_02097_),
    .B1(_03342_),
    .B2(_03343_),
    .X(_03345_));
 sky130_fd_sc_hd__and3_1 _11545_ (.A(_03342_),
    .B(_03343_),
    .C(_03309_),
    .X(_03346_));
 sky130_fd_sc_hd__o31a_1 _11546_ (.A1(_01958_),
    .A2(_02096_),
    .A3(_03100_),
    .B1(_03102_),
    .X(_03348_));
 sky130_fd_sc_hd__o21ai_1 _11547_ (.A1(_03344_),
    .A2(_03346_),
    .B1(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__a31oi_1 _11548_ (.A1(_03342_),
    .A2(_03343_),
    .A3(_03309_),
    .B1(_03348_),
    .Y(_03350_));
 sky130_fd_sc_hd__a21bo_1 _11549_ (.A1(_03345_),
    .A2(_03350_),
    .B1_N(_03349_),
    .X(_03351_));
 sky130_fd_sc_hd__a31oi_1 _11550_ (.A1(_03103_),
    .A2(_03104_),
    .A3(_03105_),
    .B1(_03110_),
    .Y(_03352_));
 sky130_fd_sc_hd__a32o_1 _11551_ (.A1(_03103_),
    .A2(_03104_),
    .A3(_03105_),
    .B1(_03109_),
    .B2(_03110_),
    .X(_03353_));
 sky130_fd_sc_hd__xnor2_1 _11552_ (.A(_03351_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__or4_1 _11553_ (.A(_04244_),
    .B(_01538_),
    .C(_01540_),
    .D(_03116_),
    .X(_03355_));
 sky130_fd_sc_hd__a211oi_1 _11554_ (.A1(_02955_),
    .A2(_03355_),
    .B1(_03906_),
    .C1(_01882_),
    .Y(_03356_));
 sky130_fd_sc_hd__a211o_1 _11555_ (.A1(_02955_),
    .A2(_03355_),
    .B1(_03906_),
    .C1(_01882_),
    .X(_03357_));
 sky130_fd_sc_hd__o32a_1 _11556_ (.A1(_04244_),
    .A2(_01542_),
    .A3(_03116_),
    .B1(_01882_),
    .B2(_03906_),
    .X(_03359_));
 sky130_fd_sc_hd__o32a_2 _11557_ (.A1(_04244_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_03356_),
    .B2(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__nor4_2 _11558_ (.A(_04244_),
    .B(_01662_),
    .C(_03356_),
    .D(_03359_),
    .Y(_03361_));
 sky130_fd_sc_hd__nor2_2 _11559_ (.A(_03360_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__or2_2 _11560_ (.A(_03360_),
    .B(_03361_),
    .X(_03363_));
 sky130_fd_sc_hd__o21bai_1 _11561_ (.A1(_03120_),
    .A2(_03121_),
    .B1_N(_03123_),
    .Y(_03364_));
 sky130_fd_sc_hd__a21boi_4 _11562_ (.A1(_03120_),
    .A2(_03121_),
    .B1_N(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__inv_2 _11563_ (.A(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__nor2_1 _11564_ (.A(_03363_),
    .B(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__or3_1 _11565_ (.A(_03360_),
    .B(_03361_),
    .C(_03366_),
    .X(_03368_));
 sky130_fd_sc_hd__o21a_1 _11566_ (.A1(_03360_),
    .A2(_03361_),
    .B1(_03366_),
    .X(_03370_));
 sky130_fd_sc_hd__nor2_1 _11567_ (.A(_03367_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__o211ai_4 _11568_ (.A1(_02747_),
    .A2(_02969_),
    .B1(_03128_),
    .C1(_03133_),
    .Y(_03372_));
 sky130_fd_sc_hd__o221ai_1 _11569_ (.A1(_03126_),
    .A2(_03127_),
    .B1(_03367_),
    .B2(_03370_),
    .C1(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__nand3_1 _11570_ (.A(_03128_),
    .B(_03135_),
    .C(_03371_),
    .Y(_03374_));
 sky130_fd_sc_hd__o211ai_1 _11571_ (.A1(_03126_),
    .A2(_03127_),
    .B1(_03371_),
    .C1(_03372_),
    .Y(_03375_));
 sky130_fd_sc_hd__o211ai_1 _11572_ (.A1(_03367_),
    .A2(_03370_),
    .B1(_03128_),
    .C1(_03135_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand3_1 _11573_ (.A(_03375_),
    .B(_03376_),
    .C(_03354_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand3b_1 _11574_ (.A_N(_03354_),
    .B(_03373_),
    .C(_03374_),
    .Y(_03378_));
 sky130_fd_sc_hd__a21oi_1 _11575_ (.A1(_03377_),
    .A2(_03378_),
    .B1(_03308_),
    .Y(_03379_));
 sky130_fd_sc_hd__o2111a_1 _11576_ (.A1(_03276_),
    .A2(_03304_),
    .B1(_03307_),
    .C1(_03377_),
    .D1(_03378_),
    .X(_03381_));
 sky130_fd_sc_hd__a21bo_1 _11577_ (.A1(_03308_),
    .A2(_03377_),
    .B1_N(_03378_),
    .X(_03382_));
 sky130_fd_sc_hd__a31o_2 _11578_ (.A1(_03308_),
    .A2(_03377_),
    .A3(_03378_),
    .B1(_03379_),
    .X(_03383_));
 sky130_fd_sc_hd__o21ai_1 _11579_ (.A1(_03379_),
    .A2(_03381_),
    .B1(_03146_),
    .Y(_03384_));
 sky130_fd_sc_hd__xor2_2 _11580_ (.A(_03146_),
    .B(_03383_),
    .X(_03385_));
 sky130_fd_sc_hd__o22ai_4 _11581_ (.A1(_03144_),
    .A2(_03148_),
    .B1(_03150_),
    .B2(_03152_),
    .Y(_03386_));
 sky130_fd_sc_hd__xor2_4 _11582_ (.A(_03385_),
    .B(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__nand3_1 _11583_ (.A(_03274_),
    .B(_03275_),
    .C(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__a21o_1 _11584_ (.A1(_03274_),
    .A2(_03275_),
    .B1(_03387_),
    .X(_03389_));
 sky130_fd_sc_hd__o21ai_1 _11585_ (.A1(_06331_),
    .A2(_01221_),
    .B1(_03197_),
    .Y(_03390_));
 sky130_fd_sc_hd__o22ai_1 _11586_ (.A1(_06331_),
    .A2(_01406_),
    .B1(_01221_),
    .B2(net152),
    .Y(_03392_));
 sky130_fd_sc_hd__nand4_2 _11587_ (.A(_01405_),
    .B(_01222_),
    .C(net151),
    .D(_06341_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(_03392_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__or4_1 _11589_ (.A(_07508_),
    .B(_07510_),
    .C(_01054_),
    .D(_01056_),
    .X(_03395_));
 sky130_fd_sc_hd__o2111ai_4 _11590_ (.A1(_00142_),
    .A2(_00144_),
    .B1(_00148_),
    .C1(_00899_),
    .D1(_00902_),
    .Y(_03396_));
 sky130_fd_sc_hd__nor2_1 _11591_ (.A(_03191_),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__or4_1 _11592_ (.A(net144),
    .B(_00898_),
    .C(_00901_),
    .D(_03191_),
    .X(_03398_));
 sky130_fd_sc_hd__o2111ai_4 _11593_ (.A1(_00142_),
    .A2(_00144_),
    .B1(_00148_),
    .C1(_00565_),
    .D1(_00566_),
    .Y(_03399_));
 sky130_fd_sc_hd__o31a_1 _11594_ (.A1(_00009_),
    .A2(_00898_),
    .A3(_00901_),
    .B1(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__a32o_1 _11595_ (.A1(_00010_),
    .A2(_00899_),
    .A3(_00902_),
    .B1(_00569_),
    .B2(_00150_),
    .X(_03401_));
 sky130_fd_sc_hd__o211ai_1 _11596_ (.A1(_03397_),
    .A2(_03400_),
    .B1(_07513_),
    .C1(net141),
    .Y(_03403_));
 sky130_fd_sc_hd__o221ai_2 _11597_ (.A1(_07512_),
    .A2(_01058_),
    .B1(_03191_),
    .B2(_03396_),
    .C1(_03401_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand3_1 _11598_ (.A(_03394_),
    .B(_03403_),
    .C(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__a21o_1 _11599_ (.A1(_03403_),
    .A2(_03404_),
    .B1(_03394_),
    .X(_03406_));
 sky130_fd_sc_hd__o2bb2ai_1 _11600_ (.A1_N(_03405_),
    .A2_N(_03406_),
    .B1(_02798_),
    .B2(_03191_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand3_1 _11601_ (.A(_03406_),
    .B(_03193_),
    .C(_03405_),
    .Y(_03408_));
 sky130_fd_sc_hd__nand4_1 _11602_ (.A(_03196_),
    .B(_03390_),
    .C(_03407_),
    .D(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__a22oi_1 _11603_ (.A1(_03196_),
    .A2(_03390_),
    .B1(_03407_),
    .B2(_03408_),
    .Y(_03410_));
 sky130_fd_sc_hd__a22o_1 _11604_ (.A1(_03196_),
    .A2(_03390_),
    .B1(_03407_),
    .B2(_03408_),
    .X(_03411_));
 sky130_fd_sc_hd__a32o_1 _11605_ (.A1(_05436_),
    .A2(_01585_),
    .A3(_01588_),
    .B1(_03409_),
    .B2(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__o2111ai_1 _11606_ (.A1(_05359_),
    .A2(_05370_),
    .B1(_01590_),
    .C1(_03409_),
    .D1(_03411_),
    .Y(_03414_));
 sky130_fd_sc_hd__a31o_1 _11607_ (.A1(_05392_),
    .A2(_05414_),
    .A3(_01405_),
    .B1(_03203_),
    .X(_03415_));
 sky130_fd_sc_hd__a221o_1 _11608_ (.A1(_03190_),
    .A2(_03202_),
    .B1(_03412_),
    .B2(_03414_),
    .C1(_03203_),
    .X(_03416_));
 sky130_fd_sc_hd__nand4_1 _11609_ (.A(_03202_),
    .B(_03412_),
    .C(_03414_),
    .D(_03415_),
    .Y(_03417_));
 sky130_fd_sc_hd__a21oi_1 _11610_ (.A1(_03208_),
    .A2(_03211_),
    .B1(_03209_),
    .Y(_03418_));
 sky130_fd_sc_hd__a21oi_1 _11611_ (.A1(_03416_),
    .A2(_03417_),
    .B1(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand3_1 _11612_ (.A(_03416_),
    .B(_03417_),
    .C(_03418_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand2b_1 _11613_ (.A_N(_03419_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__o32ai_1 _11614_ (.A1(net159),
    .A2(_02053_),
    .A3(_03215_),
    .B1(net158),
    .B2(_01589_),
    .Y(_03422_));
 sky130_fd_sc_hd__or4b_1 _11615_ (.A(_04671_),
    .B(_04693_),
    .C(_01822_),
    .D_N(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__o32a_1 _11616_ (.A1(net159),
    .A2(_02053_),
    .A3(_03215_),
    .B1(net155),
    .B2(_01822_),
    .X(_03425_));
 sky130_fd_sc_hd__a31o_1 _11617_ (.A1(_04726_),
    .A2(_01823_),
    .A3(_03422_),
    .B1(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__o21ai_1 _11618_ (.A1(net158),
    .A2(_02053_),
    .B1(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__or4_1 _11619_ (.A(_03479_),
    .B(_03522_),
    .C(_02053_),
    .D(_03426_),
    .X(_03428_));
 sky130_fd_sc_hd__and2_1 _11620_ (.A(_03427_),
    .B(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__o21ai_2 _11621_ (.A1(_03222_),
    .A2(_03225_),
    .B1(_03223_),
    .Y(_03430_));
 sky130_fd_sc_hd__nand2_1 _11622_ (.A(_03429_),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__or2_2 _11623_ (.A(_03429_),
    .B(_03430_),
    .X(_03432_));
 sky130_fd_sc_hd__nand2_1 _11624_ (.A(_03431_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__a21oi_1 _11625_ (.A1(_03226_),
    .A2(_03227_),
    .B1(_02838_),
    .Y(_03434_));
 sky130_fd_sc_hd__a21oi_1 _11626_ (.A1(_02845_),
    .A2(_03434_),
    .B1(_03229_),
    .Y(_03436_));
 sky130_fd_sc_hd__a221oi_1 _11627_ (.A1(_03431_),
    .A2(_03432_),
    .B1(_02845_),
    .B2(_03434_),
    .C1(_03229_),
    .Y(_03437_));
 sky130_fd_sc_hd__a221o_1 _11628_ (.A1(_03431_),
    .A2(_03432_),
    .B1(_02845_),
    .B2(_03434_),
    .C1(_03229_),
    .X(_03438_));
 sky130_fd_sc_hd__nor2_1 _11629_ (.A(_03433_),
    .B(_03436_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand3b_1 _11630_ (.A_N(_03436_),
    .B(_03432_),
    .C(_03431_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21ai_1 _11631_ (.A1(_03437_),
    .A2(_03439_),
    .B1(_03421_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand3b_1 _11632_ (.A_N(_03421_),
    .B(_03438_),
    .C(_03440_),
    .Y(_03442_));
 sky130_fd_sc_hd__nand4_4 _11633_ (.A(_02235_),
    .B(_02626_),
    .C(_03172_),
    .D(_00769_),
    .Y(_03443_));
 sky130_fd_sc_hd__o311a_4 _11634_ (.A1(net20),
    .A2(net21),
    .A3(_02851_),
    .B1(net22),
    .C1(net25),
    .X(_03444_));
 sky130_fd_sc_hd__o211ai_4 _11635_ (.A1(net21),
    .A2(_03174_),
    .B1(net22),
    .C1(net25),
    .Y(_03445_));
 sky130_fd_sc_hd__a21oi_4 _11636_ (.A1(_03443_),
    .A2(net25),
    .B1(net22),
    .Y(_03447_));
 sky130_fd_sc_hd__a21o_4 _11637_ (.A1(_03443_),
    .A2(net25),
    .B1(net22),
    .X(_03448_));
 sky130_fd_sc_hd__nand2_8 _11638_ (.A(_03445_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__nor2_8 _11639_ (.A(_03444_),
    .B(_03447_),
    .Y(_03450_));
 sky130_fd_sc_hd__o31a_1 _11640_ (.A1(_00900_),
    .A2(_02857_),
    .A3(_03165_),
    .B1(_03164_),
    .X(_03451_));
 sky130_fd_sc_hd__a32o_1 _11641_ (.A1(_00911_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_01303_),
    .B2(_02858_),
    .X(_03452_));
 sky130_fd_sc_hd__nand4_2 _11642_ (.A(_00911_),
    .B(_01303_),
    .C(_02858_),
    .D(_03180_),
    .Y(_03453_));
 sky130_fd_sc_hd__or4_1 _11643_ (.A(_01576_),
    .B(_01598_),
    .C(_02628_),
    .D(_02630_),
    .X(_03454_));
 sky130_fd_sc_hd__nand4_2 _11644_ (.A(_02240_),
    .B(_02356_),
    .C(_02133_),
    .D(_02866_),
    .Y(_03455_));
 sky130_fd_sc_hd__o211ai_4 _11645_ (.A1(net168),
    .A2(net163),
    .B1(net139),
    .C1(_02237_),
    .Y(_03456_));
 sky130_fd_sc_hd__o32a_1 _11646_ (.A1(_02122_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(net159),
    .B2(_02241_),
    .X(_03458_));
 sky130_fd_sc_hd__a32o_1 _11647_ (.A1(_02866_),
    .A2(net139),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_02133_),
    .X(_03459_));
 sky130_fd_sc_hd__a32o_1 _11648_ (.A1(_01631_),
    .A2(_02629_),
    .A3(_02631_),
    .B1(_03455_),
    .B2(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__nand4_1 _11649_ (.A(_01631_),
    .B(_02633_),
    .C(_03455_),
    .D(_03459_),
    .Y(_03461_));
 sky130_fd_sc_hd__a22o_1 _11650_ (.A1(_03452_),
    .A2(_03453_),
    .B1(_03460_),
    .B2(_03461_),
    .X(_03462_));
 sky130_fd_sc_hd__nand4_1 _11651_ (.A(_03452_),
    .B(_03453_),
    .C(_03460_),
    .D(_03461_),
    .Y(_03463_));
 sky130_fd_sc_hd__nand2_1 _11652_ (.A(_03163_),
    .B(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand3_1 _11653_ (.A(_03163_),
    .B(_03462_),
    .C(_03463_),
    .Y(_03465_));
 sky130_fd_sc_hd__a21o_1 _11654_ (.A1(_03462_),
    .A2(_03463_),
    .B1(_03163_),
    .X(_03466_));
 sky130_fd_sc_hd__nand3_1 _11655_ (.A(_03451_),
    .B(_03465_),
    .C(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__a21o_1 _11656_ (.A1(_03465_),
    .A2(_03466_),
    .B1(_03451_),
    .X(_03469_));
 sky130_fd_sc_hd__a32o_1 _11657_ (.A1(net33),
    .A2(_03445_),
    .A3(_03448_),
    .B1(_03467_),
    .B2(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__nand4_1 _11658_ (.A(_03450_),
    .B(_03467_),
    .C(_03469_),
    .D(net33),
    .Y(_03471_));
 sky130_fd_sc_hd__a31o_1 _11659_ (.A1(net33),
    .A2(_03169_),
    .A3(_03180_),
    .B1(_03171_),
    .X(_03472_));
 sky130_fd_sc_hd__nand3_1 _11660_ (.A(_03470_),
    .B(_03471_),
    .C(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__a21o_1 _11661_ (.A1(_03470_),
    .A2(_03471_),
    .B1(_03472_),
    .X(_03474_));
 sky130_fd_sc_hd__a21oi_1 _11662_ (.A1(_03185_),
    .A2(_03187_),
    .B1(_03183_),
    .Y(_03475_));
 sky130_fd_sc_hd__a21oi_1 _11663_ (.A1(_03473_),
    .A2(_03474_),
    .B1(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__and3_1 _11664_ (.A(_03473_),
    .B(_03474_),
    .C(_03475_),
    .X(_03477_));
 sky130_fd_sc_hd__nor2_1 _11665_ (.A(_03476_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__nand3_1 _11666_ (.A(_03441_),
    .B(_03442_),
    .C(_03478_),
    .Y(_03480_));
 sky130_fd_sc_hd__a21o_1 _11667_ (.A1(_03441_),
    .A2(_03442_),
    .B1(_03478_),
    .X(_03481_));
 sky130_fd_sc_hd__nand2_1 _11668_ (.A(_03480_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__or2_1 _11669_ (.A(_03241_),
    .B(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__nand2_1 _11670_ (.A(_03241_),
    .B(_03482_),
    .Y(_03484_));
 sky130_fd_sc_hd__and2_1 _11671_ (.A(_03483_),
    .B(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__nand3_1 _11672_ (.A(_02875_),
    .B(_02880_),
    .C(_03243_),
    .Y(_03486_));
 sky130_fd_sc_hd__nand2_1 _11673_ (.A(_03242_),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__xor2_2 _11674_ (.A(_03485_),
    .B(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__and3_1 _11675_ (.A(_03388_),
    .B(_03389_),
    .C(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__a21oi_1 _11676_ (.A1(_03388_),
    .A2(_03389_),
    .B1(_03488_),
    .Y(_03491_));
 sky130_fd_sc_hd__nor2_1 _11677_ (.A(_03489_),
    .B(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__o211a_1 _11678_ (.A1(_03156_),
    .A2(_03246_),
    .B1(_03158_),
    .C1(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__or3_2 _11679_ (.A(_03258_),
    .B(_03489_),
    .C(_03491_),
    .X(_03494_));
 sky130_fd_sc_hd__o21a_1 _11680_ (.A1(_03489_),
    .A2(_03491_),
    .B1(_03258_),
    .X(_03495_));
 sky130_fd_sc_hd__a211o_1 _11681_ (.A1(_03251_),
    .A2(_03257_),
    .B1(_03493_),
    .C1(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__o211ai_1 _11682_ (.A1(_03493_),
    .A2(_03495_),
    .B1(_03251_),
    .C1(_03257_),
    .Y(_03497_));
 sky130_fd_sc_hd__o211a_1 _11683_ (.A1(_03260_),
    .A2(_03492_),
    .B1(_03251_),
    .C1(_03257_),
    .X(_03498_));
 sky130_fd_sc_hd__o211ai_2 _11684_ (.A1(_03260_),
    .A2(_03492_),
    .B1(_03251_),
    .C1(_03257_),
    .Y(_03499_));
 sky130_fd_sc_hd__nand2_1 _11685_ (.A(_03496_),
    .B(_03497_),
    .Y(_03500_));
 sky130_fd_sc_hd__xor2_1 _11686_ (.A(_03256_),
    .B(_03500_),
    .X(net86));
 sky130_fd_sc_hd__and3_1 _11687_ (.A(_03023_),
    .B(_03255_),
    .C(_03500_),
    .X(_03502_));
 sky130_fd_sc_hd__a31o_1 _11688_ (.A1(_03023_),
    .A2(_03255_),
    .A3(_03500_),
    .B1(_00834_),
    .X(_03503_));
 sky130_fd_sc_hd__a21boi_2 _11689_ (.A1(_03388_),
    .A2(_03488_),
    .B1_N(_03389_),
    .Y(_03504_));
 sky130_fd_sc_hd__a21bo_1 _11690_ (.A1(_03441_),
    .A2(_03478_),
    .B1_N(_03442_),
    .X(_03505_));
 sky130_fd_sc_hd__o31a_1 _11691_ (.A1(net158),
    .A2(_02053_),
    .A3(_03425_),
    .B1(_03423_),
    .X(_03506_));
 sky130_fd_sc_hd__o31a_1 _11692_ (.A1(_04671_),
    .A2(_04693_),
    .A3(_02053_),
    .B1(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__o21ai_1 _11693_ (.A1(net155),
    .A2(_02053_),
    .B1(_03506_),
    .Y(_03508_));
 sky130_fd_sc_hd__nor4_2 _11694_ (.A(_04671_),
    .B(_04693_),
    .C(_02053_),
    .D(_03506_),
    .Y(_03509_));
 sky130_fd_sc_hd__a221o_1 _11695_ (.A1(_03429_),
    .A2(_03430_),
    .B1(_02845_),
    .B2(_03434_),
    .C1(_03229_),
    .X(_03510_));
 sky130_fd_sc_hd__o221ai_2 _11696_ (.A1(_03429_),
    .A2(_03430_),
    .B1(_03507_),
    .B2(_03509_),
    .C1(_03510_),
    .Y(_03512_));
 sky130_fd_sc_hd__a211o_1 _11697_ (.A1(_03432_),
    .A2(_03510_),
    .B1(_03509_),
    .C1(_03507_),
    .X(_03513_));
 sky130_fd_sc_hd__o31a_1 _11698_ (.A1(_05425_),
    .A2(_01589_),
    .A3(_03410_),
    .B1(_03409_),
    .X(_03514_));
 sky130_fd_sc_hd__a21boi_1 _11699_ (.A1(_03193_),
    .A2(_03405_),
    .B1_N(_03406_),
    .Y(_03515_));
 sky130_fd_sc_hd__a211oi_1 _11700_ (.A1(_03395_),
    .A2(_03398_),
    .B1(_03400_),
    .C1(_03393_),
    .Y(_03516_));
 sky130_fd_sc_hd__a211o_1 _11701_ (.A1(_03395_),
    .A2(_03398_),
    .B1(_03400_),
    .C1(_03393_),
    .X(_03517_));
 sky130_fd_sc_hd__o311a_1 _11702_ (.A1(_07512_),
    .A2(_01058_),
    .A3(_03400_),
    .B1(_03398_),
    .C1(_03393_),
    .X(_03518_));
 sky130_fd_sc_hd__a21o_1 _11703_ (.A1(_01214_),
    .A2(_01215_),
    .B1(_07512_),
    .X(_03519_));
 sky130_fd_sc_hd__a22o_2 _11704_ (.A1(_00267_),
    .A2(_00269_),
    .B1(_00567_),
    .B2(_00568_),
    .X(_03520_));
 sky130_fd_sc_hd__o21ai_2 _11705_ (.A1(_00274_),
    .A2(_00570_),
    .B1(_03396_),
    .Y(_03521_));
 sky130_fd_sc_hd__o211ai_4 _11706_ (.A1(_00266_),
    .A2(_00268_),
    .B1(_00899_),
    .C1(_00902_),
    .Y(_03523_));
 sky130_fd_sc_hd__and4_1 _11707_ (.A(_00569_),
    .B(_00904_),
    .C(_00150_),
    .D(_00275_),
    .X(_03524_));
 sky130_fd_sc_hd__o21ai_1 _11708_ (.A1(_03399_),
    .A2(_03523_),
    .B1(_03521_),
    .Y(_03525_));
 sky130_fd_sc_hd__o21ai_2 _11709_ (.A1(_00009_),
    .A2(_01058_),
    .B1(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__o2111ai_4 _11710_ (.A1(_03399_),
    .A2(_03523_),
    .B1(_03521_),
    .C1(_00010_),
    .D1(net141),
    .Y(_03527_));
 sky130_fd_sc_hd__o211ai_1 _11711_ (.A1(_07512_),
    .A2(_01221_),
    .B1(_03526_),
    .C1(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__a221o_1 _11712_ (.A1(_01214_),
    .A2(_01215_),
    .B1(_03526_),
    .B2(_03527_),
    .C1(_07512_),
    .X(_03529_));
 sky130_fd_sc_hd__a2bb2o_1 _11713_ (.A1_N(_03516_),
    .A2_N(_03518_),
    .B1(_03528_),
    .B2(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__or4bb_1 _11714_ (.A(_03516_),
    .B(_03518_),
    .C_N(_03528_),
    .D_N(_03529_),
    .X(_03531_));
 sky130_fd_sc_hd__a21o_1 _11715_ (.A1(_03530_),
    .A2(_03531_),
    .B1(_03515_),
    .X(_03532_));
 sky130_fd_sc_hd__nand3_1 _11716_ (.A(_03515_),
    .B(_03530_),
    .C(_03531_),
    .Y(_03534_));
 sky130_fd_sc_hd__and3_1 _11717_ (.A(_06341_),
    .B(_01585_),
    .C(_01588_),
    .X(_03535_));
 sky130_fd_sc_hd__and3_1 _11718_ (.A(_03535_),
    .B(net151),
    .C(_01405_),
    .X(_03536_));
 sky130_fd_sc_hd__or4_1 _11719_ (.A(_06331_),
    .B(net152),
    .C(_01406_),
    .D(_01589_),
    .X(_03537_));
 sky130_fd_sc_hd__o32a_2 _11720_ (.A1(_06331_),
    .A2(_01584_),
    .A3(_01586_),
    .B1(net152),
    .B2(_01406_),
    .X(_03538_));
 sky130_fd_sc_hd__o211a_1 _11721_ (.A1(_03536_),
    .A2(_03538_),
    .B1(_05436_),
    .C1(_01823_),
    .X(_03539_));
 sky130_fd_sc_hd__a311oi_1 _11722_ (.A1(_05436_),
    .A2(_01820_),
    .A3(_01821_),
    .B1(_03536_),
    .C1(_03538_),
    .Y(_03540_));
 sky130_fd_sc_hd__nor2_1 _11723_ (.A(_03539_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__and3_1 _11724_ (.A(_03532_),
    .B(_03534_),
    .C(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__a21oi_1 _11725_ (.A1(_03532_),
    .A2(_03534_),
    .B1(_03541_),
    .Y(_03543_));
 sky130_fd_sc_hd__nor2_1 _11726_ (.A(_03542_),
    .B(_03543_),
    .Y(_03545_));
 sky130_fd_sc_hd__nor2_1 _11727_ (.A(_03514_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand2_1 _11728_ (.A(_03545_),
    .B(_03514_),
    .Y(_03547_));
 sky130_fd_sc_hd__nand2b_1 _11729_ (.A_N(_03546_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__a21bo_1 _11730_ (.A1(_03416_),
    .A2(_03418_),
    .B1_N(_03417_),
    .X(_03549_));
 sky130_fd_sc_hd__xor2_1 _11731_ (.A(_03548_),
    .B(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__a21o_1 _11732_ (.A1(_03512_),
    .A2(_03513_),
    .B1(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__nand3_1 _11733_ (.A(_03512_),
    .B(_03513_),
    .C(_03550_),
    .Y(_03552_));
 sky130_fd_sc_hd__a311o_1 _11734_ (.A1(_03451_),
    .A2(_03465_),
    .A3(_03466_),
    .B1(_03449_),
    .C1(_00310_),
    .X(_03553_));
 sky130_fd_sc_hd__o311a_1 _11735_ (.A1(_01620_),
    .A2(_02632_),
    .A3(_03458_),
    .B1(_03455_),
    .C1(_03453_),
    .X(_03554_));
 sky130_fd_sc_hd__o311ai_1 _11736_ (.A1(_01620_),
    .A2(_02632_),
    .A3(_03458_),
    .B1(_03455_),
    .C1(_03453_),
    .Y(_03556_));
 sky130_fd_sc_hd__a211o_1 _11737_ (.A1(_03454_),
    .A2(_03455_),
    .B1(_03458_),
    .C1(_03453_),
    .X(_03557_));
 sky130_fd_sc_hd__a22o_4 _11738_ (.A1(_01543_),
    .A2(_01565_),
    .B1(_02852_),
    .B2(_02853_),
    .X(_03558_));
 sky130_fd_sc_hd__o32ai_4 _11739_ (.A1(net159),
    .A2(_02353_),
    .A3(_02354_),
    .B1(net158),
    .B2(_02241_),
    .Y(_03559_));
 sky130_fd_sc_hd__o21ai_4 _11740_ (.A1(_02350_),
    .A2(_02351_),
    .B1(net156),
    .Y(_03560_));
 sky130_fd_sc_hd__and4_1 _11741_ (.A(_02240_),
    .B(_02356_),
    .C(_02866_),
    .D(net156),
    .X(_03561_));
 sky130_fd_sc_hd__or4_1 _11742_ (.A(net158),
    .B(_02353_),
    .C(_02354_),
    .D(_03456_),
    .X(_03562_));
 sky130_fd_sc_hd__o21ai_1 _11743_ (.A1(_03456_),
    .A2(_03560_),
    .B1(_03559_),
    .Y(_03563_));
 sky130_fd_sc_hd__o2111ai_4 _11744_ (.A1(_03456_),
    .A2(_03560_),
    .B1(_03559_),
    .C1(_02133_),
    .D1(_02633_),
    .Y(_03564_));
 sky130_fd_sc_hd__o31a_1 _11745_ (.A1(_02079_),
    .A2(_02100_),
    .A3(_02632_),
    .B1(_03563_),
    .X(_03565_));
 sky130_fd_sc_hd__o21ai_1 _11746_ (.A1(_02122_),
    .A2(_02632_),
    .B1(_03563_),
    .Y(_03567_));
 sky130_fd_sc_hd__a32o_1 _11747_ (.A1(_01631_),
    .A2(_02854_),
    .A3(_02856_),
    .B1(_03564_),
    .B2(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__o2111ai_2 _11748_ (.A1(_01532_),
    .A2(_01554_),
    .B1(_02858_),
    .C1(_03564_),
    .D1(_03567_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _11749_ (.A(_03568_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__a22o_1 _11750_ (.A1(_03556_),
    .A2(_03557_),
    .B1(_03568_),
    .B2(_03569_),
    .X(_03571_));
 sky130_fd_sc_hd__or3b_1 _11751_ (.A(_03554_),
    .B(_03570_),
    .C_N(_03557_),
    .X(_03572_));
 sky130_fd_sc_hd__nand4_2 _11752_ (.A(_03462_),
    .B(_03464_),
    .C(_03571_),
    .D(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__a22o_1 _11753_ (.A1(_03462_),
    .A2(_03464_),
    .B1(_03571_),
    .B2(_03572_),
    .X(_03574_));
 sky130_fd_sc_hd__a32o_1 _11754_ (.A1(_01303_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_03450_),
    .B2(_00911_),
    .X(_03575_));
 sky130_fd_sc_hd__or3_1 _11755_ (.A(_01292_),
    .B(_03444_),
    .C(_03447_),
    .X(_03576_));
 sky130_fd_sc_hd__and4_1 _11756_ (.A(_00911_),
    .B(_01303_),
    .C(_03180_),
    .D(_03450_),
    .X(_03578_));
 sky130_fd_sc_hd__o31a_1 _11757_ (.A1(_00900_),
    .A2(_03179_),
    .A3(_03576_),
    .B1(_03575_),
    .X(_03579_));
 sky130_fd_sc_hd__nand4b_4 _11758_ (.A_N(_02851_),
    .B(_00791_),
    .C(_00769_),
    .D(_00747_),
    .Y(_03580_));
 sky130_fd_sc_hd__o311a_4 _11759_ (.A1(net21),
    .A2(net22),
    .A3(_03174_),
    .B1(net24),
    .C1(net25),
    .X(_03581_));
 sky130_fd_sc_hd__a21oi_4 _11760_ (.A1(_03580_),
    .A2(net25),
    .B1(net24),
    .Y(_03582_));
 sky130_fd_sc_hd__or2_4 _11761_ (.A(_03581_),
    .B(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__nor2_8 _11762_ (.A(_03581_),
    .B(_03582_),
    .Y(_03584_));
 sky130_fd_sc_hd__or3_1 _11763_ (.A(_03582_),
    .B(_00310_),
    .C(_03581_),
    .X(_03585_));
 sky130_fd_sc_hd__xnor2_2 _11764_ (.A(_03579_),
    .B(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__and3_1 _11765_ (.A(_03573_),
    .B(_03574_),
    .C(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__a21oi_1 _11766_ (.A1(_03573_),
    .A2(_03574_),
    .B1(_03586_),
    .Y(_03589_));
 sky130_fd_sc_hd__o211a_1 _11767_ (.A1(_03587_),
    .A2(_03589_),
    .B1(_03469_),
    .C1(_03553_),
    .X(_03590_));
 sky130_fd_sc_hd__a211o_1 _11768_ (.A1(_03469_),
    .A2(_03553_),
    .B1(_03587_),
    .C1(_03589_),
    .X(_03591_));
 sky130_fd_sc_hd__and2b_1 _11769_ (.A_N(_03590_),
    .B(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__a21boi_1 _11770_ (.A1(_03474_),
    .A2(_03475_),
    .B1_N(_03473_),
    .Y(_03593_));
 sky130_fd_sc_hd__xnor2_1 _11771_ (.A(_03592_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__a21o_1 _11772_ (.A1(_03551_),
    .A2(_03552_),
    .B1(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__nand3_1 _11773_ (.A(_03551_),
    .B(_03552_),
    .C(_03594_),
    .Y(_03596_));
 sky130_fd_sc_hd__a21o_1 _11774_ (.A1(_03595_),
    .A2(_03596_),
    .B1(_03505_),
    .X(_03597_));
 sky130_fd_sc_hd__nand3_1 _11775_ (.A(_03595_),
    .B(_03596_),
    .C(_03505_),
    .Y(_03598_));
 sky130_fd_sc_hd__nand3_2 _11776_ (.A(_03242_),
    .B(_03484_),
    .C(_03486_),
    .Y(_03600_));
 sky130_fd_sc_hd__o21ai_1 _11777_ (.A1(_03241_),
    .A2(_03482_),
    .B1(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__a22oi_1 _11778_ (.A1(_03597_),
    .A2(_03598_),
    .B1(_03600_),
    .B2(_03483_),
    .Y(_03602_));
 sky130_fd_sc_hd__o211ai_2 _11779_ (.A1(_03241_),
    .A2(_03482_),
    .B1(_03598_),
    .C1(_03600_),
    .Y(_03603_));
 sky130_fd_sc_hd__o2111ai_1 _11780_ (.A1(_03241_),
    .A2(_03482_),
    .B1(_03597_),
    .C1(_03598_),
    .D1(_03600_),
    .Y(_03604_));
 sky130_fd_sc_hd__nand2b_1 _11781_ (.A_N(_03602_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__or4_2 _11782_ (.A(_04244_),
    .B(_01658_),
    .C(_01660_),
    .D(_03359_),
    .X(_03606_));
 sky130_fd_sc_hd__a211oi_4 _11783_ (.A1(_03357_),
    .A2(_03606_),
    .B1(_04244_),
    .C1(_01882_),
    .Y(_03607_));
 sky130_fd_sc_hd__a211o_1 _11784_ (.A1(_03357_),
    .A2(_03606_),
    .B1(_04244_),
    .C1(_01882_),
    .X(_03608_));
 sky130_fd_sc_hd__o211a_2 _11785_ (.A1(_04244_),
    .A2(_01882_),
    .B1(_03357_),
    .C1(_03606_),
    .X(_03609_));
 sky130_fd_sc_hd__nor2_1 _11786_ (.A(_03607_),
    .B(_03609_),
    .Y(_03611_));
 sky130_fd_sc_hd__o211ai_2 _11787_ (.A1(_03363_),
    .A2(_03366_),
    .B1(_03128_),
    .C1(_03135_),
    .Y(_03612_));
 sky130_fd_sc_hd__o211ai_4 _11788_ (.A1(_03362_),
    .A2(_03365_),
    .B1(_03372_),
    .C1(_03130_),
    .Y(_03613_));
 sky130_fd_sc_hd__o31a_1 _11789_ (.A1(_03360_),
    .A2(_03361_),
    .A3(_03366_),
    .B1(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__o221ai_4 _11790_ (.A1(_03363_),
    .A2(_03366_),
    .B1(_03607_),
    .B2(_03609_),
    .C1(_03613_),
    .Y(_03615_));
 sky130_fd_sc_hd__o211ai_2 _11791_ (.A1(_03362_),
    .A2(_03365_),
    .B1(_03611_),
    .C1(_03612_),
    .Y(_03616_));
 sky130_fd_sc_hd__o221ai_2 _11792_ (.A1(_03362_),
    .A2(_03365_),
    .B1(_03607_),
    .B2(_03609_),
    .C1(_03612_),
    .Y(_03617_));
 sky130_fd_sc_hd__o211ai_1 _11793_ (.A1(_03363_),
    .A2(_03366_),
    .B1(_03611_),
    .C1(_03613_),
    .Y(_03618_));
 sky130_fd_sc_hd__o2bb2ai_1 _11794_ (.A1_N(_03350_),
    .A2_N(_03345_),
    .B1(_03108_),
    .B2(_03352_),
    .Y(_03619_));
 sky130_fd_sc_hd__and2_1 _11795_ (.A(_03349_),
    .B(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__a21boi_2 _11796_ (.A1(_03309_),
    .A2(_03343_),
    .B1_N(_03342_),
    .Y(_03622_));
 sky130_fd_sc_hd__and3_1 _11797_ (.A(_02647_),
    .B(_02427_),
    .C(_02428_),
    .X(_03623_));
 sky130_fd_sc_hd__o32a_1 _11798_ (.A1(_01958_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_02636_),
    .B2(_02433_),
    .X(_03624_));
 sky130_fd_sc_hd__or4_1 _11799_ (.A(_01958_),
    .B(_02636_),
    .C(_02433_),
    .D(_02696_),
    .X(_03625_));
 sky130_fd_sc_hd__nand2b_1 _11800_ (.A_N(_03624_),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__o31a_1 _11801_ (.A1(_03906_),
    .A2(_02092_),
    .A3(_02094_),
    .B1(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__nor3_1 _11802_ (.A(_03906_),
    .B(_02096_),
    .C(_03626_),
    .Y(_03628_));
 sky130_fd_sc_hd__or2_1 _11803_ (.A(_03627_),
    .B(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__inv_2 _11804_ (.A(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__o21ai_1 _11805_ (.A1(_02925_),
    .A2(_03090_),
    .B1(_03335_),
    .Y(_03631_));
 sky130_fd_sc_hd__o2bb2a_1 _11806_ (.A1_N(_03092_),
    .A2_N(_03335_),
    .B1(_03337_),
    .B2(_03327_),
    .X(_03633_));
 sky130_fd_sc_hd__o22ai_2 _11807_ (.A1(net166),
    .A2(_02925_),
    .B1(_03090_),
    .B2(_03319_),
    .Y(_03634_));
 sky130_fd_sc_hd__a21oi_1 _11808_ (.A1(_03322_),
    .A2(_03634_),
    .B1(_03332_),
    .Y(_03635_));
 sky130_fd_sc_hd__a22o_1 _11809_ (.A1(_03077_),
    .A2(_03331_),
    .B1(_03634_),
    .B2(_03322_),
    .X(_03636_));
 sky130_fd_sc_hd__and3_1 _11810_ (.A(_03332_),
    .B(_03634_),
    .C(_03322_),
    .X(_03637_));
 sky130_fd_sc_hd__nand4_2 _11811_ (.A(_03322_),
    .B(_03634_),
    .C(_03331_),
    .D(_03077_),
    .Y(_03638_));
 sky130_fd_sc_hd__and3_1 _11812_ (.A(_01499_),
    .B(_02922_),
    .C(_02924_),
    .X(_03639_));
 sky130_fd_sc_hd__o211ai_2 _11813_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_02922_),
    .C1(_02924_),
    .Y(_03640_));
 sky130_fd_sc_hd__and3_1 _11814_ (.A(net164),
    .B(_03082_),
    .C(_03084_),
    .X(_03641_));
 sky130_fd_sc_hd__a21oi_1 _11815_ (.A1(_03312_),
    .A2(_03315_),
    .B1(_00987_),
    .Y(_03642_));
 sky130_fd_sc_hd__o21ai_4 _11816_ (.A1(net54),
    .A2(_03313_),
    .B1(_03642_),
    .Y(_03644_));
 sky130_fd_sc_hd__nand4_4 _11817_ (.A(net138),
    .B(_02917_),
    .C(_03311_),
    .D(_00780_),
    .Y(_03645_));
 sky130_fd_sc_hd__a41oi_4 _11818_ (.A1(net138),
    .A2(_02917_),
    .A3(_03311_),
    .A4(_00780_),
    .B1(_00299_),
    .Y(_03646_));
 sky130_fd_sc_hd__a311o_2 _11819_ (.A1(_02918_),
    .A2(_03311_),
    .A3(_00780_),
    .B1(net56),
    .C1(_00299_),
    .X(_03647_));
 sky130_fd_sc_hd__a21bo_2 _11820_ (.A1(_03645_),
    .A2(net173),
    .B1_N(net56),
    .X(_03648_));
 sky130_fd_sc_hd__o311a_2 _11821_ (.A1(net53),
    .A2(net54),
    .A3(_03079_),
    .B1(net56),
    .C1(net173),
    .X(_03649_));
 sky130_fd_sc_hd__nand2_8 _11822_ (.A(net56),
    .B(_03646_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21o_4 _11823_ (.A1(_03645_),
    .A2(net173),
    .B1(net56),
    .X(_03651_));
 sky130_fd_sc_hd__nand2_8 _11824_ (.A(_03650_),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_8 _11825_ (.A(_03647_),
    .B(_03648_),
    .Y(_03653_));
 sky130_fd_sc_hd__o21a_1 _11826_ (.A1(net56),
    .A2(_03646_),
    .B1(net1),
    .X(_03655_));
 sky130_fd_sc_hd__o21ai_1 _11827_ (.A1(net56),
    .A2(_03646_),
    .B1(net1),
    .Y(_03656_));
 sky130_fd_sc_hd__o21ai_4 _11828_ (.A1(_03649_),
    .A2(_03656_),
    .B1(_03644_),
    .Y(_03657_));
 sky130_fd_sc_hd__o21ai_2 _11829_ (.A1(net56),
    .A2(_03646_),
    .B1(_00998_),
    .Y(_03658_));
 sky130_fd_sc_hd__a31o_2 _11830_ (.A1(net173),
    .A2(net56),
    .A3(_03645_),
    .B1(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__and4_1 _11831_ (.A(_00998_),
    .B(_03320_),
    .C(_03653_),
    .D(net1),
    .X(_03660_));
 sky130_fd_sc_hd__nand3b_2 _11832_ (.A_N(_03644_),
    .B(_03650_),
    .C(_03655_),
    .Y(_03661_));
 sky130_fd_sc_hd__o311a_1 _11833_ (.A1(_03649_),
    .A2(_03658_),
    .A3(_03321_),
    .B1(_03641_),
    .C1(_03657_),
    .X(_03662_));
 sky130_fd_sc_hd__o2111ai_4 _11834_ (.A1(_03321_),
    .A2(_03659_),
    .B1(_03657_),
    .C1(net164),
    .D1(_03087_),
    .Y(_03663_));
 sky130_fd_sc_hd__a21oi_1 _11835_ (.A1(_03657_),
    .A2(_03661_),
    .B1(_03641_),
    .Y(_03664_));
 sky130_fd_sc_hd__a32o_1 _11836_ (.A1(net164),
    .A2(_03082_),
    .A3(_03084_),
    .B1(_03657_),
    .B2(_03661_),
    .X(_03666_));
 sky130_fd_sc_hd__o21ai_1 _11837_ (.A1(_03662_),
    .A2(_03664_),
    .B1(_03639_),
    .Y(_03667_));
 sky130_fd_sc_hd__a211o_1 _11838_ (.A1(_01499_),
    .A2(_02926_),
    .B1(_03662_),
    .C1(_03664_),
    .X(_03668_));
 sky130_fd_sc_hd__o2111ai_4 _11839_ (.A1(_01423_),
    .A2(_01445_),
    .B1(_02926_),
    .C1(_03663_),
    .D1(_03666_),
    .Y(_03669_));
 sky130_fd_sc_hd__o21ai_1 _11840_ (.A1(_03662_),
    .A2(_03664_),
    .B1(_03640_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand4_2 _11841_ (.A(_03636_),
    .B(_03638_),
    .C(_03669_),
    .D(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__o211ai_2 _11842_ (.A1(_03635_),
    .A2(_03637_),
    .B1(_03667_),
    .C1(_03668_),
    .Y(_03672_));
 sky130_fd_sc_hd__and3_1 _11843_ (.A(_03671_),
    .B(_03672_),
    .C(_03633_),
    .X(_03673_));
 sky130_fd_sc_hd__nand4_1 _11844_ (.A(_03338_),
    .B(_03631_),
    .C(_03671_),
    .D(_03672_),
    .Y(_03674_));
 sky130_fd_sc_hd__a21o_1 _11845_ (.A1(_03671_),
    .A2(_03672_),
    .B1(_03633_),
    .X(_03675_));
 sky130_fd_sc_hd__a41o_1 _11846_ (.A1(_03338_),
    .A2(_03631_),
    .A3(_03671_),
    .A4(_03672_),
    .B1(_03630_),
    .X(_03677_));
 sky130_fd_sc_hd__a21o_1 _11847_ (.A1(_03674_),
    .A2(_03675_),
    .B1(_03629_),
    .X(_03678_));
 sky130_fd_sc_hd__nand3_2 _11848_ (.A(_03629_),
    .B(_03674_),
    .C(_03675_),
    .Y(_03679_));
 sky130_fd_sc_hd__nand3_2 _11849_ (.A(_03622_),
    .B(_03678_),
    .C(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__a21oi_2 _11850_ (.A1(_03678_),
    .A2(_03679_),
    .B1(_03622_),
    .Y(_03681_));
 sky130_fd_sc_hd__and4b_1 _11851_ (.A_N(_03620_),
    .B(_03622_),
    .C(_03678_),
    .D(_03679_),
    .X(_03682_));
 sky130_fd_sc_hd__nand3_1 _11852_ (.A(_03349_),
    .B(_03619_),
    .C(_03680_),
    .Y(_03683_));
 sky130_fd_sc_hd__o21ai_2 _11853_ (.A1(_03620_),
    .A2(_03681_),
    .B1(_03680_),
    .Y(_03684_));
 sky130_fd_sc_hd__a21oi_1 _11854_ (.A1(_03620_),
    .A2(_03681_),
    .B1(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__a31o_1 _11855_ (.A1(_03349_),
    .A2(_03619_),
    .A3(_03681_),
    .B1(_03684_),
    .X(_03686_));
 sky130_fd_sc_hd__o2111ai_4 _11856_ (.A1(_03620_),
    .A2(_03680_),
    .B1(_03686_),
    .C1(_03616_),
    .D1(_03615_),
    .Y(_03688_));
 sky130_fd_sc_hd__o211ai_2 _11857_ (.A1(_03682_),
    .A2(_03685_),
    .B1(_03617_),
    .C1(_03618_),
    .Y(_03689_));
 sky130_fd_sc_hd__a32o_1 _11858_ (.A1(_03278_),
    .A2(_03295_),
    .A3(_03296_),
    .B1(_03298_),
    .B2(_03277_),
    .X(_03690_));
 sky130_fd_sc_hd__or4_1 _11859_ (.A(_00361_),
    .B(_00363_),
    .C(_00576_),
    .D(_00578_),
    .X(_03691_));
 sky130_fd_sc_hd__o32a_1 _11860_ (.A1(net148),
    .A2(_01033_),
    .A3(_01035_),
    .B1(_00192_),
    .B2(_00744_),
    .X(_03692_));
 sky130_fd_sc_hd__and4_1 _11861_ (.A(_00743_),
    .B(_01038_),
    .C(_00072_),
    .D(_00193_),
    .X(_03693_));
 sky130_fd_sc_hd__or2_1 _11862_ (.A(_03692_),
    .B(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__xor2_1 _11863_ (.A(_03691_),
    .B(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__or4_1 _11864_ (.A(_07441_),
    .B(_01184_),
    .C(_01186_),
    .D(_03287_),
    .X(_03696_));
 sky130_fd_sc_hd__o311a_1 _11865_ (.A1(_07441_),
    .A2(_01188_),
    .A3(_03287_),
    .B1(_03285_),
    .C1(_03280_),
    .X(_03697_));
 sky130_fd_sc_hd__a21oi_1 _11866_ (.A1(_03285_),
    .A2(_03696_),
    .B1(_03280_),
    .Y(_03699_));
 sky130_fd_sc_hd__o221a_1 _11867_ (.A1(_00321_),
    .A2(_07537_),
    .B1(_01181_),
    .B2(_01182_),
    .C1(_07536_),
    .X(_03700_));
 sky130_fd_sc_hd__and3_1 _11868_ (.A(_01659_),
    .B(net140),
    .C(_05316_),
    .X(_03701_));
 sky130_fd_sc_hd__nand4_1 _11869_ (.A(_05272_),
    .B(_05283_),
    .C(_01659_),
    .D(net140),
    .Y(_03702_));
 sky130_fd_sc_hd__a32o_1 _11870_ (.A1(_05316_),
    .A2(_01659_),
    .A3(net140),
    .B1(_07200_),
    .B2(_01544_),
    .X(_03703_));
 sky130_fd_sc_hd__o211ai_4 _11871_ (.A1(_07125_),
    .A2(_07135_),
    .B1(_01659_),
    .C1(net140),
    .Y(_03704_));
 sky130_fd_sc_hd__and3_1 _11872_ (.A(_03701_),
    .B(_01544_),
    .C(_07200_),
    .X(_03705_));
 sky130_fd_sc_hd__nand4_1 _11873_ (.A(_07200_),
    .B(_01544_),
    .C(_01664_),
    .D(_05316_),
    .Y(_03706_));
 sky130_fd_sc_hd__and3_1 _11874_ (.A(_01269_),
    .B(_01271_),
    .C(_07440_),
    .X(_03707_));
 sky130_fd_sc_hd__o211a_1 _11875_ (.A1(_03286_),
    .A2(_03704_),
    .B1(_03707_),
    .C1(_03703_),
    .X(_03708_));
 sky130_fd_sc_hd__o2111ai_1 _11876_ (.A1(_03286_),
    .A2(_03704_),
    .B1(_07440_),
    .C1(_03703_),
    .D1(_01273_),
    .Y(_03710_));
 sky130_fd_sc_hd__a21oi_1 _11877_ (.A1(_03703_),
    .A2(_03706_),
    .B1(_03707_),
    .Y(_03711_));
 sky130_fd_sc_hd__a32o_1 _11878_ (.A1(_07440_),
    .A2(_01269_),
    .A3(_01271_),
    .B1(_03703_),
    .B2(_03706_),
    .X(_03712_));
 sky130_fd_sc_hd__o21ai_1 _11879_ (.A1(_03708_),
    .A2(_03711_),
    .B1(_03700_),
    .Y(_03713_));
 sky130_fd_sc_hd__o211ai_2 _11880_ (.A1(net149),
    .A2(_01188_),
    .B1(_03710_),
    .C1(_03712_),
    .Y(_03714_));
 sky130_fd_sc_hd__o211ai_1 _11881_ (.A1(_03697_),
    .A2(_03699_),
    .B1(_03713_),
    .C1(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__a211o_1 _11882_ (.A1(_03713_),
    .A2(_03714_),
    .B1(_03697_),
    .C1(_03699_),
    .X(_03716_));
 sky130_fd_sc_hd__a22oi_2 _11883_ (.A1(_03291_),
    .A2(_03294_),
    .B1(_03715_),
    .B2(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__and4_1 _11884_ (.A(_03291_),
    .B(_03294_),
    .C(_03715_),
    .D(_03716_),
    .X(_03718_));
 sky130_fd_sc_hd__nor3_1 _11885_ (.A(_03695_),
    .B(_03717_),
    .C(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__o21a_1 _11886_ (.A1(_03717_),
    .A2(_03718_),
    .B1(_03695_),
    .X(_03721_));
 sky130_fd_sc_hd__nor2_1 _11887_ (.A(_03719_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__and2_1 _11888_ (.A(_03722_),
    .B(_03690_),
    .X(_03723_));
 sky130_fd_sc_hd__nand2_1 _11889_ (.A(_03722_),
    .B(_03690_),
    .Y(_03724_));
 sky130_fd_sc_hd__nor2_1 _11890_ (.A(_03690_),
    .B(_03722_),
    .Y(_03725_));
 sky130_fd_sc_hd__or2_1 _11891_ (.A(_03723_),
    .B(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__xor2_2 _11892_ (.A(_03306_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__nand2b_1 _11893_ (.A_N(_03727_),
    .B(_03689_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand3_1 _11894_ (.A(_03688_),
    .B(_03689_),
    .C(_03727_),
    .Y(_03729_));
 sky130_fd_sc_hd__a21o_1 _11895_ (.A1(_03688_),
    .A2(_03689_),
    .B1(_03727_),
    .X(_03730_));
 sky130_fd_sc_hd__and2_1 _11896_ (.A(_03729_),
    .B(_03730_),
    .X(_03732_));
 sky130_fd_sc_hd__a21oi_1 _11897_ (.A1(_03729_),
    .A2(_03730_),
    .B1(_03382_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand3_1 _11898_ (.A(_03730_),
    .B(_03382_),
    .C(_03729_),
    .Y(_03734_));
 sky130_fd_sc_hd__and2b_1 _11899_ (.A_N(_03733_),
    .B(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__o221ai_4 _11900_ (.A1(_03144_),
    .A2(_03148_),
    .B1(_03150_),
    .B2(_03152_),
    .C1(_03384_),
    .Y(_03736_));
 sky130_fd_sc_hd__o21ai_2 _11901_ (.A1(_03146_),
    .A2(_03383_),
    .B1(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__xor2_4 _11902_ (.A(_03735_),
    .B(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__o21ai_1 _11903_ (.A1(_00428_),
    .A2(_00532_),
    .B1(_03264_),
    .Y(_03739_));
 sky130_fd_sc_hd__or3_2 _11904_ (.A(_00428_),
    .B(_00532_),
    .C(_03264_),
    .X(_03740_));
 sky130_fd_sc_hd__nand2_1 _11905_ (.A(_03739_),
    .B(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__o21ai_2 _11906_ (.A1(_03267_),
    .A2(_03268_),
    .B1(_03271_),
    .Y(_03743_));
 sky130_fd_sc_hd__xor2_2 _11907_ (.A(_03741_),
    .B(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__nand2_1 _11908_ (.A(_03274_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__or2_1 _11909_ (.A(_03744_),
    .B(_03274_),
    .X(_03746_));
 sky130_fd_sc_hd__o21ba_1 _11910_ (.A1(_03744_),
    .A2(_03274_),
    .B1_N(_03738_),
    .X(_03747_));
 sky130_fd_sc_hd__and3b_1 _11911_ (.A_N(_03738_),
    .B(_03745_),
    .C(_03746_),
    .X(_03748_));
 sky130_fd_sc_hd__a21boi_1 _11912_ (.A1(_03745_),
    .A2(_03746_),
    .B1_N(_03738_),
    .Y(_03749_));
 sky130_fd_sc_hd__o21ba_2 _11913_ (.A1(_03605_),
    .A2(_03748_),
    .B1_N(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__inv_2 _11914_ (.A(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__a211o_1 _11915_ (.A1(_03747_),
    .A2(_03745_),
    .B1(_03605_),
    .C1(_03749_),
    .X(_03752_));
 sky130_fd_sc_hd__o21ai_1 _11916_ (.A1(_03748_),
    .A2(_03749_),
    .B1(_03605_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2_2 _11917_ (.A(_03752_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__a211oi_1 _11918_ (.A1(_03494_),
    .A2(_03499_),
    .B1(_03504_),
    .C1(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_2 _11919_ (.A(_03755_),
    .B(_03504_),
    .Y(_03757_));
 sky130_fd_sc_hd__o211ai_4 _11920_ (.A1(_03504_),
    .A2(_03755_),
    .B1(_03494_),
    .C1(_03499_),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_1 _11921_ (.A(_03757_),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__o32a_2 _11922_ (.A1(_03493_),
    .A2(_03498_),
    .A3(_03757_),
    .B1(_03759_),
    .B2(_03756_),
    .X(_03760_));
 sky130_fd_sc_hd__xor2_1 _11923_ (.A(_03503_),
    .B(_03760_),
    .X(net88));
 sky130_fd_sc_hd__nand2_1 _11924_ (.A(_03502_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__nor2_1 _11925_ (.A(_03691_),
    .B(_03692_),
    .Y(_03762_));
 sky130_fd_sc_hd__a31o_1 _11926_ (.A1(_03703_),
    .A2(_03706_),
    .A3(_03707_),
    .B1(_03700_),
    .X(_03764_));
 sky130_fd_sc_hd__a211o_1 _11927_ (.A1(_03712_),
    .A2(_03764_),
    .B1(_03762_),
    .C1(_03693_),
    .X(_03765_));
 sky130_fd_sc_hd__o211ai_4 _11928_ (.A1(_03693_),
    .A2(_03762_),
    .B1(_03764_),
    .C1(_03712_),
    .Y(_03766_));
 sky130_fd_sc_hd__o32a_1 _11929_ (.A1(net148),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_01272_),
    .B2(net149),
    .X(_03767_));
 sky130_fd_sc_hd__and3_1 _11930_ (.A(_03700_),
    .B(_01273_),
    .C(_00072_),
    .X(_03768_));
 sky130_fd_sc_hd__or4_1 _11931_ (.A(net149),
    .B(net148),
    .C(_01188_),
    .D(_01272_),
    .X(_03769_));
 sky130_fd_sc_hd__and3_1 _11932_ (.A(_01541_),
    .B(_07440_),
    .C(_01539_),
    .X(_03770_));
 sky130_fd_sc_hd__nand3_1 _11933_ (.A(net134),
    .B(_05316_),
    .C(_01879_),
    .Y(_03771_));
 sky130_fd_sc_hd__o21ai_1 _11934_ (.A1(_07189_),
    .A2(_01662_),
    .B1(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__o211ai_4 _11935_ (.A1(_07125_),
    .A2(_07135_),
    .B1(net135),
    .C1(_01880_),
    .Y(_03773_));
 sky130_fd_sc_hd__o2bb2ai_1 _11936_ (.A1_N(_03704_),
    .A2_N(_03771_),
    .B1(_03773_),
    .B2(_03702_),
    .Y(_03775_));
 sky130_fd_sc_hd__o21ai_1 _11937_ (.A1(_07441_),
    .A2(_01542_),
    .B1(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__o2111ai_1 _11938_ (.A1(_03702_),
    .A2(_03773_),
    .B1(_07440_),
    .C1(_03772_),
    .D1(_01544_),
    .Y(_03777_));
 sky130_fd_sc_hd__nand2_1 _11939_ (.A(_03775_),
    .B(_03770_),
    .Y(_03778_));
 sky130_fd_sc_hd__a31o_1 _11940_ (.A1(_07440_),
    .A2(_01539_),
    .A3(_01541_),
    .B1(_03775_),
    .X(_03779_));
 sky130_fd_sc_hd__o211ai_2 _11941_ (.A1(_03767_),
    .A2(_03768_),
    .B1(_03778_),
    .C1(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand4b_1 _11942_ (.A_N(_03767_),
    .B(_03769_),
    .C(_03776_),
    .D(_03777_),
    .Y(_03781_));
 sky130_fd_sc_hd__a21o_1 _11943_ (.A1(_03780_),
    .A2(_03781_),
    .B1(_03705_),
    .X(_03782_));
 sky130_fd_sc_hd__nand3_1 _11944_ (.A(_03780_),
    .B(_03781_),
    .C(_03705_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand4_1 _11945_ (.A(_03765_),
    .B(_03766_),
    .C(_03782_),
    .D(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__a22o_1 _11946_ (.A1(_03765_),
    .A2(_03766_),
    .B1(_03782_),
    .B2(_03783_),
    .X(_03786_));
 sky130_fd_sc_hd__a21oi_1 _11947_ (.A1(_03713_),
    .A2(_03714_),
    .B1(_03697_),
    .Y(_03787_));
 sky130_fd_sc_hd__or2_1 _11948_ (.A(_03699_),
    .B(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__a21o_1 _11949_ (.A1(_03784_),
    .A2(_03786_),
    .B1(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__and3_1 _11950_ (.A(_03784_),
    .B(_03786_),
    .C(_03788_),
    .X(_03790_));
 sky130_fd_sc_hd__nand3_1 _11951_ (.A(_03784_),
    .B(_03786_),
    .C(_03788_),
    .Y(_03791_));
 sky130_fd_sc_hd__o32a_1 _11952_ (.A1(_00192_),
    .A2(_01033_),
    .A3(_01035_),
    .B1(_00366_),
    .B2(_00744_),
    .X(_03792_));
 sky130_fd_sc_hd__and4_1 _11953_ (.A(_00743_),
    .B(_01038_),
    .C(_00193_),
    .D(_00367_),
    .X(_03793_));
 sky130_fd_sc_hd__or4_1 _11954_ (.A(_00192_),
    .B(_00366_),
    .C(_00744_),
    .D(_01037_),
    .X(_03794_));
 sky130_fd_sc_hd__o22ai_2 _11955_ (.A1(_00532_),
    .A2(_00580_),
    .B1(_03792_),
    .B2(_03793_),
    .Y(_03795_));
 sky130_fd_sc_hd__or4_2 _11956_ (.A(_00532_),
    .B(_00580_),
    .C(_03792_),
    .D(_03793_),
    .X(_03797_));
 sky130_fd_sc_hd__nand2_1 _11957_ (.A(_03795_),
    .B(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__and3_1 _11958_ (.A(_03789_),
    .B(_03791_),
    .C(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__a21oi_1 _11959_ (.A1(_03789_),
    .A2(_03791_),
    .B1(_03798_),
    .Y(_03800_));
 sky130_fd_sc_hd__nor2_1 _11960_ (.A(_03799_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__nor2_1 _11961_ (.A(_03695_),
    .B(_03718_),
    .Y(_03802_));
 sky130_fd_sc_hd__o21a_1 _11962_ (.A1(_03717_),
    .A2(_03802_),
    .B1(_03801_),
    .X(_03803_));
 sky130_fd_sc_hd__or3_2 _11963_ (.A(_03717_),
    .B(_03801_),
    .C(_03802_),
    .X(_03804_));
 sky130_fd_sc_hd__nand2b_1 _11964_ (.A_N(_03803_),
    .B(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__a21oi_2 _11965_ (.A1(_03306_),
    .A2(_03724_),
    .B1(_03725_),
    .Y(_03806_));
 sky130_fd_sc_hd__xnor2_2 _11966_ (.A(_03805_),
    .B(_03806_),
    .Y(_03808_));
 sky130_fd_sc_hd__or3_2 _11967_ (.A(_04244_),
    .B(_02092_),
    .C(_02094_),
    .X(_03809_));
 sky130_fd_sc_hd__o32a_1 _11968_ (.A1(_02636_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_03906_),
    .B2(_02433_),
    .X(_03810_));
 sky130_fd_sc_hd__a31o_1 _11969_ (.A1(_03917_),
    .A2(_02697_),
    .A3(_03623_),
    .B1(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__xor2_2 _11970_ (.A(_03809_),
    .B(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__nand3_1 _11971_ (.A(_03636_),
    .B(_03669_),
    .C(_03670_),
    .Y(_03813_));
 sky130_fd_sc_hd__o31ai_1 _11972_ (.A1(_03906_),
    .A2(_02096_),
    .A3(_03624_),
    .B1(_03625_),
    .Y(_03814_));
 sky130_fd_sc_hd__a31o_1 _11973_ (.A1(_03661_),
    .A2(_03641_),
    .A3(_03657_),
    .B1(_03639_),
    .X(_03815_));
 sky130_fd_sc_hd__a21o_1 _11974_ (.A1(_03666_),
    .A2(_03815_),
    .B1(_03814_),
    .X(_03816_));
 sky130_fd_sc_hd__nand3_1 _11975_ (.A(_03666_),
    .B(_03814_),
    .C(_03815_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_03816_),
    .B(_03817_),
    .Y(_03819_));
 sky130_fd_sc_hd__and3_1 _11977_ (.A(_01969_),
    .B(_03082_),
    .C(_03084_),
    .X(_03820_));
 sky130_fd_sc_hd__o211ai_2 _11978_ (.A1(_01892_),
    .A2(_01914_),
    .B1(_02922_),
    .C1(_02924_),
    .Y(_03821_));
 sky130_fd_sc_hd__o21ai_1 _11979_ (.A1(_01488_),
    .A2(_03086_),
    .B1(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__o31ai_4 _11980_ (.A1(_01958_),
    .A2(_03086_),
    .A3(_03640_),
    .B1(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__a31o_1 _11981_ (.A1(_03312_),
    .A2(net54),
    .A3(net173),
    .B1(net166),
    .X(_03824_));
 sky130_fd_sc_hd__o22ai_2 _11982_ (.A1(_03317_),
    .A2(_03824_),
    .B1(_03649_),
    .B2(_03658_),
    .Y(_03825_));
 sky130_fd_sc_hd__o2111ai_4 _11983_ (.A1(_00321_),
    .A2(_01139_),
    .B1(_01172_),
    .C1(_03650_),
    .D1(_03651_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand4b_4 _11984_ (.A_N(_03644_),
    .B(_03650_),
    .C(_03651_),
    .D(net164),
    .Y(_03827_));
 sky130_fd_sc_hd__o21ai_1 _11985_ (.A1(_03644_),
    .A2(_03826_),
    .B1(_03825_),
    .Y(_03828_));
 sky130_fd_sc_hd__or2_4 _11986_ (.A(net56),
    .B(_00299_),
    .X(_03830_));
 sky130_fd_sc_hd__nor2_8 _11987_ (.A(_03645_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_4 _11988_ (.A(net53),
    .B(_03830_),
    .C(net54),
    .D(_03079_),
    .X(_03832_));
 sky130_fd_sc_hd__or4_1 _11989_ (.A(_00288_),
    .B(_03830_),
    .C(net54),
    .D(_03312_),
    .X(_03833_));
 sky130_fd_sc_hd__or4_4 _11990_ (.A(_00299_),
    .B(net54),
    .C(net56),
    .D(_03312_),
    .X(_03834_));
 sky130_fd_sc_hd__a22oi_2 _11991_ (.A1(net1),
    .A2(_03831_),
    .B1(_03827_),
    .B2(_03825_),
    .Y(_03835_));
 sky130_fd_sc_hd__a21oi_1 _11992_ (.A1(_03828_),
    .A2(_03833_),
    .B1(_03823_),
    .Y(_03836_));
 sky130_fd_sc_hd__a21o_1 _11993_ (.A1(_03828_),
    .A2(_03833_),
    .B1(_03823_),
    .X(_03837_));
 sky130_fd_sc_hd__o211a_1 _11994_ (.A1(_00288_),
    .A2(_03834_),
    .B1(_03828_),
    .C1(_03823_),
    .X(_03838_));
 sky130_fd_sc_hd__nand2_1 _11995_ (.A(_03835_),
    .B(_03823_),
    .Y(_03839_));
 sky130_fd_sc_hd__o22ai_2 _11996_ (.A1(_03321_),
    .A2(_03659_),
    .B1(_03836_),
    .B2(_03838_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand3_1 _11997_ (.A(_03837_),
    .B(_03839_),
    .C(_03660_),
    .Y(_03842_));
 sky130_fd_sc_hd__nand2_1 _11998_ (.A(_03841_),
    .B(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand3_1 _11999_ (.A(_03816_),
    .B(_03817_),
    .C(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand3_1 _12000_ (.A(_03819_),
    .B(_03841_),
    .C(_03842_),
    .Y(_03845_));
 sky130_fd_sc_hd__nand4_2 _12001_ (.A(_03638_),
    .B(_03813_),
    .C(_03844_),
    .D(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__a22oi_1 _12002_ (.A1(_03638_),
    .A2(_03813_),
    .B1(_03819_),
    .B2(_03843_),
    .Y(_03847_));
 sky130_fd_sc_hd__o21ai_1 _12003_ (.A1(_03819_),
    .A2(_03843_),
    .B1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__nand3_2 _12004_ (.A(_03846_),
    .B(_03848_),
    .C(_03812_),
    .Y(_03849_));
 sky130_fd_sc_hd__a21o_1 _12005_ (.A1(_03846_),
    .A2(_03848_),
    .B1(_03812_),
    .X(_03850_));
 sky130_fd_sc_hd__o2111ai_4 _12006_ (.A1(_03630_),
    .A2(_03673_),
    .B1(_03675_),
    .C1(_03849_),
    .D1(_03850_),
    .Y(_03852_));
 sky130_fd_sc_hd__a22o_1 _12007_ (.A1(_03675_),
    .A2(_03677_),
    .B1(_03849_),
    .B2(_03850_),
    .X(_03853_));
 sky130_fd_sc_hd__a21oi_1 _12008_ (.A1(_03852_),
    .A2(_03853_),
    .B1(_03684_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand3_1 _12009_ (.A(_03684_),
    .B(_03852_),
    .C(_03853_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2b_1 _12010_ (.A_N(_03854_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__inv_2 _12011_ (.A(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__a31oi_1 _12012_ (.A1(_03368_),
    .A2(_03608_),
    .A3(_03613_),
    .B1(_03609_),
    .Y(_03858_));
 sky130_fd_sc_hd__o211ai_2 _12013_ (.A1(_03609_),
    .A2(_03614_),
    .B1(_03608_),
    .C1(_03857_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _12014_ (.A(_03858_),
    .B(_03856_),
    .Y(_03860_));
 sky130_fd_sc_hd__a21bo_1 _12015_ (.A1(_03859_),
    .A2(_03860_),
    .B1_N(_03808_),
    .X(_03861_));
 sky130_fd_sc_hd__nand3b_1 _12016_ (.A_N(_03808_),
    .B(_03859_),
    .C(_03860_),
    .Y(_03863_));
 sky130_fd_sc_hd__a21bo_1 _12017_ (.A1(_03808_),
    .A2(_03860_),
    .B1_N(_03859_),
    .X(_03864_));
 sky130_fd_sc_hd__and2_2 _12018_ (.A(_03861_),
    .B(_03863_),
    .X(_03865_));
 sky130_fd_sc_hd__nand2_2 _12019_ (.A(_03688_),
    .B(_03728_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand3_1 _12020_ (.A(_03861_),
    .B(_03863_),
    .C(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__xnor2_2 _12021_ (.A(_03865_),
    .B(_03866_),
    .Y(_03868_));
 sky130_fd_sc_hd__o211ai_2 _12022_ (.A1(_03146_),
    .A2(_03383_),
    .B1(_03734_),
    .C1(_03736_),
    .Y(_03869_));
 sky130_fd_sc_hd__o21a_2 _12023_ (.A1(_03382_),
    .A2(_03732_),
    .B1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__xor2_4 _12024_ (.A(_03868_),
    .B(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__nand2_1 _12025_ (.A(_03739_),
    .B(_03743_),
    .Y(_03872_));
 sky130_fd_sc_hd__o211ai_4 _12026_ (.A1(_03744_),
    .A2(_03274_),
    .B1(_03740_),
    .C1(_03872_),
    .Y(_03874_));
 sky130_fd_sc_hd__and2_1 _12027_ (.A(_03874_),
    .B(_03871_),
    .X(_03875_));
 sky130_fd_sc_hd__xnor2_1 _12028_ (.A(_03871_),
    .B(_03874_),
    .Y(_03876_));
 sky130_fd_sc_hd__a21boi_1 _12029_ (.A1(_03552_),
    .A2(_03594_),
    .B1_N(_03551_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _12030_ (.A(_03574_),
    .B(_03586_),
    .Y(_03878_));
 sky130_fd_sc_hd__o21a_1 _12031_ (.A1(_03554_),
    .A2(_03570_),
    .B1(_03557_),
    .X(_03879_));
 sky130_fd_sc_hd__o31ai_1 _12032_ (.A1(_00900_),
    .A2(_03179_),
    .A3(_03576_),
    .B1(_03585_),
    .Y(_03880_));
 sky130_fd_sc_hd__a31o_1 _12033_ (.A1(_03575_),
    .A2(_03584_),
    .A3(net33),
    .B1(_03578_),
    .X(_03881_));
 sky130_fd_sc_hd__o21ai_2 _12034_ (.A1(_03558_),
    .A2(_03565_),
    .B1(_03564_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _12035_ (.A(_03881_),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__a21o_1 _12036_ (.A1(_03575_),
    .A2(_03880_),
    .B1(_03882_),
    .X(_03885_));
 sky130_fd_sc_hd__a32o_1 _12037_ (.A1(_01631_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_02133_),
    .B2(_02858_),
    .X(_03886_));
 sky130_fd_sc_hd__a211o_1 _12038_ (.A1(_02046_),
    .A2(_02068_),
    .B1(_03175_),
    .C1(_03177_),
    .X(_03887_));
 sky130_fd_sc_hd__o21ai_1 _12039_ (.A1(_03558_),
    .A2(_03887_),
    .B1(_03886_),
    .Y(_03888_));
 sky130_fd_sc_hd__and3_1 _12040_ (.A(_02866_),
    .B(_02629_),
    .C(_02631_),
    .X(_03889_));
 sky130_fd_sc_hd__o21ai_2 _12041_ (.A1(net155),
    .A2(_02241_),
    .B1(_03560_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand4_4 _12042_ (.A(net156),
    .B(_04726_),
    .C(net139),
    .D(_02237_),
    .Y(_03891_));
 sky130_fd_sc_hd__o21ai_1 _12043_ (.A1(_02355_),
    .A2(_03891_),
    .B1(_03890_),
    .Y(_03892_));
 sky130_fd_sc_hd__o21ai_1 _12044_ (.A1(net159),
    .A2(_02632_),
    .B1(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__o2111ai_4 _12045_ (.A1(_02355_),
    .A2(_03891_),
    .B1(_02633_),
    .C1(_02866_),
    .D1(_03890_),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _12046_ (.A(_03892_),
    .B(_03889_),
    .Y(_03896_));
 sky130_fd_sc_hd__o221ai_2 _12047_ (.A1(net159),
    .A2(_02632_),
    .B1(_03891_),
    .B2(_02355_),
    .C1(_03890_),
    .Y(_03897_));
 sky130_fd_sc_hd__o2111ai_4 _12048_ (.A1(_03558_),
    .A2(_03887_),
    .B1(_03893_),
    .C1(_03894_),
    .D1(_03886_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand3_2 _12049_ (.A(_03888_),
    .B(_03896_),
    .C(_03897_),
    .Y(_03899_));
 sky130_fd_sc_hd__o311a_1 _12050_ (.A1(net159),
    .A2(_02241_),
    .A3(_03560_),
    .B1(_03898_),
    .C1(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__o211ai_1 _12051_ (.A1(_03456_),
    .A2(_03560_),
    .B1(_03898_),
    .C1(_03899_),
    .Y(_03901_));
 sky130_fd_sc_hd__a21oi_1 _12052_ (.A1(_03898_),
    .A2(_03899_),
    .B1(_03562_),
    .Y(_03902_));
 sky130_fd_sc_hd__a21o_1 _12053_ (.A1(_03898_),
    .A2(_03899_),
    .B1(_03562_),
    .X(_03903_));
 sky130_fd_sc_hd__o2bb2ai_1 _12054_ (.A1_N(_03883_),
    .A2_N(_03885_),
    .B1(_03900_),
    .B2(_03902_),
    .Y(_03904_));
 sky130_fd_sc_hd__nand4_2 _12055_ (.A(_03883_),
    .B(_03885_),
    .C(_03901_),
    .D(_03903_),
    .Y(_03905_));
 sky130_fd_sc_hd__a21o_1 _12056_ (.A1(_03904_),
    .A2(_03905_),
    .B1(_03879_),
    .X(_03907_));
 sky130_fd_sc_hd__o2111ai_1 _12057_ (.A1(_03570_),
    .A2(_03554_),
    .B1(_03557_),
    .C1(_03904_),
    .D1(_03905_),
    .Y(_03908_));
 sky130_fd_sc_hd__or4_2 _12058_ (.A(_00900_),
    .B(_03581_),
    .C(_03582_),
    .D(_03576_),
    .X(_03909_));
 sky130_fd_sc_hd__a32o_1 _12059_ (.A1(_01303_),
    .A2(_03445_),
    .A3(_03448_),
    .B1(_03584_),
    .B2(_00911_),
    .X(_03910_));
 sky130_fd_sc_hd__nor4_4 _12060_ (.A(_00321_),
    .B(net22),
    .C(net24),
    .D(_03443_),
    .Y(_03911_));
 sky130_fd_sc_hd__or4_4 _12061_ (.A(_00321_),
    .B(net22),
    .C(net24),
    .D(_03443_),
    .X(_03912_));
 sky130_fd_sc_hd__a22o_1 _12062_ (.A1(net33),
    .A2(_03911_),
    .B1(_03910_),
    .B2(_03909_),
    .X(_03913_));
 sky130_fd_sc_hd__inv_2 _12063_ (.A(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__a21oi_1 _12064_ (.A1(_03907_),
    .A2(_03908_),
    .B1(_03913_),
    .Y(_03915_));
 sky130_fd_sc_hd__and3_1 _12065_ (.A(_03907_),
    .B(_03908_),
    .C(_03913_),
    .X(_03916_));
 sky130_fd_sc_hd__or2_1 _12066_ (.A(_03915_),
    .B(_03916_),
    .X(_03918_));
 sky130_fd_sc_hd__and3_1 _12067_ (.A(_03918_),
    .B(_03878_),
    .C(_03573_),
    .X(_03919_));
 sky130_fd_sc_hd__a21o_1 _12068_ (.A1(_03573_),
    .A2(_03878_),
    .B1(_03918_),
    .X(_03920_));
 sky130_fd_sc_hd__nand2b_1 _12069_ (.A_N(_03919_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__a21o_1 _12070_ (.A1(_03591_),
    .A2(_03593_),
    .B1(_03590_),
    .X(_03922_));
 sky130_fd_sc_hd__xor2_1 _12071_ (.A(_03921_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__nor3_1 _12072_ (.A(_05425_),
    .B(_01822_),
    .C(_03538_),
    .Y(_03924_));
 sky130_fd_sc_hd__o21ai_1 _12073_ (.A1(_07512_),
    .A2(_01221_),
    .B1(_03527_),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _12074_ (.A(_03526_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__o311ai_4 _12075_ (.A1(_05425_),
    .A2(_01822_),
    .A3(_03538_),
    .B1(_03926_),
    .C1(_03537_),
    .Y(_03927_));
 sky130_fd_sc_hd__o211ai_2 _12076_ (.A1(_03536_),
    .A2(_03924_),
    .B1(_03925_),
    .C1(_03526_),
    .Y(_03929_));
 sky130_fd_sc_hd__o32ai_4 _12077_ (.A1(_00009_),
    .A2(_01217_),
    .A3(_01219_),
    .B1(_07512_),
    .B2(net136),
    .Y(_03930_));
 sky130_fd_sc_hd__a211o_1 _12078_ (.A1(_01402_),
    .A2(_01397_),
    .B1(_00009_),
    .C1(_01399_),
    .X(_03931_));
 sky130_fd_sc_hd__o21ai_1 _12079_ (.A1(_03519_),
    .A2(_03931_),
    .B1(_03930_),
    .Y(_03932_));
 sky130_fd_sc_hd__o2111ai_2 _12080_ (.A1(_00299_),
    .A2(_00424_),
    .B1(_00427_),
    .C1(_00565_),
    .D1(_00566_),
    .Y(_03933_));
 sky130_fd_sc_hd__o32a_1 _12081_ (.A1(_00274_),
    .A2(_00898_),
    .A3(_00901_),
    .B1(net142),
    .B2(_00570_),
    .X(_03934_));
 sky130_fd_sc_hd__o21ai_2 _12082_ (.A1(net142),
    .A2(_00570_),
    .B1(_03523_),
    .Y(_03935_));
 sky130_fd_sc_hd__o2111ai_4 _12083_ (.A1(_00299_),
    .A2(_00424_),
    .B1(_00427_),
    .C1(_00899_),
    .D1(_00902_),
    .Y(_03936_));
 sky130_fd_sc_hd__or4_1 _12084_ (.A(net142),
    .B(_00898_),
    .C(_00901_),
    .D(_03520_),
    .X(_03937_));
 sky130_fd_sc_hd__o2bb2ai_1 _12085_ (.A1_N(_03523_),
    .A2_N(_03933_),
    .B1(_03936_),
    .B2(_03520_),
    .Y(_03938_));
 sky130_fd_sc_hd__o21ai_1 _12086_ (.A1(net144),
    .A2(_01058_),
    .B1(_03938_),
    .Y(_03940_));
 sky130_fd_sc_hd__o2111ai_4 _12087_ (.A1(_03520_),
    .A2(_03936_),
    .B1(_03935_),
    .C1(_00150_),
    .D1(net141),
    .Y(_03941_));
 sky130_fd_sc_hd__o2111ai_2 _12088_ (.A1(_00142_),
    .A2(_00144_),
    .B1(_00148_),
    .C1(net141),
    .D1(_03938_),
    .Y(_03942_));
 sky130_fd_sc_hd__o221ai_2 _12089_ (.A1(net144),
    .A2(_01058_),
    .B1(_03520_),
    .B2(_03936_),
    .C1(_03935_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand3_2 _12090_ (.A(_03932_),
    .B(_03942_),
    .C(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__o2111ai_4 _12091_ (.A1(_03519_),
    .A2(_03931_),
    .B1(_03940_),
    .C1(_03941_),
    .D1(_03930_),
    .Y(_03945_));
 sky130_fd_sc_hd__a2bb2o_1 _12092_ (.A1_N(_03396_),
    .A2_N(_03520_),
    .B1(_03944_),
    .B2(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__nand3_1 _12093_ (.A(_03944_),
    .B(_03945_),
    .C(_03524_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand4_1 _12094_ (.A(_03927_),
    .B(_03929_),
    .C(_03946_),
    .D(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__a22o_1 _12095_ (.A1(_03927_),
    .A2(_03929_),
    .B1(_03946_),
    .B2(_03947_),
    .X(_03949_));
 sky130_fd_sc_hd__nand2_1 _12096_ (.A(_03948_),
    .B(_03949_),
    .Y(_03951_));
 sky130_fd_sc_hd__a31o_1 _12097_ (.A1(_03517_),
    .A2(_03528_),
    .A3(_03529_),
    .B1(_03518_),
    .X(_03952_));
 sky130_fd_sc_hd__nand2_1 _12098_ (.A(_03951_),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__or2_1 _12099_ (.A(_03952_),
    .B(_03951_),
    .X(_03954_));
 sky130_fd_sc_hd__or4_2 _12100_ (.A(_05381_),
    .B(_05403_),
    .C(_02049_),
    .D(_02051_),
    .X(_03955_));
 sky130_fd_sc_hd__or4_1 _12101_ (.A(_06331_),
    .B(net152),
    .C(_01589_),
    .D(_01822_),
    .X(_03956_));
 sky130_fd_sc_hd__o32a_1 _12102_ (.A1(net152),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(_06331_),
    .X(_03957_));
 sky130_fd_sc_hd__a31o_1 _12103_ (.A1(net151),
    .A2(_01823_),
    .A3(_03535_),
    .B1(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__xor2_1 _12104_ (.A(_03955_),
    .B(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__a21oi_1 _12105_ (.A1(_03953_),
    .A2(_03954_),
    .B1(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand3_1 _12106_ (.A(_03953_),
    .B(_03954_),
    .C(_03959_),
    .Y(_03962_));
 sky130_fd_sc_hd__and2b_1 _12107_ (.A_N(_03960_),
    .B(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__a21boi_1 _12108_ (.A1(_03532_),
    .A2(_03541_),
    .B1_N(_03534_),
    .Y(_03964_));
 sky130_fd_sc_hd__nor2_1 _12109_ (.A(_03963_),
    .B(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_1 _12110_ (.A(_03963_),
    .B(_03964_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand2b_1 _12111_ (.A_N(_03965_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__o21ai_1 _12112_ (.A1(_03546_),
    .A2(_03549_),
    .B1(_03547_),
    .Y(_03968_));
 sky130_fd_sc_hd__xor2_1 _12113_ (.A(_03967_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__and3_1 _12114_ (.A(_03432_),
    .B(_03508_),
    .C(_03510_),
    .X(_03970_));
 sky130_fd_sc_hd__a311o_1 _12115_ (.A1(_03432_),
    .A2(_03508_),
    .A3(_03510_),
    .B1(_03969_),
    .C1(_03509_),
    .X(_03971_));
 sky130_fd_sc_hd__o21ai_1 _12116_ (.A1(_03509_),
    .A2(_03970_),
    .B1(_03969_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand3b_1 _12117_ (.A_N(_03923_),
    .B(_03971_),
    .C(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__a21bo_1 _12118_ (.A1(_03971_),
    .A2(_03973_),
    .B1_N(_03923_),
    .X(_03975_));
 sky130_fd_sc_hd__a21oi_1 _12119_ (.A1(_03974_),
    .A2(_03975_),
    .B1(_03877_),
    .Y(_03976_));
 sky130_fd_sc_hd__nand3_2 _12120_ (.A(_03877_),
    .B(_03974_),
    .C(_03975_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand2b_1 _12121_ (.A_N(_03976_),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__a32o_1 _12122_ (.A1(_03505_),
    .A2(_03595_),
    .A3(_03596_),
    .B1(_03601_),
    .B2(_03597_),
    .X(_03979_));
 sky130_fd_sc_hd__xor2_1 _12123_ (.A(_03978_),
    .B(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__o21ba_1 _12124_ (.A1(_03871_),
    .A2(_03874_),
    .B1_N(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__xnor2_2 _12125_ (.A(_03876_),
    .B(_03980_),
    .Y(_03982_));
 sky130_fd_sc_hd__inv_2 _12126_ (.A(_03982_),
    .Y(_03984_));
 sky130_fd_sc_hd__or2_1 _12127_ (.A(_03751_),
    .B(_03982_),
    .X(_03985_));
 sky130_fd_sc_hd__nand2_1 _12128_ (.A(_03982_),
    .B(_03751_),
    .Y(_03986_));
 sky130_fd_sc_hd__nand2_1 _12129_ (.A(_03985_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__xor2_1 _12130_ (.A(_03759_),
    .B(_03987_),
    .X(_03988_));
 sky130_fd_sc_hd__a21oi_1 _12131_ (.A1(_00845_),
    .A2(_03761_),
    .B1(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__and3_1 _12132_ (.A(_00845_),
    .B(_03761_),
    .C(_03988_),
    .X(_03990_));
 sky130_fd_sc_hd__or2_1 _12133_ (.A(_03989_),
    .B(_03990_),
    .X(net89));
 sky130_fd_sc_hd__a31o_1 _12134_ (.A1(_03502_),
    .A2(_03760_),
    .A3(_03988_),
    .B1(_00834_),
    .X(_03991_));
 sky130_fd_sc_hd__or3_2 _12135_ (.A(_05327_),
    .B(_02092_),
    .C(_02094_),
    .X(_03992_));
 sky130_fd_sc_hd__a21bo_1 _12136_ (.A1(_03812_),
    .A2(_03846_),
    .B1_N(_03848_),
    .X(_03994_));
 sky130_fd_sc_hd__nand3_1 _12137_ (.A(_03816_),
    .B(_03841_),
    .C(_03842_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_1 _12138_ (.A(_03817_),
    .B(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__and3_1 _12139_ (.A(_02647_),
    .B(_02922_),
    .C(_02924_),
    .X(_03997_));
 sky130_fd_sc_hd__nand2_2 _12140_ (.A(_03820_),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__a32o_1 _12141_ (.A1(_02647_),
    .A2(_02922_),
    .A3(_02924_),
    .B1(_03087_),
    .B2(_01969_),
    .X(_03999_));
 sky130_fd_sc_hd__o31a_1 _12142_ (.A1(_02636_),
    .A2(_03086_),
    .A3(_03821_),
    .B1(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__nand2_1 _12143_ (.A(_03998_),
    .B(_03999_),
    .Y(_04001_));
 sky130_fd_sc_hd__and3_2 _12144_ (.A(_03831_),
    .B(_00976_),
    .C(_00965_),
    .X(_04002_));
 sky130_fd_sc_hd__a21oi_1 _12145_ (.A1(_03312_),
    .A2(_03315_),
    .B1(_01488_),
    .Y(_04003_));
 sky130_fd_sc_hd__o21ai_2 _12146_ (.A1(net54),
    .A2(_03313_),
    .B1(_04003_),
    .Y(_04005_));
 sky130_fd_sc_hd__a32o_1 _12147_ (.A1(net164),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_04003_),
    .B2(_03318_),
    .X(_04006_));
 sky130_fd_sc_hd__o2111a_1 _12148_ (.A1(net54),
    .A2(_03313_),
    .B1(_03650_),
    .C1(_04003_),
    .D1(_03651_),
    .X(_04007_));
 sky130_fd_sc_hd__nand3b_1 _12149_ (.A_N(_04005_),
    .B(_03653_),
    .C(net164),
    .Y(_04008_));
 sky130_fd_sc_hd__a22oi_2 _12150_ (.A1(_03826_),
    .A2(_04005_),
    .B1(_04007_),
    .B2(net164),
    .Y(_04009_));
 sky130_fd_sc_hd__nand2_1 _12151_ (.A(_04006_),
    .B(_04008_),
    .Y(_04010_));
 sky130_fd_sc_hd__o211a_1 _12152_ (.A1(_03834_),
    .A2(_00987_),
    .B1(_04010_),
    .C1(_04001_),
    .X(_04011_));
 sky130_fd_sc_hd__o211ai_2 _12153_ (.A1(_03834_),
    .A2(_00987_),
    .B1(_04010_),
    .C1(_04001_),
    .Y(_04012_));
 sky130_fd_sc_hd__o21ai_4 _12154_ (.A1(_04002_),
    .A2(_04009_),
    .B1(_04000_),
    .Y(_04013_));
 sky130_fd_sc_hd__o311a_1 _12155_ (.A1(net166),
    .A2(_03319_),
    .A3(_03659_),
    .B1(_04012_),
    .C1(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__a21oi_2 _12156_ (.A1(_04012_),
    .A2(_04013_),
    .B1(_03827_),
    .Y(_04016_));
 sky130_fd_sc_hd__a21o_1 _12157_ (.A1(_04012_),
    .A2(_04013_),
    .B1(_03827_),
    .X(_04017_));
 sky130_fd_sc_hd__o41a_1 _12158_ (.A1(_02636_),
    .A2(_03906_),
    .A3(_02433_),
    .A4(_02696_),
    .B1(_03809_),
    .X(_04018_));
 sky130_fd_sc_hd__nor2_1 _12159_ (.A(_03810_),
    .B(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__o21ai_1 _12160_ (.A1(_03823_),
    .A2(_03835_),
    .B1(_03661_),
    .Y(_04020_));
 sky130_fd_sc_hd__and4b_1 _12161_ (.A_N(_03321_),
    .B(_03653_),
    .C(_03839_),
    .D(_00998_),
    .X(_04021_));
 sky130_fd_sc_hd__o22ai_2 _12162_ (.A1(_03810_),
    .A2(_04018_),
    .B1(_03823_),
    .B2(_03835_),
    .Y(_04022_));
 sky130_fd_sc_hd__a21o_1 _12163_ (.A1(_03839_),
    .A2(_03660_),
    .B1(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__and3_1 _12164_ (.A(_03839_),
    .B(_04019_),
    .C(_04020_),
    .X(_04024_));
 sky130_fd_sc_hd__nand3_2 _12165_ (.A(_03839_),
    .B(_04019_),
    .C(_04020_),
    .Y(_04025_));
 sky130_fd_sc_hd__nand2_1 _12166_ (.A(_04023_),
    .B(_04025_),
    .Y(_04027_));
 sky130_fd_sc_hd__nand4b_1 _12167_ (.A_N(_04014_),
    .B(_04017_),
    .C(_04023_),
    .D(_04025_),
    .Y(_04028_));
 sky130_fd_sc_hd__o21ai_1 _12168_ (.A1(_04014_),
    .A2(_04016_),
    .B1(_04027_),
    .Y(_04029_));
 sky130_fd_sc_hd__o221ai_2 _12169_ (.A1(_04014_),
    .A2(_04016_),
    .B1(_04022_),
    .B2(_04021_),
    .C1(_04025_),
    .Y(_04030_));
 sky130_fd_sc_hd__a211o_1 _12170_ (.A1(_04023_),
    .A2(_04025_),
    .B1(_04014_),
    .C1(_04016_),
    .X(_04031_));
 sky130_fd_sc_hd__nand3_1 _12171_ (.A(_04031_),
    .B(_03996_),
    .C(_04030_),
    .Y(_04032_));
 sky130_fd_sc_hd__nand4_1 _12172_ (.A(_03817_),
    .B(_03995_),
    .C(_04028_),
    .D(_04029_),
    .Y(_04033_));
 sky130_fd_sc_hd__and3_1 _12173_ (.A(_04255_),
    .B(_02427_),
    .C(_02428_),
    .X(_04034_));
 sky130_fd_sc_hd__and4_1 _12174_ (.A(_03639_),
    .B(_03820_),
    .C(_03917_),
    .D(_02697_),
    .X(_04035_));
 sky130_fd_sc_hd__a32o_1 _12175_ (.A1(_03820_),
    .A2(_02926_),
    .A3(_01499_),
    .B1(_02697_),
    .B2(_03917_),
    .X(_04036_));
 sky130_fd_sc_hd__nand2b_1 _12176_ (.A_N(_04035_),
    .B(_04036_),
    .Y(_04038_));
 sky130_fd_sc_hd__xnor2_1 _12177_ (.A(_04034_),
    .B(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__a21o_1 _12178_ (.A1(_04032_),
    .A2(_04033_),
    .B1(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__nand3_1 _12179_ (.A(_04032_),
    .B(_04033_),
    .C(_04039_),
    .Y(_04041_));
 sky130_fd_sc_hd__nand3_1 _12180_ (.A(_03994_),
    .B(_04040_),
    .C(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__inv_2 _12181_ (.A(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__a21o_1 _12182_ (.A1(_04040_),
    .A2(_04041_),
    .B1(_03994_),
    .X(_04044_));
 sky130_fd_sc_hd__nand2_1 _12183_ (.A(_04042_),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand3b_2 _12184_ (.A_N(_03681_),
    .B(_03683_),
    .C(_03852_),
    .Y(_04046_));
 sky130_fd_sc_hd__and3_1 _12185_ (.A(_03853_),
    .B(_04045_),
    .C(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__a21oi_1 _12186_ (.A1(_03853_),
    .A2(_04046_),
    .B1(_04045_),
    .Y(_04049_));
 sky130_fd_sc_hd__nor2_1 _12187_ (.A(_04047_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__or4_2 _12188_ (.A(_05327_),
    .B(_02092_),
    .C(_02094_),
    .D(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__o31a_2 _12189_ (.A1(_05327_),
    .A2(_02092_),
    .A3(_02094_),
    .B1(_04050_),
    .X(_04052_));
 sky130_fd_sc_hd__xnor2_1 _12190_ (.A(_03992_),
    .B(_04050_),
    .Y(_04053_));
 sky130_fd_sc_hd__a31oi_4 _12191_ (.A1(_03789_),
    .A2(_03795_),
    .A3(_03797_),
    .B1(_03790_),
    .Y(_04054_));
 sky130_fd_sc_hd__o31ai_1 _12192_ (.A1(_00532_),
    .A2(_00580_),
    .A3(_03792_),
    .B1(_03794_),
    .Y(_04055_));
 sky130_fd_sc_hd__o21ai_1 _12193_ (.A1(_03286_),
    .A2(_03704_),
    .B1(_03781_),
    .Y(_04056_));
 sky130_fd_sc_hd__a21o_1 _12194_ (.A1(_03780_),
    .A2(_04056_),
    .B1(_04055_),
    .X(_04057_));
 sky130_fd_sc_hd__nand3_1 _12195_ (.A(_03780_),
    .B(_04055_),
    .C(_04056_),
    .Y(_04058_));
 sky130_fd_sc_hd__and3_1 _12196_ (.A(_00193_),
    .B(_01185_),
    .C(_01187_),
    .X(_04060_));
 sky130_fd_sc_hd__o32a_1 _12197_ (.A1(_00192_),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_01272_),
    .B2(net148),
    .X(_04061_));
 sky130_fd_sc_hd__and3_1 _12198_ (.A(_04060_),
    .B(_01273_),
    .C(_00072_),
    .X(_04062_));
 sky130_fd_sc_hd__or4_1 _12199_ (.A(net148),
    .B(_00192_),
    .C(_01188_),
    .D(_01272_),
    .X(_04063_));
 sky130_fd_sc_hd__nor2_1 _12200_ (.A(_04061_),
    .B(_04062_),
    .Y(_04064_));
 sky130_fd_sc_hd__o21ai_2 _12201_ (.A1(_07441_),
    .A2(_01662_),
    .B1(_03773_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand4_2 _12202_ (.A(net162),
    .B(_07437_),
    .C(_01879_),
    .D(net134),
    .Y(_04066_));
 sky130_fd_sc_hd__o21ai_1 _12203_ (.A1(_03704_),
    .A2(_04066_),
    .B1(_04065_),
    .Y(_04067_));
 sky130_fd_sc_hd__o21ai_1 _12204_ (.A1(net149),
    .A2(_01542_),
    .B1(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__o2111ai_1 _12205_ (.A1(_03704_),
    .A2(_04066_),
    .B1(_04065_),
    .C1(_07540_),
    .D1(_01544_),
    .Y(_04069_));
 sky130_fd_sc_hd__a2bb2o_1 _12206_ (.A1_N(_04061_),
    .A2_N(_04062_),
    .B1(_04068_),
    .B2(_04069_),
    .X(_04071_));
 sky130_fd_sc_hd__nand3_1 _12207_ (.A(_04068_),
    .B(_04069_),
    .C(_04064_),
    .Y(_04072_));
 sky130_fd_sc_hd__a32o_1 _12208_ (.A1(_03701_),
    .A2(_01883_),
    .A3(_07200_),
    .B1(_03772_),
    .B2(_03770_),
    .X(_04073_));
 sky130_fd_sc_hd__a21o_1 _12209_ (.A1(_04071_),
    .A2(_04072_),
    .B1(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__nand3_1 _12210_ (.A(_04071_),
    .B(_04072_),
    .C(_04073_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_1 _12211_ (.A(_04074_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__a22o_1 _12212_ (.A1(_04057_),
    .A2(_04058_),
    .B1(_04074_),
    .B2(_04075_),
    .X(_04077_));
 sky130_fd_sc_hd__nand4_1 _12213_ (.A(_04057_),
    .B(_04058_),
    .C(_04074_),
    .D(_04075_),
    .Y(_04078_));
 sky130_fd_sc_hd__nand2_1 _12214_ (.A(_04077_),
    .B(_04078_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand3_1 _12215_ (.A(_03765_),
    .B(_03782_),
    .C(_03783_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21oi_1 _12216_ (.A1(_03766_),
    .A2(_04080_),
    .B1(_04079_),
    .Y(_04082_));
 sky130_fd_sc_hd__a21o_1 _12217_ (.A1(_03766_),
    .A2(_04080_),
    .B1(_04079_),
    .X(_04083_));
 sky130_fd_sc_hd__nand3_1 _12218_ (.A(_03766_),
    .B(_04079_),
    .C(_04080_),
    .Y(_04084_));
 sky130_fd_sc_hd__and3_1 _12219_ (.A(_03768_),
    .B(_00364_),
    .C(_00362_),
    .X(_04085_));
 sky130_fd_sc_hd__or4_1 _12220_ (.A(_00361_),
    .B(_00363_),
    .C(_01037_),
    .D(_03769_),
    .X(_04086_));
 sky130_fd_sc_hd__a31o_1 _12221_ (.A1(_00362_),
    .A2(_00364_),
    .A3(_01038_),
    .B1(_03768_),
    .X(_04087_));
 sky130_fd_sc_hd__o211ai_1 _12222_ (.A1(_00744_),
    .A2(_00532_),
    .B1(_04087_),
    .C1(_04086_),
    .Y(_04088_));
 sky130_fd_sc_hd__a221o_1 _12223_ (.A1(_00741_),
    .A2(_00742_),
    .B1(_04086_),
    .B2(_04087_),
    .C1(_00532_),
    .X(_04089_));
 sky130_fd_sc_hd__nand2_1 _12224_ (.A(_04088_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__nand3_1 _12225_ (.A(_04083_),
    .B(_04084_),
    .C(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a21o_1 _12226_ (.A1(_04083_),
    .A2(_04084_),
    .B1(_04090_),
    .X(_04093_));
 sky130_fd_sc_hd__nand2_1 _12227_ (.A(_04091_),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_1 _12228_ (.A(_04094_),
    .B(_04054_),
    .Y(_04095_));
 sky130_fd_sc_hd__nor2_1 _12229_ (.A(_04054_),
    .B(_04094_),
    .Y(_04096_));
 sky130_fd_sc_hd__xnor2_2 _12230_ (.A(_04054_),
    .B(_04094_),
    .Y(_04097_));
 sky130_fd_sc_hd__a21oi_4 _12231_ (.A1(_03804_),
    .A2(_03806_),
    .B1(_03803_),
    .Y(_04098_));
 sky130_fd_sc_hd__xor2_4 _12232_ (.A(_04097_),
    .B(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__xnor2_1 _12233_ (.A(_04053_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__or2_2 _12234_ (.A(_03864_),
    .B(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__nand2_1 _12235_ (.A(_03864_),
    .B(_04100_),
    .Y(_04102_));
 sky130_fd_sc_hd__o211ai_2 _12236_ (.A1(_03382_),
    .A2(_03732_),
    .B1(_03867_),
    .C1(_03869_),
    .Y(_04104_));
 sky130_fd_sc_hd__o21bai_1 _12237_ (.A1(_03865_),
    .A2(_03866_),
    .B1_N(_03870_),
    .Y(_04105_));
 sky130_fd_sc_hd__a22o_1 _12238_ (.A1(_04101_),
    .A2(_04102_),
    .B1(_04105_),
    .B2(_03867_),
    .X(_04106_));
 sky130_fd_sc_hd__nand4_1 _12239_ (.A(_03867_),
    .B(_04101_),
    .C(_04102_),
    .D(_04105_),
    .Y(_04107_));
 sky130_fd_sc_hd__and2_2 _12240_ (.A(_04106_),
    .B(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__o21ai_4 _12241_ (.A1(_00570_),
    .A2(_00580_),
    .B1(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__or4_2 _12242_ (.A(_00570_),
    .B(_00576_),
    .C(_00578_),
    .D(_04108_),
    .X(_04110_));
 sky130_fd_sc_hd__a21oi_1 _12243_ (.A1(_03922_),
    .A2(_03920_),
    .B1(_03919_),
    .Y(_04111_));
 sky130_fd_sc_hd__a31o_1 _12244_ (.A1(_03879_),
    .A2(_03904_),
    .A3(_03905_),
    .B1(_03914_),
    .X(_04112_));
 sky130_fd_sc_hd__o32a_1 _12245_ (.A1(_02122_),
    .A2(_03558_),
    .A3(_03179_),
    .B1(_01292_),
    .B2(_03583_),
    .X(_04113_));
 sky130_fd_sc_hd__and4bb_1 _12246_ (.A_N(_03558_),
    .B_N(_03887_),
    .C(_03584_),
    .D(_01303_),
    .X(_04115_));
 sky130_fd_sc_hd__a2bb2o_1 _12247_ (.A1_N(_04113_),
    .A2_N(_04115_),
    .B1(_00911_),
    .B2(_03911_),
    .X(_04116_));
 sky130_fd_sc_hd__o22a_1 _12248_ (.A1(_03882_),
    .A2(_03881_),
    .B1(_03902_),
    .B2(_03900_),
    .X(_04117_));
 sky130_fd_sc_hd__a21oi_1 _12249_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(_03899_),
    .B(_03561_),
    .Y(_04119_));
 sky130_fd_sc_hd__a21oi_1 _12251_ (.A1(_03898_),
    .A2(_04119_),
    .B1(_03909_),
    .Y(_04120_));
 sky130_fd_sc_hd__inv_2 _12252_ (.A(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__and3_1 _12253_ (.A(_03898_),
    .B(_03909_),
    .C(_04119_),
    .X(_04122_));
 sky130_fd_sc_hd__nand3_1 _12254_ (.A(_03898_),
    .B(_03909_),
    .C(_04119_),
    .Y(_04123_));
 sky130_fd_sc_hd__or4_1 _12255_ (.A(_02210_),
    .B(_03175_),
    .C(_03177_),
    .D(_03449_),
    .X(_04124_));
 sky130_fd_sc_hd__o22ai_2 _12256_ (.A1(_02122_),
    .A2(_03179_),
    .B1(_03449_),
    .B2(_01620_),
    .Y(_04126_));
 sky130_fd_sc_hd__o31ai_4 _12257_ (.A1(_02210_),
    .A2(_03179_),
    .A3(_03449_),
    .B1(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__and3_1 _12258_ (.A(_02866_),
    .B(_02854_),
    .C(_02856_),
    .X(_04128_));
 sky130_fd_sc_hd__o2111ai_4 _12259_ (.A1(_04606_),
    .A2(_04660_),
    .B1(_04704_),
    .C1(_02629_),
    .D1(_02631_),
    .Y(_04129_));
 sky130_fd_sc_hd__o22ai_4 _12260_ (.A1(net155),
    .A2(_02355_),
    .B1(_02632_),
    .B2(net158),
    .Y(_04130_));
 sky130_fd_sc_hd__o21ai_1 _12261_ (.A1(_03560_),
    .A2(_04129_),
    .B1(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _12262_ (.A(_04131_),
    .B(_04128_),
    .Y(_04132_));
 sky130_fd_sc_hd__o221ai_4 _12263_ (.A1(net159),
    .A2(_02857_),
    .B1(_03560_),
    .B2(_04129_),
    .C1(_04130_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand3_1 _12264_ (.A(_04127_),
    .B(_04132_),
    .C(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__a21o_1 _12265_ (.A1(_04132_),
    .A2(_04133_),
    .B1(_04127_),
    .X(_04135_));
 sky130_fd_sc_hd__o2bb2a_1 _12266_ (.A1_N(_03889_),
    .A2_N(_03890_),
    .B1(_03891_),
    .B2(_02355_),
    .X(_04137_));
 sky130_fd_sc_hd__nand3_1 _12267_ (.A(_04134_),
    .B(_04135_),
    .C(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__a21o_1 _12268_ (.A1(_04134_),
    .A2(_04135_),
    .B1(_04137_),
    .X(_04139_));
 sky130_fd_sc_hd__a22o_1 _12269_ (.A1(_04121_),
    .A2(_04123_),
    .B1(_04138_),
    .B2(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__nand4_1 _12270_ (.A(_04121_),
    .B(_04123_),
    .C(_04138_),
    .D(_04139_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand3_1 _12271_ (.A(_04118_),
    .B(_04140_),
    .C(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__a21o_1 _12272_ (.A1(_04140_),
    .A2(_04141_),
    .B1(_04118_),
    .X(_04143_));
 sky130_fd_sc_hd__a21oi_1 _12273_ (.A1(_04142_),
    .A2(_04143_),
    .B1(_04116_),
    .Y(_04144_));
 sky130_fd_sc_hd__a21boi_1 _12274_ (.A1(_04116_),
    .A2(_04142_),
    .B1_N(_04143_),
    .Y(_04145_));
 sky130_fd_sc_hd__a31o_1 _12275_ (.A1(_04116_),
    .A2(_04142_),
    .A3(_04143_),
    .B1(_04144_),
    .X(_04146_));
 sky130_fd_sc_hd__a21oi_1 _12276_ (.A1(_03907_),
    .A2(_04112_),
    .B1(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand3_1 _12277_ (.A(_03907_),
    .B(_04112_),
    .C(_04146_),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2b_1 _12278_ (.A_N(_04147_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__a21o_1 _12279_ (.A1(_04111_),
    .A2(_04148_),
    .B1(_04147_),
    .X(_04150_));
 sky130_fd_sc_hd__xnor2_1 _12280_ (.A(_04111_),
    .B(_04149_),
    .Y(_04151_));
 sky130_fd_sc_hd__and3_1 _12281_ (.A(_05436_),
    .B(net139),
    .C(_02237_),
    .X(_04152_));
 sky130_fd_sc_hd__o21ai_1 _12282_ (.A1(_03957_),
    .A2(_03955_),
    .B1(_03956_),
    .Y(_04153_));
 sky130_fd_sc_hd__o21ai_1 _12283_ (.A1(_03396_),
    .A2(_03520_),
    .B1(_03945_),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _12284_ (.A(_03944_),
    .B(_03524_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand3_2 _12285_ (.A(_04153_),
    .B(_04154_),
    .C(_03944_),
    .Y(_04156_));
 sky130_fd_sc_hd__o2111a_1 _12286_ (.A1(_03957_),
    .A2(_03955_),
    .B1(_03945_),
    .C1(_03956_),
    .D1(_04155_),
    .X(_04158_));
 sky130_fd_sc_hd__a21o_1 _12287_ (.A1(_03944_),
    .A2(_04154_),
    .B1(_04153_),
    .X(_04159_));
 sky130_fd_sc_hd__a32o_1 _12288_ (.A1(_07513_),
    .A2(_01585_),
    .A3(_01588_),
    .B1(_01405_),
    .B2(_00010_),
    .X(_04160_));
 sky130_fd_sc_hd__and4_1 _12289_ (.A(_01405_),
    .B(_01590_),
    .C(_07513_),
    .D(_00010_),
    .X(_04161_));
 sky130_fd_sc_hd__nand4_2 _12290_ (.A(_01405_),
    .B(_01590_),
    .C(_07513_),
    .D(_00010_),
    .Y(_04162_));
 sky130_fd_sc_hd__and3_1 _12291_ (.A(_00150_),
    .B(net145),
    .C(_01220_),
    .X(_04163_));
 sky130_fd_sc_hd__o2111ai_4 _12292_ (.A1(_00299_),
    .A2(_00424_),
    .B1(_00427_),
    .C1(_01055_),
    .D1(_01057_),
    .Y(_04164_));
 sky130_fd_sc_hd__nor2_1 _12293_ (.A(_03523_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__o21ai_2 _12294_ (.A1(_00274_),
    .A2(_01058_),
    .B1(_03936_),
    .Y(_04166_));
 sky130_fd_sc_hd__o21ai_1 _12295_ (.A1(_03523_),
    .A2(_04164_),
    .B1(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__o21ai_1 _12296_ (.A1(net144),
    .A2(_01221_),
    .B1(_04167_),
    .Y(_04169_));
 sky130_fd_sc_hd__o2111ai_2 _12297_ (.A1(_03523_),
    .A2(_04164_),
    .B1(_04166_),
    .C1(_01222_),
    .D1(_00150_),
    .Y(_04170_));
 sky130_fd_sc_hd__a22o_1 _12298_ (.A1(_04160_),
    .A2(_04162_),
    .B1(_04169_),
    .B2(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__nand4_2 _12299_ (.A(_04160_),
    .B(_04162_),
    .C(_04169_),
    .D(_04170_),
    .Y(_04172_));
 sky130_fd_sc_hd__o31ai_1 _12300_ (.A1(net144),
    .A2(_01058_),
    .A3(_03934_),
    .B1(_03937_),
    .Y(_04173_));
 sky130_fd_sc_hd__a21o_1 _12301_ (.A1(_04171_),
    .A2(_04172_),
    .B1(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__nand3_1 _12302_ (.A(_04171_),
    .B(_04172_),
    .C(_04173_),
    .Y(_04175_));
 sky130_fd_sc_hd__nand2_1 _12303_ (.A(_04174_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__a22o_1 _12304_ (.A1(_04156_),
    .A2(_04159_),
    .B1(_04174_),
    .B2(_04175_),
    .X(_04177_));
 sky130_fd_sc_hd__nand4_1 _12305_ (.A(_04156_),
    .B(_04159_),
    .C(_04174_),
    .D(_04175_),
    .Y(_04178_));
 sky130_fd_sc_hd__a21bo_1 _12306_ (.A1(_03946_),
    .A2(_03947_),
    .B1_N(_03929_),
    .X(_04180_));
 sky130_fd_sc_hd__a22o_1 _12307_ (.A1(_04177_),
    .A2(_04178_),
    .B1(_04180_),
    .B2(_03927_),
    .X(_04181_));
 sky130_fd_sc_hd__nand4_1 _12308_ (.A(_03927_),
    .B(_04177_),
    .C(_04178_),
    .D(_04180_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2_1 _12309_ (.A(_04181_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__or3_1 _12310_ (.A(_06331_),
    .B(_02049_),
    .C(_02051_),
    .X(_04184_));
 sky130_fd_sc_hd__o32a_1 _12311_ (.A1(_00009_),
    .A2(_01406_),
    .A3(_03519_),
    .B1(_01822_),
    .B2(net152),
    .X(_04185_));
 sky130_fd_sc_hd__or4_1 _12312_ (.A(net152),
    .B(_03519_),
    .C(_03931_),
    .D(_01822_),
    .X(_04186_));
 sky130_fd_sc_hd__nand2b_1 _12313_ (.A_N(_04185_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__xnor2_1 _12314_ (.A(_04184_),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__and2_1 _12315_ (.A(_04183_),
    .B(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__nor2_1 _12316_ (.A(_04183_),
    .B(_04188_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_1 _12317_ (.A(_04182_),
    .B(_04188_),
    .Y(_04192_));
 sky130_fd_sc_hd__a21boi_1 _12318_ (.A1(_03953_),
    .A2(_03959_),
    .B1_N(_03954_),
    .Y(_04193_));
 sky130_fd_sc_hd__nor3_1 _12319_ (.A(_04193_),
    .B(_04191_),
    .C(_04189_),
    .Y(_04194_));
 sky130_fd_sc_hd__o21ai_1 _12320_ (.A1(_04189_),
    .A2(_04191_),
    .B1(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2b_1 _12321_ (.A_N(_04194_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__a21oi_2 _12322_ (.A1(_03968_),
    .A2(_03966_),
    .B1(_03965_),
    .Y(_04197_));
 sky130_fd_sc_hd__xnor2_1 _12323_ (.A(_04196_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__xnor2_1 _12324_ (.A(_04152_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__a31o_1 _12325_ (.A1(_05436_),
    .A2(_02240_),
    .A3(_04198_),
    .B1(_04151_),
    .X(_04200_));
 sky130_fd_sc_hd__o21ai_1 _12326_ (.A1(_04152_),
    .A2(_04198_),
    .B1(_04200_),
    .Y(_04202_));
 sky130_fd_sc_hd__xnor2_1 _12327_ (.A(_04151_),
    .B(_04199_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21bo_1 _12328_ (.A1(_03971_),
    .A2(_03923_),
    .B1_N(_03973_),
    .X(_04204_));
 sky130_fd_sc_hd__nor2_1 _12329_ (.A(_04204_),
    .B(_04203_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand2_1 _12330_ (.A(_04203_),
    .B(_04204_),
    .Y(_04206_));
 sky130_fd_sc_hd__and2b_1 _12331_ (.A_N(_04205_),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__a31oi_4 _12332_ (.A1(_03597_),
    .A2(_03603_),
    .A3(_03977_),
    .B1(_03976_),
    .Y(_04208_));
 sky130_fd_sc_hd__xnor2_2 _12333_ (.A(_04207_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__a21o_1 _12334_ (.A1(_04109_),
    .A2(_04110_),
    .B1(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__nand3_1 _12335_ (.A(_04109_),
    .B(_04110_),
    .C(_04209_),
    .Y(_04211_));
 sky130_fd_sc_hd__a221o_1 _12336_ (.A1(_03871_),
    .A2(_03874_),
    .B1(_04210_),
    .B2(_04211_),
    .C1(_03981_),
    .X(_04213_));
 sky130_fd_sc_hd__o211ai_4 _12337_ (.A1(_03875_),
    .A2(_03981_),
    .B1(_04210_),
    .C1(_04211_),
    .Y(_04214_));
 sky130_fd_sc_hd__o211ai_4 _12338_ (.A1(_03982_),
    .A2(_03751_),
    .B1(_03757_),
    .C1(_03758_),
    .Y(_04215_));
 sky130_fd_sc_hd__a22o_1 _12339_ (.A1(_04213_),
    .A2(_04214_),
    .B1(_04215_),
    .B2(_03986_),
    .X(_04216_));
 sky130_fd_sc_hd__o2111ai_1 _12340_ (.A1(_03750_),
    .A2(_03984_),
    .B1(_04213_),
    .C1(_04214_),
    .D1(_04215_),
    .Y(_04217_));
 sky130_fd_sc_hd__and2_1 _12341_ (.A(_04216_),
    .B(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__xnor2_1 _12342_ (.A(_03991_),
    .B(_04218_),
    .Y(net90));
 sky130_fd_sc_hd__and4b_2 _12343_ (.A_N(_04218_),
    .B(_03988_),
    .C(_03760_),
    .D(_03502_),
    .X(_04219_));
 sky130_fd_sc_hd__o211ai_4 _12344_ (.A1(_03750_),
    .A2(_03984_),
    .B1(_04213_),
    .C1(_04215_),
    .Y(_04220_));
 sky130_fd_sc_hd__a21boi_4 _12345_ (.A1(_04109_),
    .A2(_04209_),
    .B1_N(_04110_),
    .Y(_04221_));
 sky130_fd_sc_hd__inv_2 _12346_ (.A(_04221_),
    .Y(_04223_));
 sky130_fd_sc_hd__and4_1 _12347_ (.A(_01631_),
    .B(_02133_),
    .C(_03450_),
    .D(_03584_),
    .X(_04224_));
 sky130_fd_sc_hd__o32a_1 _12348_ (.A1(_01620_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(_02122_),
    .B2(_03449_),
    .X(_04225_));
 sky130_fd_sc_hd__o22a_1 _12349_ (.A1(_03912_),
    .A2(_01292_),
    .B1(_04225_),
    .B2(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__a31o_1 _12350_ (.A1(_04121_),
    .A2(_04138_),
    .A3(_04139_),
    .B1(_04122_),
    .X(_04227_));
 sky130_fd_sc_hd__a32oi_4 _12351_ (.A1(_04127_),
    .A2(_04132_),
    .A3(_04133_),
    .B1(_04135_),
    .B2(_04137_),
    .Y(_04228_));
 sky130_fd_sc_hd__xor2_1 _12352_ (.A(_04115_),
    .B(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__a41o_1 _12353_ (.A1(net156),
    .A2(_04726_),
    .A3(_02356_),
    .A4(_02633_),
    .B1(_04128_),
    .X(_04230_));
 sky130_fd_sc_hd__a32o_1 _12354_ (.A1(_04726_),
    .A2(_02629_),
    .A3(_02631_),
    .B1(_02858_),
    .B2(net156),
    .X(_04231_));
 sky130_fd_sc_hd__or3_1 _12355_ (.A(net158),
    .B(_02857_),
    .C(_04129_),
    .X(_04232_));
 sky130_fd_sc_hd__a32o_1 _12356_ (.A1(_02866_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_04231_),
    .B2(_04232_),
    .X(_04234_));
 sky130_fd_sc_hd__nand4_1 _12357_ (.A(_02866_),
    .B(_03180_),
    .C(_04231_),
    .D(_04232_),
    .Y(_04235_));
 sky130_fd_sc_hd__a22o_1 _12358_ (.A1(_04130_),
    .A2(_04230_),
    .B1(_04234_),
    .B2(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__nand4_2 _12359_ (.A(_04130_),
    .B(_04230_),
    .C(_04234_),
    .D(_04235_),
    .Y(_04237_));
 sky130_fd_sc_hd__a21o_1 _12360_ (.A1(_04236_),
    .A2(_04237_),
    .B1(_04124_),
    .X(_04238_));
 sky130_fd_sc_hd__nand3_1 _12361_ (.A(_04124_),
    .B(_04236_),
    .C(_04237_),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_1 _12362_ (.A(_04238_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__xnor2_2 _12363_ (.A(_04229_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__a311o_1 _12364_ (.A1(_04121_),
    .A2(_04138_),
    .A3(_04139_),
    .B1(_04241_),
    .C1(_04122_),
    .X(_04242_));
 sky130_fd_sc_hd__a21o_1 _12365_ (.A1(_04227_),
    .A2(_04241_),
    .B1(_04226_),
    .X(_04243_));
 sky130_fd_sc_hd__and3_1 _12366_ (.A(_04226_),
    .B(_04227_),
    .C(_04241_),
    .X(_04245_));
 sky130_fd_sc_hd__o21ai_1 _12367_ (.A1(_04227_),
    .A2(_04241_),
    .B1(_04243_),
    .Y(_04246_));
 sky130_fd_sc_hd__o22a_1 _12368_ (.A1(_04226_),
    .A2(_04242_),
    .B1(_04245_),
    .B2(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__nand2_1 _12369_ (.A(_04145_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__nor2_1 _12370_ (.A(_04145_),
    .B(_04247_),
    .Y(_04249_));
 sky130_fd_sc_hd__xnor2_1 _12371_ (.A(_04145_),
    .B(_04247_),
    .Y(_04250_));
 sky130_fd_sc_hd__xnor2_1 _12372_ (.A(_04150_),
    .B(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__and3_1 _12373_ (.A(_04152_),
    .B(_02356_),
    .C(_06341_),
    .X(_04252_));
 sky130_fd_sc_hd__or4_1 _12374_ (.A(_05425_),
    .B(_06331_),
    .C(_02241_),
    .D(_02355_),
    .X(_04253_));
 sky130_fd_sc_hd__o32a_1 _12375_ (.A1(_05425_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_06331_),
    .B2(_02241_),
    .X(_04254_));
 sky130_fd_sc_hd__a21o_1 _12376_ (.A1(_04195_),
    .A2(_04197_),
    .B1(_04194_),
    .X(_04256_));
 sky130_fd_sc_hd__a21oi_1 _12377_ (.A1(_04195_),
    .A2(_04197_),
    .B1(_04194_),
    .Y(_04257_));
 sky130_fd_sc_hd__or2_1 _12378_ (.A(_04158_),
    .B(_04176_),
    .X(_04258_));
 sky130_fd_sc_hd__o21ai_1 _12379_ (.A1(_04184_),
    .A2(_04185_),
    .B1(_04186_),
    .Y(_04259_));
 sky130_fd_sc_hd__o311ai_2 _12380_ (.A1(net144),
    .A2(_01058_),
    .A3(_03934_),
    .B1(_03937_),
    .C1(_04172_),
    .Y(_04260_));
 sky130_fd_sc_hd__nand3_1 _12381_ (.A(_04259_),
    .B(_04260_),
    .C(_04171_),
    .Y(_04261_));
 sky130_fd_sc_hd__a21o_1 _12382_ (.A1(_04171_),
    .A2(_04260_),
    .B1(_04259_),
    .X(_04262_));
 sky130_fd_sc_hd__nand2_1 _12383_ (.A(_04261_),
    .B(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__o21ai_1 _12384_ (.A1(_04163_),
    .A2(_04165_),
    .B1(_04166_),
    .Y(_04264_));
 sky130_fd_sc_hd__o31ai_2 _12385_ (.A1(_00274_),
    .A2(_01217_),
    .A3(_01219_),
    .B1(_04164_),
    .Y(_04265_));
 sky130_fd_sc_hd__a211o_1 _12386_ (.A1(_01214_),
    .A2(_01215_),
    .B1(_00274_),
    .C1(_04164_),
    .X(_04267_));
 sky130_fd_sc_hd__a31o_1 _12387_ (.A1(_00275_),
    .A2(net145),
    .A3(_01220_),
    .B1(_04164_),
    .X(_04268_));
 sky130_fd_sc_hd__o2111ai_4 _12388_ (.A1(net142),
    .A2(_01058_),
    .B1(net145),
    .C1(_01220_),
    .D1(_00275_),
    .Y(_04269_));
 sky130_fd_sc_hd__o211ai_2 _12389_ (.A1(_01406_),
    .A2(net144),
    .B1(_04269_),
    .C1(_04268_),
    .Y(_04270_));
 sky130_fd_sc_hd__nand4_1 _12390_ (.A(_00150_),
    .B(_04267_),
    .C(_01405_),
    .D(_04265_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand4_1 _12391_ (.A(_00150_),
    .B(_04268_),
    .C(_04269_),
    .D(_01405_),
    .Y(_04272_));
 sky130_fd_sc_hd__a22o_1 _12392_ (.A1(_00150_),
    .A2(_01405_),
    .B1(_04268_),
    .B2(_04269_),
    .X(_04273_));
 sky130_fd_sc_hd__nand3_1 _12393_ (.A(_04272_),
    .B(_04273_),
    .C(_04264_),
    .Y(_04274_));
 sky130_fd_sc_hd__o2111ai_4 _12394_ (.A1(_04163_),
    .A2(_04165_),
    .B1(_04166_),
    .C1(_04270_),
    .D1(_04271_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand3_1 _12395_ (.A(_04162_),
    .B(_04274_),
    .C(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__a21o_1 _12396_ (.A1(_04274_),
    .A2(_04275_),
    .B1(_04162_),
    .X(_04278_));
 sky130_fd_sc_hd__and2_1 _12397_ (.A(_04276_),
    .B(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__nor2_1 _12398_ (.A(_04263_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__and2_1 _12399_ (.A(_04263_),
    .B(_04279_),
    .X(_04281_));
 sky130_fd_sc_hd__o221a_1 _12400_ (.A1(_04158_),
    .A2(_04176_),
    .B1(_04280_),
    .B2(_04281_),
    .C1(_04156_),
    .X(_04282_));
 sky130_fd_sc_hd__o221ai_2 _12401_ (.A1(_04158_),
    .A2(_04176_),
    .B1(_04280_),
    .B2(_04281_),
    .C1(_04156_),
    .Y(_04283_));
 sky130_fd_sc_hd__a211oi_1 _12402_ (.A1(_04156_),
    .A2(_04258_),
    .B1(_04280_),
    .C1(_04281_),
    .Y(_04284_));
 sky130_fd_sc_hd__nor2_1 _12403_ (.A(_04282_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__a32o_1 _12404_ (.A1(_07513_),
    .A2(_01820_),
    .A3(_01821_),
    .B1(_00010_),
    .B2(_01590_),
    .X(_04286_));
 sky130_fd_sc_hd__or4_2 _12405_ (.A(_07512_),
    .B(_00009_),
    .C(_01589_),
    .D(_01822_),
    .X(_04287_));
 sky130_fd_sc_hd__a211o_1 _12406_ (.A1(_04286_),
    .A2(_04287_),
    .B1(net152),
    .C1(_02053_),
    .X(_04289_));
 sky130_fd_sc_hd__o211ai_1 _12407_ (.A1(net152),
    .A2(_02053_),
    .B1(_04286_),
    .C1(_04287_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _12408_ (.A(_04289_),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__xor2_1 _12409_ (.A(_04285_),
    .B(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__a21o_1 _12410_ (.A1(_04181_),
    .A2(_04192_),
    .B1(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__nand3_1 _12411_ (.A(_04292_),
    .B(_04192_),
    .C(_04181_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand4_1 _12412_ (.A(_04256_),
    .B(_04292_),
    .C(_04181_),
    .D(_04192_),
    .Y(_04295_));
 sky130_fd_sc_hd__a21boi_2 _12413_ (.A1(_04257_),
    .A2(_04294_),
    .B1_N(_04293_),
    .Y(_04296_));
 sky130_fd_sc_hd__o2bb2ai_1 _12414_ (.A1_N(_04295_),
    .A2_N(_04296_),
    .B1(_04256_),
    .B2(_04293_),
    .Y(_04297_));
 sky130_fd_sc_hd__o21ai_2 _12415_ (.A1(_04252_),
    .A2(_04254_),
    .B1(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__a311oi_2 _12416_ (.A1(_06341_),
    .A2(_02356_),
    .A3(_04152_),
    .B1(_04254_),
    .C1(_04297_),
    .Y(_04300_));
 sky130_fd_sc_hd__inv_2 _12417_ (.A(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21oi_1 _12418_ (.A1(_04298_),
    .A2(_04301_),
    .B1(_04251_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand3_1 _12419_ (.A(_04251_),
    .B(_04298_),
    .C(_04301_),
    .Y(_04303_));
 sky130_fd_sc_hd__nand2b_1 _12420_ (.A_N(_04302_),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__nand2_1 _12421_ (.A(_04202_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__nor2_1 _12422_ (.A(_04202_),
    .B(_04304_),
    .Y(_04306_));
 sky130_fd_sc_hd__or3b_1 _12423_ (.A(_04202_),
    .B(_04302_),
    .C_N(_04303_),
    .X(_04307_));
 sky130_fd_sc_hd__and2_1 _12424_ (.A(_04305_),
    .B(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__o21ai_4 _12425_ (.A1(_04205_),
    .A2(_04208_),
    .B1(_04206_),
    .Y(_04309_));
 sky130_fd_sc_hd__xnor2_4 _12426_ (.A(_04308_),
    .B(_04309_),
    .Y(_04311_));
 sky130_fd_sc_hd__and4_1 _12427_ (.A(_00569_),
    .B(_00743_),
    .C(_00904_),
    .D(_00581_),
    .X(_04312_));
 sky130_fd_sc_hd__o32a_1 _12428_ (.A1(_00576_),
    .A2(_00578_),
    .A3(_00903_),
    .B1(_00744_),
    .B2(_00570_),
    .X(_04313_));
 sky130_fd_sc_hd__o211ai_4 _12429_ (.A1(_03865_),
    .A2(_03866_),
    .B1(_04102_),
    .C1(_04104_),
    .Y(_04314_));
 sky130_fd_sc_hd__o21a_1 _12430_ (.A1(_03864_),
    .A2(_04100_),
    .B1(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__or4_1 _12431_ (.A(_05327_),
    .B(_07189_),
    .C(_02433_),
    .D(_02096_),
    .X(_04316_));
 sky130_fd_sc_hd__a32o_1 _12432_ (.A1(_05316_),
    .A2(_02427_),
    .A3(_02428_),
    .B1(_07200_),
    .B2(_02097_),
    .X(_04317_));
 sky130_fd_sc_hd__or3_1 _12433_ (.A(_04244_),
    .B(_02692_),
    .C(_02694_),
    .X(_04318_));
 sky130_fd_sc_hd__o32a_1 _12434_ (.A1(_02636_),
    .A2(net132),
    .A3(net130),
    .B1(_03906_),
    .B2(_02925_),
    .X(_04319_));
 sky130_fd_sc_hd__or4_1 _12435_ (.A(_02636_),
    .B(_03906_),
    .C(_02925_),
    .D(_03086_),
    .X(_04320_));
 sky130_fd_sc_hd__a31o_1 _12436_ (.A1(_03917_),
    .A2(_03087_),
    .A3(_03997_),
    .B1(_04319_),
    .X(_04322_));
 sky130_fd_sc_hd__xnor2_1 _12437_ (.A(_04318_),
    .B(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__o32a_1 _12438_ (.A1(_04014_),
    .A2(_04016_),
    .A3(_04024_),
    .B1(_04022_),
    .B2(_04021_),
    .X(_04324_));
 sky130_fd_sc_hd__a21oi_2 _12439_ (.A1(_04036_),
    .A2(_04034_),
    .B1(_04035_),
    .Y(_04325_));
 sky130_fd_sc_hd__o311ai_4 _12440_ (.A1(_03644_),
    .A2(_03826_),
    .A3(_04011_),
    .B1(_04013_),
    .C1(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__a211o_1 _12441_ (.A1(_03827_),
    .A2(_04013_),
    .B1(_04325_),
    .C1(_04011_),
    .X(_04327_));
 sky130_fd_sc_hd__a32o_1 _12442_ (.A1(_01499_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_01969_),
    .B2(_03320_),
    .X(_04328_));
 sky130_fd_sc_hd__nand3b_1 _12443_ (.A_N(_04005_),
    .B(_03653_),
    .C(_01969_),
    .Y(_04329_));
 sky130_fd_sc_hd__nand2_1 _12444_ (.A(_04328_),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__or4_1 _12445_ (.A(_00299_),
    .B(net56),
    .C(net166),
    .D(_03645_),
    .X(_04331_));
 sky130_fd_sc_hd__a21o_1 _12446_ (.A1(_04330_),
    .A2(_04331_),
    .B1(_04008_),
    .X(_04333_));
 sky130_fd_sc_hd__and3_1 _12447_ (.A(_04008_),
    .B(_04330_),
    .C(_04331_),
    .X(_04334_));
 sky130_fd_sc_hd__o211ai_1 _12448_ (.A1(net166),
    .A2(_03834_),
    .B1(_04008_),
    .C1(_04330_),
    .Y(_04335_));
 sky130_fd_sc_hd__a22o_1 _12449_ (.A1(_03820_),
    .A2(_03997_),
    .B1(_04333_),
    .B2(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__nand4_1 _12450_ (.A(_03997_),
    .B(_04335_),
    .C(_01969_),
    .D(_03087_),
    .Y(_04337_));
 sky130_fd_sc_hd__o21ai_1 _12451_ (.A1(_03998_),
    .A2(_04334_),
    .B1(_04336_),
    .Y(_04338_));
 sky130_fd_sc_hd__o2111ai_2 _12452_ (.A1(_03998_),
    .A2(_04334_),
    .B1(_04336_),
    .C1(_04326_),
    .D1(_04327_),
    .Y(_04339_));
 sky130_fd_sc_hd__a22o_1 _12453_ (.A1(_04326_),
    .A2(_04327_),
    .B1(_04336_),
    .B2(_04337_),
    .X(_04340_));
 sky130_fd_sc_hd__nand3_1 _12454_ (.A(_04340_),
    .B(_04324_),
    .C(_04339_),
    .Y(_04341_));
 sky130_fd_sc_hd__a21o_1 _12455_ (.A1(_04339_),
    .A2(_04340_),
    .B1(_04324_),
    .X(_04342_));
 sky130_fd_sc_hd__and3_1 _12456_ (.A(_04323_),
    .B(_04341_),
    .C(_04342_),
    .X(_04344_));
 sky130_fd_sc_hd__a21oi_1 _12457_ (.A1(_04341_),
    .A2(_04342_),
    .B1(_04323_),
    .Y(_04345_));
 sky130_fd_sc_hd__a32o_1 _12458_ (.A1(_03996_),
    .A2(_04030_),
    .A3(_04031_),
    .B1(_04033_),
    .B2(_04039_),
    .X(_04346_));
 sky130_fd_sc_hd__nor3_1 _12459_ (.A(_04346_),
    .B(_04345_),
    .C(_04344_),
    .Y(_04347_));
 sky130_fd_sc_hd__o21a_1 _12460_ (.A1(_04344_),
    .A2(_04345_),
    .B1(_04346_),
    .X(_04348_));
 sky130_fd_sc_hd__nor2_1 _12461_ (.A(_04347_),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__a31oi_2 _12462_ (.A1(_03853_),
    .A2(_04044_),
    .A3(_04046_),
    .B1(_04043_),
    .Y(_04350_));
 sky130_fd_sc_hd__xnor2_1 _12463_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__o311a_1 _12464_ (.A1(_07189_),
    .A2(_02433_),
    .A3(_03992_),
    .B1(_04317_),
    .C1(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__a21o_1 _12465_ (.A1(_04316_),
    .A2(_04317_),
    .B1(_04351_),
    .X(_04353_));
 sky130_fd_sc_hd__nand2b_1 _12466_ (.A_N(_04352_),
    .B(_04353_),
    .Y(_04355_));
 sky130_fd_sc_hd__a21bo_1 _12467_ (.A1(_04058_),
    .A2(_04076_),
    .B1_N(_04057_),
    .X(_04356_));
 sky130_fd_sc_hd__a32o_1 _12468_ (.A1(_00533_),
    .A2(_04087_),
    .A3(_00743_),
    .B1(_01038_),
    .B2(_04085_),
    .X(_04357_));
 sky130_fd_sc_hd__nand2b_1 _12469_ (.A_N(_04073_),
    .B(_04072_),
    .Y(_04358_));
 sky130_fd_sc_hd__nand3_1 _12470_ (.A(_04357_),
    .B(_04358_),
    .C(_04071_),
    .Y(_04359_));
 sky130_fd_sc_hd__a21o_1 _12471_ (.A1(_04071_),
    .A2(_04358_),
    .B1(_04357_),
    .X(_04360_));
 sky130_fd_sc_hd__a2bb2o_1 _12472_ (.A1_N(_03704_),
    .A2_N(_04066_),
    .B1(_07540_),
    .B2(_01544_),
    .X(_04361_));
 sky130_fd_sc_hd__and3_1 _12473_ (.A(_00072_),
    .B(_01539_),
    .C(_01541_),
    .X(_04362_));
 sky130_fd_sc_hd__o21ai_2 _12474_ (.A1(net149),
    .A2(_01662_),
    .B1(_04066_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand4_2 _12475_ (.A(_07540_),
    .B(_01879_),
    .C(net134),
    .D(_07440_),
    .Y(_04364_));
 sky130_fd_sc_hd__o21ai_1 _12476_ (.A1(_01662_),
    .A2(_04364_),
    .B1(_04363_),
    .Y(_04366_));
 sky130_fd_sc_hd__o21ai_2 _12477_ (.A1(net148),
    .A2(_01542_),
    .B1(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__o2111ai_4 _12478_ (.A1(_04364_),
    .A2(_01662_),
    .B1(_01544_),
    .C1(_00072_),
    .D1(_04363_),
    .Y(_04368_));
 sky130_fd_sc_hd__a22oi_2 _12479_ (.A1(_04065_),
    .A2(_04361_),
    .B1(_04367_),
    .B2(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__a22o_1 _12480_ (.A1(_04065_),
    .A2(_04361_),
    .B1(_04367_),
    .B2(_04368_),
    .X(_04370_));
 sky130_fd_sc_hd__nand4_2 _12481_ (.A(_04065_),
    .B(_04361_),
    .C(_04367_),
    .D(_04368_),
    .Y(_04371_));
 sky130_fd_sc_hd__a21o_1 _12482_ (.A1(_04370_),
    .A2(_04371_),
    .B1(_04063_),
    .X(_04372_));
 sky130_fd_sc_hd__or3b_1 _12483_ (.A(_04062_),
    .B(_04369_),
    .C_N(_04371_),
    .X(_04373_));
 sky130_fd_sc_hd__nand4_1 _12484_ (.A(_04359_),
    .B(_04360_),
    .C(_04372_),
    .D(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__a22o_1 _12485_ (.A1(_04359_),
    .A2(_04360_),
    .B1(_04372_),
    .B2(_04373_),
    .X(_04375_));
 sky130_fd_sc_hd__nand3_1 _12486_ (.A(_04375_),
    .B(_04356_),
    .C(_04374_),
    .Y(_04377_));
 sky130_fd_sc_hd__a21o_1 _12487_ (.A1(_04374_),
    .A2(_04375_),
    .B1(_04356_),
    .X(_04378_));
 sky130_fd_sc_hd__or4_1 _12488_ (.A(_00192_),
    .B(_00366_),
    .C(_01188_),
    .D(_01272_),
    .X(_04379_));
 sky130_fd_sc_hd__o32a_1 _12489_ (.A1(_00366_),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_01272_),
    .B2(_00192_),
    .X(_04380_));
 sky130_fd_sc_hd__a31o_1 _12490_ (.A1(_00367_),
    .A2(_01273_),
    .A3(_04060_),
    .B1(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__o21ai_1 _12491_ (.A1(_00532_),
    .A2(_01037_),
    .B1(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__or4_1 _12492_ (.A(_00532_),
    .B(_01033_),
    .C(_01035_),
    .D(_04381_),
    .X(_04383_));
 sky130_fd_sc_hd__nand2_1 _12493_ (.A(_04382_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a21oi_1 _12494_ (.A1(_04377_),
    .A2(_04378_),
    .B1(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _12495_ (.A(_04378_),
    .B(_04384_),
    .Y(_04386_));
 sky130_fd_sc_hd__nand3_1 _12496_ (.A(_04377_),
    .B(_04378_),
    .C(_04384_),
    .Y(_04388_));
 sky130_fd_sc_hd__nand2b_1 _12497_ (.A_N(_04385_),
    .B(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__and2_1 _12498_ (.A(_04084_),
    .B(_04090_),
    .X(_04390_));
 sky130_fd_sc_hd__a211oi_1 _12499_ (.A1(_04084_),
    .A2(_04090_),
    .B1(_04082_),
    .C1(_04389_),
    .Y(_04391_));
 sky130_fd_sc_hd__o21ai_1 _12500_ (.A1(_04082_),
    .A2(_04390_),
    .B1(_04389_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2b_2 _12501_ (.A_N(_04391_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__o21ai_4 _12502_ (.A1(_04096_),
    .A2(_04098_),
    .B1(_04095_),
    .Y(_04394_));
 sky130_fd_sc_hd__xor2_4 _12503_ (.A(_04393_),
    .B(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__inv_2 _12504_ (.A(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__nand3b_2 _12505_ (.A_N(_04352_),
    .B(_04353_),
    .C(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _12506_ (.A(_04355_),
    .B(_04395_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2_2 _12507_ (.A(_04397_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__a21oi_4 _12508_ (.A1(_04051_),
    .A2(_04099_),
    .B1(_04052_),
    .Y(_04401_));
 sky130_fd_sc_hd__a221oi_4 _12509_ (.A1(_04051_),
    .A2(_04099_),
    .B1(_04397_),
    .B2(_04399_),
    .C1(_04052_),
    .Y(_04402_));
 sky130_fd_sc_hd__xnor2_1 _12510_ (.A(_04400_),
    .B(_04401_),
    .Y(_04403_));
 sky130_fd_sc_hd__xor2_2 _12511_ (.A(_04315_),
    .B(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__or3b_4 _12512_ (.A(_04312_),
    .B(_04313_),
    .C_N(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__o21ba_2 _12513_ (.A1(_04312_),
    .A2(_04313_),
    .B1_N(_04404_),
    .X(_04406_));
 sky130_fd_sc_hd__or2_1 _12514_ (.A(_04311_),
    .B(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__o21ai_1 _12515_ (.A1(_04311_),
    .A2(_04406_),
    .B1(_04405_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21o_1 _12516_ (.A1(_04311_),
    .A2(_04406_),
    .B1(_04408_),
    .X(_04410_));
 sky130_fd_sc_hd__o21ai_2 _12517_ (.A1(_04311_),
    .A2(_04405_),
    .B1(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__inv_2 _12518_ (.A(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__nor2_1 _12519_ (.A(_04221_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__a22oi_1 _12520_ (.A1(_04412_),
    .A2(_04221_),
    .B1(_04220_),
    .B2(_04214_),
    .Y(_04414_));
 sky130_fd_sc_hd__o211ai_2 _12521_ (.A1(_04221_),
    .A2(_04412_),
    .B1(_04214_),
    .C1(_04220_),
    .Y(_04415_));
 sky130_fd_sc_hd__o21ai_1 _12522_ (.A1(_04223_),
    .A2(_04411_),
    .B1(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__a21oi_1 _12523_ (.A1(_04214_),
    .A2(_04220_),
    .B1(_04412_),
    .Y(_04417_));
 sky130_fd_sc_hd__o2bb2a_1 _12524_ (.A1_N(_04223_),
    .A2_N(_04417_),
    .B1(_04414_),
    .B2(_04413_),
    .X(_04418_));
 sky130_fd_sc_hd__a41o_1 _12525_ (.A1(_04214_),
    .A2(_04220_),
    .A3(_04221_),
    .A4(_04412_),
    .B1(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__or3_1 _12526_ (.A(_00834_),
    .B(_04219_),
    .C(_04419_),
    .X(_04421_));
 sky130_fd_sc_hd__o21ai_1 _12527_ (.A1(_00834_),
    .A2(_04219_),
    .B1(_04419_),
    .Y(_04422_));
 sky130_fd_sc_hd__and2_1 _12528_ (.A(_04421_),
    .B(_04422_),
    .X(net91));
 sky130_fd_sc_hd__a2bb2o_1 _12529_ (.A1_N(_00812_),
    .A2_N(_00823_),
    .B1(_04219_),
    .B2(_04419_),
    .X(_04423_));
 sky130_fd_sc_hd__o32a_1 _12530_ (.A1(_01033_),
    .A2(_01035_),
    .A3(_00570_),
    .B1(_00903_),
    .B2(_00744_),
    .X(_04424_));
 sky130_fd_sc_hd__and4_1 _12531_ (.A(_01038_),
    .B(_00743_),
    .C(_00569_),
    .D(_00904_),
    .X(_04425_));
 sky130_fd_sc_hd__o22ai_1 _12532_ (.A1(_00580_),
    .A2(_01058_),
    .B1(_04424_),
    .B2(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__or4_1 _12533_ (.A(_00580_),
    .B(_01058_),
    .C(_04424_),
    .D(_04425_),
    .X(_04427_));
 sky130_fd_sc_hd__nand2_1 _12534_ (.A(_04426_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_1 _12535_ (.A(_04428_),
    .B(_04312_),
    .Y(_04429_));
 sky130_fd_sc_hd__a41o_1 _12536_ (.A1(_00569_),
    .A2(_00581_),
    .A3(_00743_),
    .A4(_00904_),
    .B1(_04428_),
    .X(_04431_));
 sky130_fd_sc_hd__a21bo_1 _12537_ (.A1(_04372_),
    .A2(_04373_),
    .B1_N(_04360_),
    .X(_04432_));
 sky130_fd_sc_hd__or4_1 _12538_ (.A(_00532_),
    .B(_01033_),
    .C(_01035_),
    .D(_04380_),
    .X(_04433_));
 sky130_fd_sc_hd__o21a_1 _12539_ (.A1(_04063_),
    .A2(_04369_),
    .B1(_04371_),
    .X(_04434_));
 sky130_fd_sc_hd__a21oi_1 _12540_ (.A1(_04379_),
    .A2(_04433_),
    .B1(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__o2111ai_1 _12541_ (.A1(_04063_),
    .A2(_04369_),
    .B1(_04371_),
    .C1(_04379_),
    .D1(_04433_),
    .Y(_04436_));
 sky130_fd_sc_hd__and2b_1 _12542_ (.A_N(_04435_),
    .B(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__and3_1 _12543_ (.A(_00072_),
    .B(_01659_),
    .C(net140),
    .X(_04438_));
 sky130_fd_sc_hd__o2bb2a_1 _12544_ (.A1_N(_04363_),
    .A2_N(_04362_),
    .B1(_01662_),
    .B2(_07441_),
    .X(_04439_));
 sky130_fd_sc_hd__a211oi_1 _12545_ (.A1(_07534_),
    .A2(_07535_),
    .B1(_01882_),
    .C1(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__a32o_1 _12546_ (.A1(_07540_),
    .A2(_01879_),
    .A3(net134),
    .B1(_04363_),
    .B2(_04362_),
    .X(_04442_));
 sky130_fd_sc_hd__o31ai_1 _12547_ (.A1(net149),
    .A2(_01882_),
    .A3(_04439_),
    .B1(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__xnor2_1 _12548_ (.A(_04438_),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__xnor2_1 _12549_ (.A(_04437_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__nand3_1 _12550_ (.A(_04445_),
    .B(_04432_),
    .C(_04359_),
    .Y(_04446_));
 sky130_fd_sc_hd__a21o_1 _12551_ (.A1(_04359_),
    .A2(_04432_),
    .B1(_04445_),
    .X(_04447_));
 sky130_fd_sc_hd__and3_1 _12552_ (.A(_00533_),
    .B(_01185_),
    .C(_01187_),
    .X(_04448_));
 sky130_fd_sc_hd__and3_1 _12553_ (.A(_00367_),
    .B(_01539_),
    .C(_01541_),
    .X(_04449_));
 sky130_fd_sc_hd__and3_1 _12554_ (.A(_04449_),
    .B(_01273_),
    .C(_00193_),
    .X(_04450_));
 sky130_fd_sc_hd__o32a_1 _12555_ (.A1(_00192_),
    .A2(_01538_),
    .A3(_01540_),
    .B1(_00366_),
    .B2(_01272_),
    .X(_04451_));
 sky130_fd_sc_hd__a32o_1 _12556_ (.A1(_00193_),
    .A2(_01539_),
    .A3(_01541_),
    .B1(_00367_),
    .B2(_01273_),
    .X(_04453_));
 sky130_fd_sc_hd__o32a_1 _12557_ (.A1(_00532_),
    .A2(_01184_),
    .A3(_01186_),
    .B1(_04450_),
    .B2(_04451_),
    .X(_04454_));
 sky130_fd_sc_hd__or4_1 _12558_ (.A(_00532_),
    .B(_01188_),
    .C(_04450_),
    .D(_04451_),
    .X(_04455_));
 sky130_fd_sc_hd__and2b_1 _12559_ (.A_N(_04454_),
    .B(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__nand3_1 _12560_ (.A(_04446_),
    .B(_04447_),
    .C(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__a21o_1 _12561_ (.A1(_04446_),
    .A2(_04447_),
    .B1(_04456_),
    .X(_04458_));
 sky130_fd_sc_hd__and4_1 _12562_ (.A(_04377_),
    .B(_04386_),
    .C(_04457_),
    .D(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__a22o_1 _12563_ (.A1(_04377_),
    .A2(_04386_),
    .B1(_04457_),
    .B2(_04458_),
    .X(_04460_));
 sky130_fd_sc_hd__o21ai_2 _12564_ (.A1(_04391_),
    .A2(_04394_),
    .B1(_04392_),
    .Y(_04461_));
 sky130_fd_sc_hd__a21oi_2 _12565_ (.A1(_04461_),
    .A2(_04460_),
    .B1(_04459_),
    .Y(_04462_));
 sky130_fd_sc_hd__o21a_1 _12566_ (.A1(_04460_),
    .A2(_04461_),
    .B1(_04462_),
    .X(_04464_));
 sky130_fd_sc_hd__a21oi_2 _12567_ (.A1(_04459_),
    .A2(_04461_),
    .B1(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__or3_1 _12568_ (.A(_05327_),
    .B(_02692_),
    .C(_02694_),
    .X(_04466_));
 sky130_fd_sc_hd__o32a_1 _12569_ (.A1(_05327_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_07189_),
    .B2(_02433_),
    .X(_04467_));
 sky130_fd_sc_hd__and4_1 _12570_ (.A(_05316_),
    .B(_02432_),
    .C(_02697_),
    .D(_07200_),
    .X(_04468_));
 sky130_fd_sc_hd__or4_1 _12571_ (.A(_07441_),
    .B(_02096_),
    .C(_04467_),
    .D(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__o32a_1 _12572_ (.A1(_07441_),
    .A2(_02092_),
    .A3(_02094_),
    .B1(_04467_),
    .B2(_04468_),
    .X(_04470_));
 sky130_fd_sc_hd__a2bb2o_1 _12573_ (.A1_N(_04467_),
    .A2_N(_04468_),
    .B1(_07440_),
    .B2(_02097_),
    .X(_04471_));
 sky130_fd_sc_hd__a21oi_1 _12574_ (.A1(_04469_),
    .A2(_04471_),
    .B1(_04316_),
    .Y(_04472_));
 sky130_fd_sc_hd__o311a_1 _12575_ (.A1(_07189_),
    .A2(_02433_),
    .A3(_03992_),
    .B1(_04469_),
    .C1(_04471_),
    .X(_04473_));
 sky130_fd_sc_hd__or2_1 _12576_ (.A(_04472_),
    .B(_04473_),
    .X(_04475_));
 sky130_fd_sc_hd__a21boi_1 _12577_ (.A1(_04323_),
    .A2(_04341_),
    .B1_N(_04342_),
    .Y(_04476_));
 sky130_fd_sc_hd__a21bo_1 _12578_ (.A1(_04338_),
    .A2(_04327_),
    .B1_N(_04326_),
    .X(_04477_));
 sky130_fd_sc_hd__a32oi_4 _12579_ (.A1(_01969_),
    .A2(_03653_),
    .A3(_04005_),
    .B1(_03831_),
    .B2(_01499_),
    .Y(_04478_));
 sky130_fd_sc_hd__o31a_1 _12580_ (.A1(_04244_),
    .A2(_02696_),
    .A3(_04319_),
    .B1(_04320_),
    .X(_04479_));
 sky130_fd_sc_hd__o211ai_2 _12581_ (.A1(_03998_),
    .A2(_04334_),
    .B1(_04479_),
    .C1(_04333_),
    .Y(_04480_));
 sky130_fd_sc_hd__a21o_1 _12582_ (.A1(_04333_),
    .A2(_04337_),
    .B1(_04479_),
    .X(_04481_));
 sky130_fd_sc_hd__a21boi_1 _12583_ (.A1(_04481_),
    .A2(_04478_),
    .B1_N(_04480_),
    .Y(_04482_));
 sky130_fd_sc_hd__nand3_1 _12584_ (.A(_04481_),
    .B(_04478_),
    .C(_04480_),
    .Y(_04483_));
 sky130_fd_sc_hd__a21o_1 _12585_ (.A1(_04480_),
    .A2(_04481_),
    .B1(_04478_),
    .X(_04484_));
 sky130_fd_sc_hd__nand3_1 _12586_ (.A(_04477_),
    .B(_04483_),
    .C(_04484_),
    .Y(_04486_));
 sky130_fd_sc_hd__a21oi_1 _12587_ (.A1(_04483_),
    .A2(_04484_),
    .B1(_04477_),
    .Y(_04487_));
 sky130_fd_sc_hd__a21o_1 _12588_ (.A1(_04483_),
    .A2(_04484_),
    .B1(_04477_),
    .X(_04488_));
 sky130_fd_sc_hd__nand2_1 _12589_ (.A(_04486_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__or3_2 _12590_ (.A(_04244_),
    .B(_02920_),
    .C(_02923_),
    .X(_04490_));
 sky130_fd_sc_hd__and3_1 _12591_ (.A(_03917_),
    .B(_03316_),
    .C(_03318_),
    .X(_04491_));
 sky130_fd_sc_hd__or4_1 _12592_ (.A(_02636_),
    .B(_03906_),
    .C(_03086_),
    .D(_03319_),
    .X(_04492_));
 sky130_fd_sc_hd__o32a_1 _12593_ (.A1(_03906_),
    .A2(net132),
    .A3(net130),
    .B1(_03319_),
    .B2(_02636_),
    .X(_04493_));
 sky130_fd_sc_hd__a31o_1 _12594_ (.A1(_02647_),
    .A2(_03087_),
    .A3(_04491_),
    .B1(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__xor2_2 _12595_ (.A(_04490_),
    .B(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__and2_1 _12596_ (.A(_04489_),
    .B(_04495_),
    .X(_04497_));
 sky130_fd_sc_hd__nor2_1 _12597_ (.A(_04495_),
    .B(_04489_),
    .Y(_04498_));
 sky130_fd_sc_hd__o21a_1 _12598_ (.A1(_04497_),
    .A2(_04498_),
    .B1(_04476_),
    .X(_04499_));
 sky130_fd_sc_hd__o21ai_1 _12599_ (.A1(_04497_),
    .A2(_04498_),
    .B1(_04476_),
    .Y(_04500_));
 sky130_fd_sc_hd__a21o_1 _12600_ (.A1(_04489_),
    .A2(_04495_),
    .B1(_04476_),
    .X(_04501_));
 sky130_fd_sc_hd__o21ai_1 _12601_ (.A1(_04498_),
    .A2(_04501_),
    .B1(_04500_),
    .Y(_04502_));
 sky130_fd_sc_hd__o21bai_2 _12602_ (.A1(_04347_),
    .A2(_04350_),
    .B1_N(_04348_),
    .Y(_04503_));
 sky130_fd_sc_hd__xnor2_1 _12603_ (.A(_04502_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__nand2_1 _12604_ (.A(_04504_),
    .B(_04475_),
    .Y(_04505_));
 sky130_fd_sc_hd__nor2_1 _12605_ (.A(_04475_),
    .B(_04504_),
    .Y(_04506_));
 sky130_fd_sc_hd__xnor2_1 _12606_ (.A(_04475_),
    .B(_04504_),
    .Y(_04508_));
 sky130_fd_sc_hd__and2_1 _12607_ (.A(_04465_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__nor2_1 _12608_ (.A(_04465_),
    .B(_04508_),
    .Y(_04510_));
 sky130_fd_sc_hd__o21a_1 _12609_ (.A1(_04506_),
    .A2(_04465_),
    .B1(_04505_),
    .X(_04511_));
 sky130_fd_sc_hd__a21o_1 _12610_ (.A1(_04395_),
    .A2(_04353_),
    .B1(_04352_),
    .X(_04512_));
 sky130_fd_sc_hd__o21bai_4 _12611_ (.A1(_04509_),
    .A2(_04510_),
    .B1_N(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__nor3b_1 _12612_ (.A(_04509_),
    .B(_04510_),
    .C_N(_04512_),
    .Y(_04514_));
 sky130_fd_sc_hd__or3b_2 _12613_ (.A(_04509_),
    .B(_04510_),
    .C_N(_04512_),
    .X(_04515_));
 sky130_fd_sc_hd__a2bb2oi_4 _12614_ (.A1_N(_04400_),
    .A2_N(_04401_),
    .B1(_04101_),
    .B2(_04314_),
    .Y(_04516_));
 sky130_fd_sc_hd__a221oi_4 _12615_ (.A1(_04401_),
    .A2(_04400_),
    .B1(_04515_),
    .B2(_04513_),
    .C1(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__o211a_2 _12616_ (.A1(_04402_),
    .A2(_04516_),
    .B1(_04515_),
    .C1(_04513_),
    .X(_04519_));
 sky130_fd_sc_hd__o211a_1 _12617_ (.A1(_04517_),
    .A2(_04519_),
    .B1(_04429_),
    .C1(_04431_),
    .X(_04520_));
 sky130_fd_sc_hd__a211o_2 _12618_ (.A1(_04429_),
    .A2(_04431_),
    .B1(_04517_),
    .C1(_04519_),
    .X(_04521_));
 sky130_fd_sc_hd__and2b_1 _12619_ (.A_N(_04520_),
    .B(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__a21oi_2 _12620_ (.A1(_04251_),
    .A2(_04298_),
    .B1(_04300_),
    .Y(_04523_));
 sky130_fd_sc_hd__o21a_1 _12621_ (.A1(_04115_),
    .A2(_04228_),
    .B1(_04240_),
    .X(_04524_));
 sky130_fd_sc_hd__a21oi_1 _12622_ (.A1(_04115_),
    .A2(_04228_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__and3_1 _12623_ (.A(net156),
    .B(_03176_),
    .C(_03178_),
    .X(_04526_));
 sky130_fd_sc_hd__a32o_1 _12624_ (.A1(_02866_),
    .A2(_03180_),
    .A3(_04231_),
    .B1(net156),
    .B2(_02633_),
    .X(_04527_));
 sky130_fd_sc_hd__a32oi_2 _12625_ (.A1(_02866_),
    .A2(_03180_),
    .A3(_04231_),
    .B1(_04726_),
    .B2(_02858_),
    .Y(_04528_));
 sky130_fd_sc_hd__a31o_1 _12626_ (.A1(_04726_),
    .A2(_02858_),
    .A3(_04527_),
    .B1(_04528_),
    .X(_04530_));
 sky130_fd_sc_hd__xnor2_1 _12627_ (.A(_04526_),
    .B(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__nand4_1 _12628_ (.A(_03180_),
    .B(_03450_),
    .C(_04236_),
    .D(_02199_),
    .Y(_04532_));
 sky130_fd_sc_hd__a21bo_1 _12629_ (.A1(_04237_),
    .A2(_04532_),
    .B1_N(_04224_),
    .X(_04533_));
 sky130_fd_sc_hd__nand3b_1 _12630_ (.A_N(_04224_),
    .B(_04237_),
    .C(_04532_),
    .Y(_04534_));
 sky130_fd_sc_hd__and3b_1 _12631_ (.A_N(_04531_),
    .B(_04533_),
    .C(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__a21boi_1 _12632_ (.A1(_04533_),
    .A2(_04534_),
    .B1_N(_04531_),
    .Y(_04536_));
 sky130_fd_sc_hd__o21bai_1 _12633_ (.A1(_04535_),
    .A2(_04536_),
    .B1_N(_04525_),
    .Y(_04537_));
 sky130_fd_sc_hd__o32a_1 _12634_ (.A1(_02122_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(net159),
    .B2(_03449_),
    .X(_04538_));
 sky130_fd_sc_hd__or4_2 _12635_ (.A(_02811_),
    .B(_02833_),
    .C(_03581_),
    .D(_03582_),
    .X(_04539_));
 sky130_fd_sc_hd__and4_1 _12636_ (.A(_02133_),
    .B(_02866_),
    .C(_03450_),
    .D(_03584_),
    .X(_04541_));
 sky130_fd_sc_hd__o22a_1 _12637_ (.A1(_01620_),
    .A2(_03912_),
    .B1(_04538_),
    .B2(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__or3b_1 _12638_ (.A(_04535_),
    .B(_04536_),
    .C_N(_04525_),
    .X(_04543_));
 sky130_fd_sc_hd__nand2_1 _12639_ (.A(_04537_),
    .B(_04542_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _12640_ (.A(_04543_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand2_1 _12641_ (.A(_04537_),
    .B(_04543_),
    .Y(_04546_));
 sky130_fd_sc_hd__xnor2_1 _12642_ (.A(_04542_),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__o211ai_2 _12643_ (.A1(_04227_),
    .A2(_04241_),
    .B1(_04243_),
    .C1(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__a21o_1 _12644_ (.A1(_04242_),
    .A2(_04243_),
    .B1(_04547_),
    .X(_04549_));
 sky130_fd_sc_hd__a21o_1 _12645_ (.A1(_04150_),
    .A2(_04248_),
    .B1(_04249_),
    .X(_04550_));
 sky130_fd_sc_hd__nand3_1 _12646_ (.A(_04550_),
    .B(_04549_),
    .C(_04548_),
    .Y(_04552_));
 sky130_fd_sc_hd__a221o_1 _12647_ (.A1(_04248_),
    .A2(_04150_),
    .B1(_04549_),
    .B2(_04548_),
    .C1(_04249_),
    .X(_04553_));
 sky130_fd_sc_hd__nand2_2 _12648_ (.A(_04552_),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__or2_1 _12649_ (.A(_04284_),
    .B(_04291_),
    .X(_04555_));
 sky130_fd_sc_hd__nand2_1 _12650_ (.A(_04261_),
    .B(_04279_),
    .Y(_04556_));
 sky130_fd_sc_hd__nand2_1 _12651_ (.A(_04262_),
    .B(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__or3b_1 _12652_ (.A(net152),
    .B(_02053_),
    .C_N(_04286_),
    .X(_04558_));
 sky130_fd_sc_hd__nand2_1 _12653_ (.A(_04274_),
    .B(_04161_),
    .Y(_04559_));
 sky130_fd_sc_hd__a22o_1 _12654_ (.A1(_04287_),
    .A2(_04558_),
    .B1(_04559_),
    .B2(_04275_),
    .X(_04560_));
 sky130_fd_sc_hd__and4_1 _12655_ (.A(_04275_),
    .B(_04287_),
    .C(_04558_),
    .D(_04559_),
    .X(_04561_));
 sky130_fd_sc_hd__nand4_1 _12656_ (.A(_04275_),
    .B(_04287_),
    .C(_04558_),
    .D(_04559_),
    .Y(_04563_));
 sky130_fd_sc_hd__and3_1 _12657_ (.A(_00429_),
    .B(net145),
    .C(_01220_),
    .X(_04564_));
 sky130_fd_sc_hd__a32o_1 _12658_ (.A1(_00150_),
    .A2(_04265_),
    .A3(_01405_),
    .B1(net141),
    .B2(_00275_),
    .X(_04565_));
 sky130_fd_sc_hd__nand2_1 _12659_ (.A(_04565_),
    .B(_04564_),
    .Y(_04566_));
 sky130_fd_sc_hd__a31o_1 _12660_ (.A1(_00150_),
    .A2(_04265_),
    .A3(_01405_),
    .B1(_04564_),
    .X(_04567_));
 sky130_fd_sc_hd__a211o_1 _12661_ (.A1(_04566_),
    .A2(_04567_),
    .B1(_00274_),
    .C1(_01406_),
    .X(_04568_));
 sky130_fd_sc_hd__o211ai_2 _12662_ (.A1(_01406_),
    .A2(_00274_),
    .B1(_04567_),
    .C1(_04566_),
    .Y(_04569_));
 sky130_fd_sc_hd__and4_1 _12663_ (.A(_04560_),
    .B(_04563_),
    .C(_04568_),
    .D(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__a22oi_1 _12664_ (.A1(_04560_),
    .A2(_04563_),
    .B1(_04568_),
    .B2(_04569_),
    .Y(_04571_));
 sky130_fd_sc_hd__nor2_1 _12665_ (.A(_04570_),
    .B(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__xnor2_1 _12666_ (.A(_04557_),
    .B(_04572_),
    .Y(_04574_));
 sky130_fd_sc_hd__or4_1 _12667_ (.A(_07508_),
    .B(_07510_),
    .C(_02049_),
    .D(_02051_),
    .X(_04575_));
 sky130_fd_sc_hd__and3_1 _12668_ (.A(_00010_),
    .B(_00150_),
    .C(_01590_),
    .X(_04576_));
 sky130_fd_sc_hd__o32a_1 _12669_ (.A1(net144),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(_00009_),
    .X(_04577_));
 sky130_fd_sc_hd__a31o_1 _12670_ (.A1(_04576_),
    .A2(_01821_),
    .A3(_01820_),
    .B1(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__xnor2_1 _12671_ (.A(_04575_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__xor2_1 _12672_ (.A(_04574_),
    .B(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__a21oi_1 _12673_ (.A1(_04283_),
    .A2(_04555_),
    .B1(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__inv_2 _12674_ (.A(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__and3_1 _12675_ (.A(_04580_),
    .B(_04555_),
    .C(_04283_),
    .X(_04583_));
 sky130_fd_sc_hd__o21a_1 _12676_ (.A1(_04581_),
    .A2(_04583_),
    .B1(_04296_),
    .X(_04585_));
 sky130_fd_sc_hd__nor3_1 _12677_ (.A(_04581_),
    .B(_04583_),
    .C(_04296_),
    .Y(_04586_));
 sky130_fd_sc_hd__nor2_1 _12678_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__a32o_1 _12679_ (.A1(net151),
    .A2(net139),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_06341_),
    .X(_04588_));
 sky130_fd_sc_hd__or4_2 _12680_ (.A(_06331_),
    .B(net152),
    .C(_02241_),
    .D(_02355_),
    .X(_04589_));
 sky130_fd_sc_hd__a22oi_2 _12681_ (.A1(_05436_),
    .A2(_02633_),
    .B1(_04588_),
    .B2(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand4_1 _12682_ (.A(_05436_),
    .B(_02633_),
    .C(_04588_),
    .D(_04589_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand2b_1 _12683_ (.A_N(_04590_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__xor2_1 _12684_ (.A(_04252_),
    .B(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__or2_1 _12685_ (.A(_04593_),
    .B(_04587_),
    .X(_04594_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(_04587_),
    .B(_04593_),
    .Y(_04596_));
 sky130_fd_sc_hd__inv_2 _12687_ (.A(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand3_2 _12688_ (.A(_04554_),
    .B(_04594_),
    .C(_04596_),
    .Y(_04598_));
 sky130_fd_sc_hd__a21o_1 _12689_ (.A1(_04594_),
    .A2(_04596_),
    .B1(_04554_),
    .X(_04599_));
 sky130_fd_sc_hd__a21o_1 _12690_ (.A1(_04598_),
    .A2(_04599_),
    .B1(_04523_),
    .X(_04600_));
 sky130_fd_sc_hd__nand3_1 _12691_ (.A(_04599_),
    .B(_04523_),
    .C(_04598_),
    .Y(_04601_));
 sky130_fd_sc_hd__nand2_1 _12692_ (.A(_04600_),
    .B(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_2 _12693_ (.A1(_04306_),
    .A2(_04309_),
    .B1(_04305_),
    .Y(_04603_));
 sky130_fd_sc_hd__xnor2_2 _12694_ (.A(_04602_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__or2_1 _12695_ (.A(_04604_),
    .B(_04522_),
    .X(_04605_));
 sky130_fd_sc_hd__nand2_1 _12696_ (.A(_04522_),
    .B(_04604_),
    .Y(_04607_));
 sky130_fd_sc_hd__a22o_2 _12697_ (.A1(_04405_),
    .A2(_04407_),
    .B1(_04605_),
    .B2(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__o2111ai_4 _12698_ (.A1(_04406_),
    .A2(_04311_),
    .B1(_04405_),
    .C1(_04605_),
    .D1(_04607_),
    .Y(_04609_));
 sky130_fd_sc_hd__o211ai_4 _12699_ (.A1(_04411_),
    .A2(_04223_),
    .B1(_04609_),
    .C1(_04415_),
    .Y(_04610_));
 sky130_fd_sc_hd__o311a_1 _12700_ (.A1(_04413_),
    .A2(_04609_),
    .A3(_04414_),
    .B1(_04608_),
    .C1(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__o21ba_1 _12701_ (.A1(_04416_),
    .A2(_04608_),
    .B1_N(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__xor2_1 _12702_ (.A(_04423_),
    .B(_04612_),
    .X(net92));
 sky130_fd_sc_hd__nand3_1 _12703_ (.A(_04612_),
    .B(_04219_),
    .C(_04419_),
    .Y(_04613_));
 sky130_fd_sc_hd__a21oi_1 _12704_ (.A1(_04486_),
    .A2(_04495_),
    .B1(_04487_),
    .Y(_04614_));
 sky130_fd_sc_hd__or3_1 _12705_ (.A(_04244_),
    .B(net132),
    .C(net130),
    .X(_04615_));
 sky130_fd_sc_hd__o311a_1 _12706_ (.A1(_04244_),
    .A2(_02925_),
    .A3(_04493_),
    .B1(_04492_),
    .C1(_04329_),
    .X(_04617_));
 sky130_fd_sc_hd__a211oi_1 _12707_ (.A1(_04490_),
    .A2(_04492_),
    .B1(_04329_),
    .C1(_04493_),
    .Y(_04618_));
 sky130_fd_sc_hd__a31o_1 _12708_ (.A1(_02647_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_04491_),
    .X(_04619_));
 sky130_fd_sc_hd__or4_2 _12709_ (.A(_02636_),
    .B(_03906_),
    .C(_03319_),
    .D(_03652_),
    .X(_04620_));
 sky130_fd_sc_hd__a32o_1 _12710_ (.A1(_01936_),
    .A2(_03831_),
    .A3(_01947_),
    .B1(_04620_),
    .B2(_04619_),
    .X(_04621_));
 sky130_fd_sc_hd__o21a_1 _12711_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__nor3_1 _12712_ (.A(_04617_),
    .B(_04618_),
    .C(_04621_),
    .Y(_04623_));
 sky130_fd_sc_hd__or2_1 _12713_ (.A(_04622_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__and2_1 _12714_ (.A(_04482_),
    .B(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__nor2_1 _12715_ (.A(_04482_),
    .B(_04624_),
    .Y(_04626_));
 sky130_fd_sc_hd__o21ai_1 _12716_ (.A1(_04625_),
    .A2(_04626_),
    .B1(_04615_),
    .Y(_04628_));
 sky130_fd_sc_hd__or4_1 _12717_ (.A(_04244_),
    .B(_03086_),
    .C(_04625_),
    .D(_04626_),
    .X(_04629_));
 sky130_fd_sc_hd__a221oi_1 _12718_ (.A1(_04495_),
    .A2(_04486_),
    .B1(_04629_),
    .B2(_04628_),
    .C1(_04487_),
    .Y(_04630_));
 sky130_fd_sc_hd__a221o_1 _12719_ (.A1(_04495_),
    .A2(_04486_),
    .B1(_04629_),
    .B2(_04628_),
    .C1(_04487_),
    .X(_04631_));
 sky130_fd_sc_hd__nand3b_1 _12720_ (.A_N(_04614_),
    .B(_04628_),
    .C(_04629_),
    .Y(_04632_));
 sky130_fd_sc_hd__o21ai_1 _12721_ (.A1(_04498_),
    .A2(_04501_),
    .B1(_04503_),
    .Y(_04633_));
 sky130_fd_sc_hd__o22ai_1 _12722_ (.A1(_04501_),
    .A2(_04498_),
    .B1(_04499_),
    .B2(_04503_),
    .Y(_04634_));
 sky130_fd_sc_hd__nand4_1 _12723_ (.A(_04500_),
    .B(_04631_),
    .C(_04632_),
    .D(_04633_),
    .Y(_04635_));
 sky130_fd_sc_hd__a22o_1 _12724_ (.A1(_04631_),
    .A2(_04632_),
    .B1(_04633_),
    .B2(_04500_),
    .X(_04636_));
 sky130_fd_sc_hd__o32a_1 _12725_ (.A1(_05327_),
    .A2(_02920_),
    .A3(_02923_),
    .B1(_07189_),
    .B2(_02696_),
    .X(_04637_));
 sky130_fd_sc_hd__and3_1 _12726_ (.A(_07200_),
    .B(_02922_),
    .C(_02924_),
    .X(_04639_));
 sky130_fd_sc_hd__a31o_1 _12727_ (.A1(_05316_),
    .A2(_02697_),
    .A3(_04639_),
    .B1(_04637_),
    .X(_04640_));
 sky130_fd_sc_hd__o21a_1 _12728_ (.A1(_07441_),
    .A2(_02433_),
    .B1(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__or3_1 _12729_ (.A(_07441_),
    .B(_02433_),
    .C(_04640_),
    .X(_04642_));
 sky130_fd_sc_hd__nand2b_1 _12730_ (.A_N(_04641_),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__a21oi_1 _12731_ (.A1(_07540_),
    .A2(_02097_),
    .B1(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__and3_1 _12732_ (.A(_07540_),
    .B(_02097_),
    .C(_04643_),
    .X(_04645_));
 sky130_fd_sc_hd__or2_1 _12733_ (.A(_04644_),
    .B(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__a41o_1 _12734_ (.A1(_05316_),
    .A2(_07200_),
    .A3(_02432_),
    .A4(_02697_),
    .B1(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__or4b_1 _12735_ (.A(_07189_),
    .B(_02433_),
    .C(_04466_),
    .D_N(_04646_),
    .X(_04648_));
 sky130_fd_sc_hd__o41a_1 _12736_ (.A1(_07189_),
    .A2(_02433_),
    .A3(_03992_),
    .A4(_04470_),
    .B1(_04469_),
    .X(_04650_));
 sky130_fd_sc_hd__a21oi_1 _12737_ (.A1(_04647_),
    .A2(_04648_),
    .B1(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__and3_1 _12738_ (.A(_04647_),
    .B(_04648_),
    .C(_04650_),
    .X(_04652_));
 sky130_fd_sc_hd__nor2_1 _12739_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__a21o_1 _12740_ (.A1(_04635_),
    .A2(_04636_),
    .B1(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__inv_2 _12741_ (.A(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__and2_1 _12742_ (.A(_04635_),
    .B(_04653_),
    .X(_04656_));
 sky130_fd_sc_hd__and3_1 _12743_ (.A(_04635_),
    .B(_04636_),
    .C(_04653_),
    .X(_04657_));
 sky130_fd_sc_hd__a21boi_1 _12744_ (.A1(_04446_),
    .A2(_04456_),
    .B1_N(_04447_),
    .Y(_04658_));
 sky130_fd_sc_hd__a221o_1 _12745_ (.A1(net25),
    .A2(_00530_),
    .B1(_01266_),
    .B2(_01267_),
    .C1(_00527_),
    .X(_04659_));
 sky130_fd_sc_hd__a21o_1 _12746_ (.A1(_04444_),
    .A2(_04436_),
    .B1(_04435_),
    .X(_04661_));
 sky130_fd_sc_hd__a31o_1 _12747_ (.A1(_00072_),
    .A2(_01664_),
    .A3(_04442_),
    .B1(_04440_),
    .X(_04662_));
 sky130_fd_sc_hd__a31o_1 _12748_ (.A1(_00533_),
    .A2(_01189_),
    .A3(_04453_),
    .B1(_04450_),
    .X(_04663_));
 sky130_fd_sc_hd__o211a_1 _12749_ (.A1(_04448_),
    .A2(_04450_),
    .B1(_04453_),
    .C1(_04662_),
    .X(_04664_));
 sky130_fd_sc_hd__inv_2 _12750_ (.A(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__nor2_1 _12751_ (.A(_04662_),
    .B(_04663_),
    .Y(_04666_));
 sky130_fd_sc_hd__nor2_1 _12752_ (.A(_04664_),
    .B(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__or4_1 _12753_ (.A(net148),
    .B(_00192_),
    .C(_01662_),
    .D(_01882_),
    .X(_04668_));
 sky130_fd_sc_hd__o32a_1 _12754_ (.A1(_00192_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_01882_),
    .B2(net148),
    .X(_04669_));
 sky130_fd_sc_hd__a31o_1 _12755_ (.A1(_00193_),
    .A2(_01883_),
    .A3(_04438_),
    .B1(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__xnor2_1 _12756_ (.A(_04449_),
    .B(_04670_),
    .Y(_04672_));
 sky130_fd_sc_hd__xor2_1 _12757_ (.A(_04667_),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__nor2_1 _12758_ (.A(_04661_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_1 _12759_ (.A(_04673_),
    .B(_04661_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand2b_1 _12760_ (.A_N(_04674_),
    .B(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__xnor2_1 _12761_ (.A(_04659_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__and2_1 _12762_ (.A(_04658_),
    .B(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__nor2_1 _12763_ (.A(_04658_),
    .B(_04677_),
    .Y(_04679_));
 sky130_fd_sc_hd__nor2_1 _12764_ (.A(_04678_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__xor2_2 _12765_ (.A(_04462_),
    .B(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__o21ai_1 _12766_ (.A1(_04655_),
    .A2(_04657_),
    .B1(_04681_),
    .Y(_04683_));
 sky130_fd_sc_hd__a211o_1 _12767_ (.A1(_04636_),
    .A2(_04656_),
    .B1(_04655_),
    .C1(_04681_),
    .X(_04684_));
 sky130_fd_sc_hd__nand3b_2 _12768_ (.A_N(_04511_),
    .B(_04683_),
    .C(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__a21bo_1 _12769_ (.A1(_04683_),
    .A2(_04684_),
    .B1_N(_04511_),
    .X(_04686_));
 sky130_fd_sc_hd__o31a_1 _12770_ (.A1(_04402_),
    .A2(_04514_),
    .A3(_04516_),
    .B1(_04513_),
    .X(_04687_));
 sky130_fd_sc_hd__a21oi_1 _12771_ (.A1(_04685_),
    .A2(_04686_),
    .B1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__and3_1 _12772_ (.A(_04687_),
    .B(_04686_),
    .C(_04685_),
    .X(_04689_));
 sky130_fd_sc_hd__or2_2 _12773_ (.A(_04688_),
    .B(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__a32o_1 _12774_ (.A1(_00569_),
    .A2(_01185_),
    .A3(_01187_),
    .B1(_00904_),
    .B2(_01038_),
    .X(_04691_));
 sky130_fd_sc_hd__and4_1 _12775_ (.A(_00904_),
    .B(_01038_),
    .C(_01189_),
    .D(_00569_),
    .X(_04692_));
 sky130_fd_sc_hd__nand4_1 _12776_ (.A(_00904_),
    .B(_01038_),
    .C(_01189_),
    .D(_00569_),
    .Y(_04694_));
 sky130_fd_sc_hd__a32o_1 _12777_ (.A1(_00743_),
    .A2(_01055_),
    .A3(_01057_),
    .B1(_04691_),
    .B2(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__and4_1 _12778_ (.A(_01059_),
    .B(_04691_),
    .C(_04694_),
    .D(_00743_),
    .X(_04696_));
 sky130_fd_sc_hd__nand4_1 _12779_ (.A(_01059_),
    .B(_04691_),
    .C(_04694_),
    .D(_00743_),
    .Y(_04697_));
 sky130_fd_sc_hd__a32o_1 _12780_ (.A1(_00577_),
    .A2(_00579_),
    .A3(_01222_),
    .B1(_04695_),
    .B2(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__nand4_1 _12781_ (.A(_00581_),
    .B(_01222_),
    .C(_04695_),
    .D(_04697_),
    .Y(_04699_));
 sky130_fd_sc_hd__and3_1 _12782_ (.A(_04698_),
    .B(_04699_),
    .C(_04425_),
    .X(_04700_));
 sky130_fd_sc_hd__a21o_1 _12783_ (.A1(_04698_),
    .A2(_04699_),
    .B1(_04425_),
    .X(_04701_));
 sky130_fd_sc_hd__and2b_1 _12784_ (.A_N(_04700_),
    .B(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__a21bo_1 _12785_ (.A1(_04312_),
    .A2(_04426_),
    .B1_N(_04427_),
    .X(_04703_));
 sky130_fd_sc_hd__xnor2_2 _12786_ (.A(_04702_),
    .B(_04703_),
    .Y(_04705_));
 sky130_fd_sc_hd__nor2_1 _12787_ (.A(_04705_),
    .B(_04690_),
    .Y(_04706_));
 sky130_fd_sc_hd__nand2_1 _12788_ (.A(_04690_),
    .B(_04705_),
    .Y(_04707_));
 sky130_fd_sc_hd__and2b_1 _12789_ (.A_N(_04706_),
    .B(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__a32oi_4 _12790_ (.A1(_04523_),
    .A2(_04598_),
    .A3(_04599_),
    .B1(_04603_),
    .B2(_04600_),
    .Y(_04709_));
 sky130_fd_sc_hd__o21a_1 _12791_ (.A1(_04587_),
    .A2(_04593_),
    .B1(_04554_),
    .X(_04710_));
 sky130_fd_sc_hd__or4_1 _12792_ (.A(_00270_),
    .B(_00272_),
    .C(_01584_),
    .D(_01586_),
    .X(_04711_));
 sky130_fd_sc_hd__o32a_1 _12793_ (.A1(_00274_),
    .A2(_01584_),
    .A3(_01586_),
    .B1(net142),
    .B2(_01406_),
    .X(_04712_));
 sky130_fd_sc_hd__and4_1 _12794_ (.A(_01405_),
    .B(_01590_),
    .C(_00275_),
    .D(_00429_),
    .X(_04713_));
 sky130_fd_sc_hd__or4_1 _12795_ (.A(_00274_),
    .B(net142),
    .C(_01406_),
    .D(_01589_),
    .X(_04714_));
 sky130_fd_sc_hd__a311oi_1 _12796_ (.A1(_00150_),
    .A2(_01820_),
    .A3(_01821_),
    .B1(_04712_),
    .C1(_04713_),
    .Y(_04716_));
 sky130_fd_sc_hd__o211a_1 _12797_ (.A1(_04712_),
    .A2(_04713_),
    .B1(_00150_),
    .C1(_01823_),
    .X(_04717_));
 sky130_fd_sc_hd__nor2_1 _12798_ (.A(_04716_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__or3b_1 _12799_ (.A(_00274_),
    .B(_01406_),
    .C_N(_04567_),
    .X(_04719_));
 sky130_fd_sc_hd__o2bb2a_1 _12800_ (.A1_N(_01823_),
    .A2_N(_04576_),
    .B1(_04577_),
    .B2(_04575_),
    .X(_04720_));
 sky130_fd_sc_hd__a21oi_1 _12801_ (.A1(_04566_),
    .A2(_04719_),
    .B1(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__o21a_1 _12802_ (.A1(_04716_),
    .A2(_04717_),
    .B1(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__and3_1 _12803_ (.A(_04720_),
    .B(_04719_),
    .C(_04566_),
    .X(_04723_));
 sky130_fd_sc_hd__nand2_1 _12804_ (.A(_04723_),
    .B(_04718_),
    .Y(_04724_));
 sky130_fd_sc_hd__o21ba_1 _12805_ (.A1(_04718_),
    .A2(_04723_),
    .B1_N(_04721_),
    .X(_04725_));
 sky130_fd_sc_hd__a21oi_1 _12806_ (.A1(_04724_),
    .A2(_04725_),
    .B1(_04722_),
    .Y(_04727_));
 sky130_fd_sc_hd__a31o_1 _12807_ (.A1(_04560_),
    .A2(_04568_),
    .A3(_04569_),
    .B1(_04561_),
    .X(_04728_));
 sky130_fd_sc_hd__xnor2_1 _12808_ (.A(_04727_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__a21oi_1 _12809_ (.A1(_00010_),
    .A2(_02054_),
    .B1(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__and3_1 _12810_ (.A(_00010_),
    .B(_02054_),
    .C(_04729_),
    .X(_04731_));
 sky130_fd_sc_hd__nor2_1 _12811_ (.A(_04730_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__a21o_1 _12812_ (.A1(_04557_),
    .A2(_04572_),
    .B1(_04579_),
    .X(_04733_));
 sky130_fd_sc_hd__o21a_1 _12813_ (.A1(_04557_),
    .A2(_04572_),
    .B1(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__nor2_1 _12814_ (.A(_04732_),
    .B(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__and2_1 _12815_ (.A(_04732_),
    .B(_04734_),
    .X(_04736_));
 sky130_fd_sc_hd__nor2_1 _12816_ (.A(_04735_),
    .B(_04736_),
    .Y(_04738_));
 sky130_fd_sc_hd__a21oi_1 _12817_ (.A1(_04296_),
    .A2(_04582_),
    .B1(_04583_),
    .Y(_04739_));
 sky130_fd_sc_hd__xnor2_1 _12818_ (.A(_04738_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__a32o_1 _12819_ (.A1(_07513_),
    .A2(net139),
    .A3(_02237_),
    .B1(_02356_),
    .B2(net151),
    .X(_04741_));
 sky130_fd_sc_hd__or4_1 _12820_ (.A(net152),
    .B(_07512_),
    .C(_02241_),
    .D(_02355_),
    .X(_04742_));
 sky130_fd_sc_hd__a22oi_1 _12821_ (.A1(_06341_),
    .A2(_02633_),
    .B1(_04741_),
    .B2(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__o2111ai_1 _12822_ (.A1(_06265_),
    .A2(_06287_),
    .B1(_02633_),
    .C1(_04741_),
    .D1(_04742_),
    .Y(_04744_));
 sky130_fd_sc_hd__and2b_1 _12823_ (.A_N(_04743_),
    .B(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__a21oi_1 _12824_ (.A1(_05436_),
    .A2(_02858_),
    .B1(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__and3_1 _12825_ (.A(_04745_),
    .B(_02858_),
    .C(_05436_),
    .X(_04747_));
 sky130_fd_sc_hd__nor3_1 _12826_ (.A(_04589_),
    .B(_04746_),
    .C(_04747_),
    .Y(_04749_));
 sky130_fd_sc_hd__o21a_1 _12827_ (.A1(_04746_),
    .A2(_04747_),
    .B1(_04589_),
    .X(_04750_));
 sky130_fd_sc_hd__o21a_1 _12828_ (.A1(_04253_),
    .A2(_04590_),
    .B1(_04591_),
    .X(_04751_));
 sky130_fd_sc_hd__o221a_1 _12829_ (.A1(_04253_),
    .A2(_04590_),
    .B1(_04749_),
    .B2(_04750_),
    .C1(_04591_),
    .X(_04752_));
 sky130_fd_sc_hd__nor3_1 _12830_ (.A(_04749_),
    .B(_04751_),
    .C(_04750_),
    .Y(_04753_));
 sky130_fd_sc_hd__nor2_1 _12831_ (.A(_04752_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__xnor2_1 _12832_ (.A(_04740_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__o32a_1 _12833_ (.A1(net158),
    .A2(_03444_),
    .A3(_03447_),
    .B1(net155),
    .B2(_03179_),
    .X(_04756_));
 sky130_fd_sc_hd__or4_1 _12834_ (.A(net158),
    .B(net155),
    .C(_03179_),
    .D(_03449_),
    .X(_04757_));
 sky130_fd_sc_hd__a31o_1 _12835_ (.A1(_04726_),
    .A2(_03450_),
    .A3(_04526_),
    .B1(_04756_),
    .X(_04758_));
 sky130_fd_sc_hd__xor2_1 _12836_ (.A(_04539_),
    .B(_04758_),
    .X(_04760_));
 sky130_fd_sc_hd__a211oi_1 _12837_ (.A1(_03446_),
    .A2(_03468_),
    .B1(_03179_),
    .C1(_04528_),
    .Y(_04761_));
 sky130_fd_sc_hd__a31o_1 _12838_ (.A1(_04726_),
    .A2(_02858_),
    .A3(_04527_),
    .B1(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__nor2_1 _12839_ (.A(_04541_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__or4b_1 _12840_ (.A(_02122_),
    .B(_03449_),
    .C(_04539_),
    .D_N(_04762_),
    .X(_04764_));
 sky130_fd_sc_hd__nand2b_1 _12841_ (.A_N(_04763_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__a21oi_1 _12842_ (.A1(_04541_),
    .A2(_04762_),
    .B1(_04760_),
    .Y(_04766_));
 sky130_fd_sc_hd__xor2_1 _12843_ (.A(_04760_),
    .B(_04765_),
    .X(_04767_));
 sky130_fd_sc_hd__nand2_1 _12844_ (.A(_04531_),
    .B(_04534_),
    .Y(_04768_));
 sky130_fd_sc_hd__and2_1 _12845_ (.A(_04533_),
    .B(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__nor2_1 _12846_ (.A(_04769_),
    .B(_04767_),
    .Y(_04771_));
 sky130_fd_sc_hd__xnor2_1 _12847_ (.A(_04767_),
    .B(_04769_),
    .Y(_04772_));
 sky130_fd_sc_hd__or4_1 _12848_ (.A(_00321_),
    .B(net24),
    .C(_02122_),
    .D(_03580_),
    .X(_04773_));
 sky130_fd_sc_hd__o311a_1 _12849_ (.A1(_02079_),
    .A2(_02100_),
    .A3(_03912_),
    .B1(_04545_),
    .C1(_04772_),
    .X(_04774_));
 sky130_fd_sc_hd__a21o_1 _12850_ (.A1(_04772_),
    .A2(_04773_),
    .B1(_04545_),
    .X(_04775_));
 sky130_fd_sc_hd__nand2b_1 _12851_ (.A_N(_04774_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__a21boi_2 _12852_ (.A1(_04550_),
    .A2(_04548_),
    .B1_N(_04549_),
    .Y(_04777_));
 sky130_fd_sc_hd__xnor2_2 _12853_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__xnor2_1 _12854_ (.A(_04755_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__o21a_1 _12855_ (.A1(_04597_),
    .A2(_04710_),
    .B1(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__a211oi_1 _12856_ (.A1(_04554_),
    .A2(_04594_),
    .B1(_04597_),
    .C1(_04779_),
    .Y(_04782_));
 sky130_fd_sc_hd__nor2_1 _12857_ (.A(_04780_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__o21bai_1 _12858_ (.A1(_04709_),
    .A2(_04782_),
    .B1_N(_04780_),
    .Y(_04784_));
 sky130_fd_sc_hd__xor2_4 _12859_ (.A(_04709_),
    .B(_04783_),
    .X(_04785_));
 sky130_fd_sc_hd__xnor2_4 _12860_ (.A(_04708_),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__inv_2 _12861_ (.A(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__a21oi_2 _12862_ (.A1(_04521_),
    .A2(_04604_),
    .B1(_04520_),
    .Y(_04788_));
 sky130_fd_sc_hd__inv_2 _12863_ (.A(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__nor2_1 _12864_ (.A(_04788_),
    .B(_04787_),
    .Y(_04790_));
 sky130_fd_sc_hd__a211o_1 _12865_ (.A1(_04521_),
    .A2(_04604_),
    .B1(_04520_),
    .C1(_04786_),
    .X(_04791_));
 sky130_fd_sc_hd__nand2b_1 _12866_ (.A_N(_04790_),
    .B(_04791_),
    .Y(_04793_));
 sky130_fd_sc_hd__a21oi_1 _12867_ (.A1(_04608_),
    .A2(_04610_),
    .B1(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__a22o_1 _12868_ (.A1(_04789_),
    .A2(_04786_),
    .B1(_04610_),
    .B2(_04608_),
    .X(_04795_));
 sky130_fd_sc_hd__o211ai_2 _12869_ (.A1(_04786_),
    .A2(_04789_),
    .B1(_04608_),
    .C1(_04610_),
    .Y(_04796_));
 sky130_fd_sc_hd__a31oi_2 _12870_ (.A1(_04608_),
    .A2(_04610_),
    .A3(_04793_),
    .B1(_04794_),
    .Y(_04797_));
 sky130_fd_sc_hd__a31o_1 _12871_ (.A1(_04608_),
    .A2(_04610_),
    .A3(_04793_),
    .B1(_04794_),
    .X(_04798_));
 sky130_fd_sc_hd__and3_1 _12872_ (.A(_00845_),
    .B(_04613_),
    .C(_04797_),
    .X(_04799_));
 sky130_fd_sc_hd__a21oi_1 _12873_ (.A1(_00845_),
    .A2(_04613_),
    .B1(_04797_),
    .Y(_04800_));
 sky130_fd_sc_hd__nor2_1 _12874_ (.A(_04799_),
    .B(_04800_),
    .Y(net93));
 sky130_fd_sc_hd__a41o_1 _12875_ (.A1(_04612_),
    .A2(_04219_),
    .A3(_04419_),
    .A4(_04798_),
    .B1(_00834_),
    .X(_04801_));
 sky130_fd_sc_hd__o21ai_1 _12876_ (.A1(_04706_),
    .A2(_04785_),
    .B1(_04707_),
    .Y(_04803_));
 sky130_fd_sc_hd__o21a_1 _12877_ (.A1(_04657_),
    .A2(_04681_),
    .B1(_04654_),
    .X(_04804_));
 sky130_fd_sc_hd__o31ai_1 _12878_ (.A1(_00366_),
    .A2(_01542_),
    .A3(_04669_),
    .B1(_04668_),
    .Y(_04805_));
 sky130_fd_sc_hd__o21ai_1 _12879_ (.A1(_04662_),
    .A2(_04663_),
    .B1(_04672_),
    .Y(_04806_));
 sky130_fd_sc_hd__and3_1 _12880_ (.A(_00533_),
    .B(_01539_),
    .C(_01541_),
    .X(_04807_));
 sky130_fd_sc_hd__o32a_1 _12881_ (.A1(_00366_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_01882_),
    .B2(_00192_),
    .X(_04808_));
 sky130_fd_sc_hd__and4_1 _12882_ (.A(_00193_),
    .B(_00367_),
    .C(_01664_),
    .D(_01883_),
    .X(_04809_));
 sky130_fd_sc_hd__nor2_1 _12883_ (.A(_04808_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__xnor2_1 _12884_ (.A(_04807_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__a21oi_1 _12885_ (.A1(_04665_),
    .A2(_04806_),
    .B1(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__and3_1 _12886_ (.A(_04665_),
    .B(_04806_),
    .C(_04811_),
    .X(_04814_));
 sky130_fd_sc_hd__nor2_1 _12887_ (.A(_04805_),
    .B(_04812_),
    .Y(_04815_));
 sky130_fd_sc_hd__nor3_1 _12888_ (.A(_04812_),
    .B(_04814_),
    .C(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21ba_1 _12889_ (.A1(_04812_),
    .A2(_04814_),
    .B1_N(_04805_),
    .X(_04817_));
 sky130_fd_sc_hd__o31a_1 _12890_ (.A1(_00532_),
    .A2(_01272_),
    .A3(_04674_),
    .B1(_04675_),
    .X(_04818_));
 sky130_fd_sc_hd__o221a_1 _12891_ (.A1(_04816_),
    .A2(_04817_),
    .B1(_04659_),
    .B2(_04674_),
    .C1(_04675_),
    .X(_04819_));
 sky130_fd_sc_hd__or3_1 _12892_ (.A(_04816_),
    .B(_04817_),
    .C(_04818_),
    .X(_04820_));
 sky130_fd_sc_hd__nand2b_1 _12893_ (.A_N(_04819_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__o21ba_1 _12894_ (.A1(_04678_),
    .A2(_04462_),
    .B1_N(_04679_),
    .X(_04822_));
 sky130_fd_sc_hd__xnor2_2 _12895_ (.A(_04821_),
    .B(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__o21bai_1 _12896_ (.A1(_04618_),
    .A2(_04621_),
    .B1_N(_04617_),
    .Y(_04825_));
 sky130_fd_sc_hd__o22a_1 _12897_ (.A1(_04244_),
    .A2(_03319_),
    .B1(_03652_),
    .B2(_03906_),
    .X(_04826_));
 sky130_fd_sc_hd__and3_1 _12898_ (.A(_04491_),
    .B(_03653_),
    .C(_04255_),
    .X(_04827_));
 sky130_fd_sc_hd__o22a_1 _12899_ (.A1(_02636_),
    .A2(_03832_),
    .B1(_04826_),
    .B2(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__or2_1 _12900_ (.A(_04828_),
    .B(_04825_),
    .X(_04829_));
 sky130_fd_sc_hd__nand2_1 _12901_ (.A(_04825_),
    .B(_04828_),
    .Y(_04830_));
 sky130_fd_sc_hd__a21oi_1 _12902_ (.A1(_04829_),
    .A2(_04830_),
    .B1(_04620_),
    .Y(_04831_));
 sky130_fd_sc_hd__and3_1 _12903_ (.A(_04620_),
    .B(_04829_),
    .C(_04830_),
    .X(_04832_));
 sky130_fd_sc_hd__a21o_1 _12904_ (.A1(_04825_),
    .A2(_04828_),
    .B1(_04620_),
    .X(_04833_));
 sky130_fd_sc_hd__o21ba_1 _12905_ (.A1(_04615_),
    .A2(_04626_),
    .B1_N(_04625_),
    .X(_04834_));
 sky130_fd_sc_hd__or3b_1 _12906_ (.A(_04831_),
    .B(_04832_),
    .C_N(_04834_),
    .X(_04836_));
 sky130_fd_sc_hd__o21bai_1 _12907_ (.A1(_04831_),
    .A2(_04832_),
    .B1_N(_04834_),
    .Y(_04837_));
 sky130_fd_sc_hd__o21ai_1 _12908_ (.A1(_04630_),
    .A2(_04634_),
    .B1(_04632_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21oi_1 _12909_ (.A1(_04836_),
    .A2(_04837_),
    .B1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__and3_1 _12910_ (.A(_04838_),
    .B(_04837_),
    .C(_04836_),
    .X(_04840_));
 sky130_fd_sc_hd__or4_2 _12911_ (.A(_00067_),
    .B(_00069_),
    .C(_02092_),
    .D(_02094_),
    .X(_04841_));
 sky130_fd_sc_hd__and3_1 _12912_ (.A(_07540_),
    .B(_02427_),
    .C(_02428_),
    .X(_04842_));
 sky130_fd_sc_hd__and3_1 _12913_ (.A(_05316_),
    .B(_04639_),
    .C(_03087_),
    .X(_04843_));
 sky130_fd_sc_hd__nand4_1 _12914_ (.A(_07200_),
    .B(_02926_),
    .C(_03087_),
    .D(_05316_),
    .Y(_04844_));
 sky130_fd_sc_hd__a32o_1 _12915_ (.A1(_07200_),
    .A2(_02922_),
    .A3(_02924_),
    .B1(_03087_),
    .B2(_05316_),
    .X(_04845_));
 sky130_fd_sc_hd__a32o_1 _12916_ (.A1(_07440_),
    .A2(_02693_),
    .A3(_02695_),
    .B1(_04844_),
    .B2(_04845_),
    .X(_04847_));
 sky130_fd_sc_hd__nand4_2 _12917_ (.A(_02697_),
    .B(_04844_),
    .C(_04845_),
    .D(_07440_),
    .Y(_04848_));
 sky130_fd_sc_hd__a221o_1 _12918_ (.A1(_02430_),
    .A2(_02431_),
    .B1(_04847_),
    .B2(_04848_),
    .C1(net149),
    .X(_04849_));
 sky130_fd_sc_hd__o211ai_1 _12919_ (.A1(_02433_),
    .A2(net149),
    .B1(_04848_),
    .C1(_04847_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _12920_ (.A(_04849_),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__a31oi_1 _12921_ (.A1(_05316_),
    .A2(_02697_),
    .A3(_04639_),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__or4b_1 _12922_ (.A(_07189_),
    .B(_02925_),
    .C(_04466_),
    .D_N(_04851_),
    .X(_04853_));
 sky130_fd_sc_hd__nand2b_1 _12923_ (.A_N(_04852_),
    .B(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__xnor2_1 _12924_ (.A(_04841_),
    .B(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__o31a_1 _12925_ (.A1(net149),
    .A2(_02096_),
    .A3(_04641_),
    .B1(_04642_),
    .X(_04856_));
 sky130_fd_sc_hd__o311a_1 _12926_ (.A1(net149),
    .A2(_02096_),
    .A3(_04641_),
    .B1(_04642_),
    .C1(_04855_),
    .X(_04858_));
 sky130_fd_sc_hd__nand2_1 _12927_ (.A(_04855_),
    .B(_04856_),
    .Y(_04859_));
 sky130_fd_sc_hd__nor2_1 _12928_ (.A(_04855_),
    .B(_04856_),
    .Y(_04860_));
 sky130_fd_sc_hd__or2_1 _12929_ (.A(_04858_),
    .B(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__a21boi_2 _12930_ (.A1(_04648_),
    .A2(_04650_),
    .B1_N(_04647_),
    .Y(_04862_));
 sky130_fd_sc_hd__xor2_1 _12931_ (.A(_04861_),
    .B(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__nor3_1 _12932_ (.A(_04839_),
    .B(_04840_),
    .C(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__or3_1 _12933_ (.A(_04839_),
    .B(_04840_),
    .C(_04863_),
    .X(_04865_));
 sky130_fd_sc_hd__o21a_1 _12934_ (.A1(_04839_),
    .A2(_04840_),
    .B1(_04863_),
    .X(_04866_));
 sky130_fd_sc_hd__nor2_1 _12935_ (.A(_04866_),
    .B(_04823_),
    .Y(_04867_));
 sky130_fd_sc_hd__o21a_1 _12936_ (.A1(_04864_),
    .A2(_04866_),
    .B1(_04823_),
    .X(_04869_));
 sky130_fd_sc_hd__a21o_1 _12937_ (.A1(_04867_),
    .A2(_04865_),
    .B1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__nor2_1 _12938_ (.A(_04804_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand2_1 _12939_ (.A(_04870_),
    .B(_04804_),
    .Y(_04872_));
 sky130_fd_sc_hd__nand2b_2 _12940_ (.A_N(_04871_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__o311ai_4 _12941_ (.A1(_04402_),
    .A2(_04514_),
    .A3(_04516_),
    .B1(_04686_),
    .C1(_04513_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_2 _12942_ (.A(_04685_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__xnor2_4 _12943_ (.A(_04873_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21oi_2 _12944_ (.A1(_04701_),
    .A2(_04703_),
    .B1(_04700_),
    .Y(_04877_));
 sky130_fd_sc_hd__o22ai_4 _12945_ (.A1(_00903_),
    .A2(_01188_),
    .B1(_01272_),
    .B2(_00570_),
    .Y(_04878_));
 sky130_fd_sc_hd__nand4_4 _12946_ (.A(_00904_),
    .B(_01269_),
    .C(_01271_),
    .D(_00569_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand4_4 _12947_ (.A(_00904_),
    .B(_01189_),
    .C(_01273_),
    .D(_00569_),
    .Y(_04881_));
 sky130_fd_sc_hd__a22oi_4 _12948_ (.A1(_01038_),
    .A2(_01059_),
    .B1(_04878_),
    .B2(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__and4_1 _12949_ (.A(_01038_),
    .B(_01059_),
    .C(_04878_),
    .D(_04881_),
    .X(_04883_));
 sky130_fd_sc_hd__o2111ai_2 _12950_ (.A1(_04880_),
    .A2(_01188_),
    .B1(_01059_),
    .C1(_01038_),
    .D1(_04878_),
    .Y(_04884_));
 sky130_fd_sc_hd__o22ai_4 _12951_ (.A1(_00744_),
    .A2(_01221_),
    .B1(_04882_),
    .B2(_04883_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand4b_2 _12952_ (.A_N(_04882_),
    .B(_00743_),
    .C(_01222_),
    .D(_04884_),
    .Y(_04886_));
 sky130_fd_sc_hd__a21oi_2 _12953_ (.A1(_04885_),
    .A2(_04886_),
    .B1(_04692_),
    .Y(_04887_));
 sky130_fd_sc_hd__a21o_1 _12954_ (.A1(_04885_),
    .A2(_04886_),
    .B1(_04692_),
    .X(_04888_));
 sky130_fd_sc_hd__and3_1 _12955_ (.A(_04885_),
    .B(_04886_),
    .C(_04692_),
    .X(_04889_));
 sky130_fd_sc_hd__nand3_2 _12956_ (.A(_04885_),
    .B(_04886_),
    .C(_04692_),
    .Y(_04891_));
 sky130_fd_sc_hd__o2111ai_2 _12957_ (.A1(_04887_),
    .A2(_04889_),
    .B1(_00577_),
    .C1(_00579_),
    .D1(net137),
    .Y(_04892_));
 sky130_fd_sc_hd__o211ai_2 _12958_ (.A1(net136),
    .A2(_00580_),
    .B1(_04891_),
    .C1(_04888_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand2_1 _12959_ (.A(_04892_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__a31o_1 _12960_ (.A1(_00581_),
    .A2(_01222_),
    .A3(_04695_),
    .B1(_04696_),
    .X(_04895_));
 sky130_fd_sc_hd__inv_2 _12961_ (.A(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__xnor2_1 _12962_ (.A(_04894_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__a31oi_2 _12963_ (.A1(_04892_),
    .A2(_04893_),
    .A3(_04896_),
    .B1(_04877_),
    .Y(_04898_));
 sky130_fd_sc_hd__xnor2_2 _12964_ (.A(_04877_),
    .B(_04897_),
    .Y(_04899_));
 sky130_fd_sc_hd__nor2_1 _12965_ (.A(_04876_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__and2_1 _12966_ (.A(_04876_),
    .B(_04899_),
    .X(_04902_));
 sky130_fd_sc_hd__and4_1 _12967_ (.A(net156),
    .B(_04726_),
    .C(_03450_),
    .D(_03584_),
    .X(_04903_));
 sky130_fd_sc_hd__o32a_1 _12968_ (.A1(net158),
    .A2(_03581_),
    .A3(_03582_),
    .B1(net155),
    .B2(_03449_),
    .X(_04904_));
 sky130_fd_sc_hd__o22a_1 _12969_ (.A1(_03912_),
    .A2(net159),
    .B1(_04904_),
    .B2(_04903_),
    .X(_04905_));
 sky130_fd_sc_hd__o21a_1 _12970_ (.A1(_04763_),
    .A2(_04766_),
    .B1(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__or3_1 _12971_ (.A(_04763_),
    .B(_04766_),
    .C(_04905_),
    .X(_04907_));
 sky130_fd_sc_hd__and2b_1 _12972_ (.A_N(_04906_),
    .B(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__o31a_1 _12973_ (.A1(net159),
    .A2(_03583_),
    .A3(_04756_),
    .B1(_04757_),
    .X(_04909_));
 sky130_fd_sc_hd__xnor2_1 _12974_ (.A(_04908_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__or2_1 _12975_ (.A(_04771_),
    .B(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__or3b_1 _12976_ (.A(_04767_),
    .B(_04769_),
    .C_N(_04910_),
    .X(_04913_));
 sky130_fd_sc_hd__and2_1 _12977_ (.A(_04911_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__o21ai_2 _12978_ (.A1(_04774_),
    .A2(_04777_),
    .B1(_04775_),
    .Y(_04915_));
 sky130_fd_sc_hd__o21ai_1 _12979_ (.A1(_04771_),
    .A2(_04910_),
    .B1(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__xor2_2 _12980_ (.A(_04914_),
    .B(_04915_),
    .X(_04917_));
 sky130_fd_sc_hd__o32a_2 _12981_ (.A1(net142),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(_00274_),
    .X(_04918_));
 sky130_fd_sc_hd__and4_1 _12982_ (.A(_00275_),
    .B(_00429_),
    .C(_01590_),
    .D(_01823_),
    .X(_04919_));
 sky130_fd_sc_hd__o2111ai_2 _12983_ (.A1(_04918_),
    .A2(_04919_),
    .B1(_00146_),
    .C1(_00148_),
    .D1(_02054_),
    .Y(_04920_));
 sky130_fd_sc_hd__a311o_1 _12984_ (.A1(_00146_),
    .A2(_00148_),
    .A3(_02054_),
    .B1(_04918_),
    .C1(_04919_),
    .X(_04921_));
 sky130_fd_sc_hd__and3_1 _12985_ (.A(_04725_),
    .B(_04920_),
    .C(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__a21o_1 _12986_ (.A1(_04920_),
    .A2(_04921_),
    .B1(_04725_),
    .X(_04924_));
 sky130_fd_sc_hd__and2b_1 _12987_ (.A_N(_04922_),
    .B(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__o31a_1 _12988_ (.A1(net144),
    .A2(_01822_),
    .A3(_04712_),
    .B1(_04714_),
    .X(_04926_));
 sky130_fd_sc_hd__xnor2_1 _12989_ (.A(_04925_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__inv_2 _12990_ (.A(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__a2bb2o_1 _12991_ (.A1_N(_04728_),
    .A2_N(_04727_),
    .B1(_02054_),
    .B2(_00010_),
    .X(_04929_));
 sky130_fd_sc_hd__a21bo_1 _12992_ (.A1(_04727_),
    .A2(_04728_),
    .B1_N(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__nor2_1 _12993_ (.A(_04928_),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand2_1 _12994_ (.A(_04928_),
    .B(_04930_),
    .Y(_04932_));
 sky130_fd_sc_hd__o21bai_1 _12995_ (.A1(_04736_),
    .A2(_04739_),
    .B1_N(_04735_),
    .Y(_04933_));
 sky130_fd_sc_hd__and2b_1 _12996_ (.A_N(_04931_),
    .B(_04932_),
    .X(_04935_));
 sky130_fd_sc_hd__xnor2_1 _12997_ (.A(_04933_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__o31ai_1 _12998_ (.A1(_05425_),
    .A2(_02857_),
    .A3(_04743_),
    .B1(_04744_),
    .Y(_04937_));
 sky130_fd_sc_hd__a22o_2 _12999_ (.A1(_06276_),
    .A2(_06298_),
    .B1(_02852_),
    .B2(_02853_),
    .X(_04938_));
 sky130_fd_sc_hd__and3_1 _13000_ (.A(_00010_),
    .B(net139),
    .C(_02237_),
    .X(_04939_));
 sky130_fd_sc_hd__a31o_1 _13001_ (.A1(_07509_),
    .A2(_07511_),
    .A3(_02356_),
    .B1(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__or4_1 _13002_ (.A(_07512_),
    .B(_00009_),
    .C(_02241_),
    .D(_02355_),
    .X(_04941_));
 sky130_fd_sc_hd__and4_1 _13003_ (.A(net151),
    .B(_02633_),
    .C(_04940_),
    .D(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__a22oi_2 _13004_ (.A1(net151),
    .A2(_02633_),
    .B1(_04940_),
    .B2(_04941_),
    .Y(_04943_));
 sky130_fd_sc_hd__a311o_1 _13005_ (.A1(_06309_),
    .A2(_06320_),
    .A3(_02858_),
    .B1(_04942_),
    .C1(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__o221ai_1 _13006_ (.A1(_06265_),
    .A2(_06287_),
    .B1(_04942_),
    .B2(_04943_),
    .C1(_02858_),
    .Y(_04946_));
 sky130_fd_sc_hd__nand2_1 _13007_ (.A(_04944_),
    .B(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__a41o_1 _13008_ (.A1(net151),
    .A2(_07513_),
    .A3(_02240_),
    .A4(_02356_),
    .B1(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__nand2b_1 _13009_ (.A_N(_04742_),
    .B(_04947_),
    .Y(_04949_));
 sky130_fd_sc_hd__inv_2 _13010_ (.A(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nand2_1 _13011_ (.A(_04948_),
    .B(_04949_),
    .Y(_04951_));
 sky130_fd_sc_hd__o31a_1 _13012_ (.A1(_05425_),
    .A2(_03175_),
    .A3(_03177_),
    .B1(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__inv_2 _13013_ (.A(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__or4_1 _13014_ (.A(_05425_),
    .B(_03175_),
    .C(_03177_),
    .D(_04951_),
    .X(_04954_));
 sky130_fd_sc_hd__and3_1 _13015_ (.A(_04954_),
    .B(_04937_),
    .C(_04953_),
    .X(_04955_));
 sky130_fd_sc_hd__a21oi_1 _13016_ (.A1(_04953_),
    .A2(_04954_),
    .B1(_04937_),
    .Y(_04957_));
 sky130_fd_sc_hd__o21ba_1 _13017_ (.A1(_04751_),
    .A2(_04750_),
    .B1_N(_04749_),
    .X(_04958_));
 sky130_fd_sc_hd__or3b_1 _13018_ (.A(_04955_),
    .B(_04957_),
    .C_N(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__o21bai_1 _13019_ (.A1(_04955_),
    .A2(_04957_),
    .B1_N(_04958_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand3_1 _13020_ (.A(_04936_),
    .B(_04959_),
    .C(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__a21o_1 _13021_ (.A1(_04959_),
    .A2(_04960_),
    .B1(_04936_),
    .X(_04962_));
 sky130_fd_sc_hd__and2_1 _13022_ (.A(_04961_),
    .B(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__xnor2_1 _13023_ (.A(_04917_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__a21bo_1 _13024_ (.A1(_04740_),
    .A2(_04754_),
    .B1_N(_04778_),
    .X(_04965_));
 sky130_fd_sc_hd__o21ai_1 _13025_ (.A1(_04740_),
    .A2(_04754_),
    .B1(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__and2_1 _13026_ (.A(_04964_),
    .B(_04966_),
    .X(_04968_));
 sky130_fd_sc_hd__nor2_1 _13027_ (.A(_04966_),
    .B(_04964_),
    .Y(_04969_));
 sky130_fd_sc_hd__o21ai_1 _13028_ (.A1(_04968_),
    .A2(_04969_),
    .B1(_04784_),
    .Y(_04970_));
 sky130_fd_sc_hd__or3_1 _13029_ (.A(_04784_),
    .B(_04968_),
    .C(_04969_),
    .X(_04971_));
 sky130_fd_sc_hd__nand2_1 _13030_ (.A(_04970_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__o21ba_1 _13031_ (.A1(_04900_),
    .A2(_04902_),
    .B1_N(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__or3b_1 _13032_ (.A(_04900_),
    .B(_04902_),
    .C_N(_04972_),
    .X(_04974_));
 sky130_fd_sc_hd__and2b_1 _13033_ (.A_N(_04973_),
    .B(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__or2_2 _13034_ (.A(_04803_),
    .B(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__nand2_2 _13035_ (.A(_04803_),
    .B(_04975_),
    .Y(_04977_));
 sky130_fd_sc_hd__o211ai_4 _13036_ (.A1(_04788_),
    .A2(_04787_),
    .B1(_04977_),
    .C1(_04796_),
    .Y(_04979_));
 sky130_fd_sc_hd__a22o_1 _13037_ (.A1(_04791_),
    .A2(_04795_),
    .B1(_04976_),
    .B2(_04977_),
    .X(_04980_));
 sky130_fd_sc_hd__o2111ai_2 _13038_ (.A1(_04789_),
    .A2(_04786_),
    .B1(_04976_),
    .C1(_04795_),
    .D1(_04977_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2_1 _13039_ (.A(_04980_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__xnor2_1 _13040_ (.A(_04801_),
    .B(_04982_),
    .Y(net94));
 sky130_fd_sc_hd__nand4b_2 _13041_ (.A_N(_04613_),
    .B(_04798_),
    .C(_04980_),
    .D(_04981_),
    .Y(_04983_));
 sky130_fd_sc_hd__o21ba_1 _13042_ (.A1(_04900_),
    .A2(_04972_),
    .B1_N(_04902_),
    .X(_04984_));
 sky130_fd_sc_hd__o21bai_1 _13043_ (.A1(_04784_),
    .A2(_04968_),
    .B1_N(_04969_),
    .Y(_04985_));
 sky130_fd_sc_hd__a21bo_1 _13044_ (.A1(_04917_),
    .A2(_04961_),
    .B1_N(_04962_),
    .X(_04986_));
 sky130_fd_sc_hd__o21bai_1 _13045_ (.A1(_04938_),
    .A2(_04943_),
    .B1_N(_04942_),
    .Y(_04987_));
 sky130_fd_sc_hd__a32o_1 _13046_ (.A1(_06341_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(net151),
    .B2(_02858_),
    .X(_04989_));
 sky130_fd_sc_hd__o31a_1 _13047_ (.A1(net152),
    .A2(_03179_),
    .A3(_04938_),
    .B1(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__or4_1 _13048_ (.A(_00009_),
    .B(net144),
    .C(_02241_),
    .D(_02355_),
    .X(_04991_));
 sky130_fd_sc_hd__o32a_1 _13049_ (.A1(_00009_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(net144),
    .B2(_02241_),
    .X(_04992_));
 sky130_fd_sc_hd__a31o_1 _13050_ (.A1(_00150_),
    .A2(_02356_),
    .A3(_04939_),
    .B1(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__o31a_1 _13051_ (.A1(_07512_),
    .A2(_02628_),
    .A3(_02630_),
    .B1(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__and4b_1 _13052_ (.A_N(_04993_),
    .B(_02631_),
    .C(_02629_),
    .D(_07513_),
    .X(_04995_));
 sky130_fd_sc_hd__nor2_1 _13053_ (.A(_04994_),
    .B(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__or2_1 _13054_ (.A(_04990_),
    .B(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__o311a_1 _13055_ (.A1(net152),
    .A2(_03179_),
    .A3(_04938_),
    .B1(_04989_),
    .C1(_04996_),
    .X(_04998_));
 sky130_fd_sc_hd__nand2_1 _13056_ (.A(_04990_),
    .B(_04996_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _13057_ (.A(_04997_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__a31oi_1 _13058_ (.A1(_07513_),
    .A2(_02356_),
    .A3(_04939_),
    .B1(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__and4_1 _13059_ (.A(_04939_),
    .B(_05001_),
    .C(_07513_),
    .D(_02356_),
    .X(_05003_));
 sky130_fd_sc_hd__o21ai_1 _13060_ (.A1(_05002_),
    .A2(_05003_),
    .B1(_04987_),
    .Y(_05004_));
 sky130_fd_sc_hd__nor3_1 _13061_ (.A(_04987_),
    .B(_05002_),
    .C(_05003_),
    .Y(_05005_));
 sky130_fd_sc_hd__or3_1 _13062_ (.A(_04987_),
    .B(_05002_),
    .C(_05003_),
    .X(_05006_));
 sky130_fd_sc_hd__a211o_1 _13063_ (.A1(_05004_),
    .A2(_05006_),
    .B1(_05425_),
    .C1(_03449_),
    .X(_05007_));
 sky130_fd_sc_hd__o211ai_1 _13064_ (.A1(_05425_),
    .A2(_03449_),
    .B1(_05004_),
    .C1(_05006_),
    .Y(_05008_));
 sky130_fd_sc_hd__nand2_1 _13065_ (.A(_05007_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__a31o_1 _13066_ (.A1(_05436_),
    .A2(_03180_),
    .A3(_04948_),
    .B1(_04950_),
    .X(_05011_));
 sky130_fd_sc_hd__a311o_1 _13067_ (.A1(_05436_),
    .A2(_03180_),
    .A3(_04948_),
    .B1(_04950_),
    .C1(_05009_),
    .X(_05012_));
 sky130_fd_sc_hd__nand2_1 _13068_ (.A(_05009_),
    .B(_05011_),
    .Y(_05013_));
 sky130_fd_sc_hd__o21ba_1 _13069_ (.A1(_04957_),
    .A2(_04958_),
    .B1_N(_04955_),
    .X(_05014_));
 sky130_fd_sc_hd__nand3b_1 _13070_ (.A_N(_05014_),
    .B(_05013_),
    .C(_05012_),
    .Y(_05015_));
 sky130_fd_sc_hd__a21bo_1 _13071_ (.A1(_05012_),
    .A2(_05013_),
    .B1_N(_05014_),
    .X(_05016_));
 sky130_fd_sc_hd__or4_1 _13072_ (.A(_00145_),
    .B(_00147_),
    .C(_02053_),
    .D(_04918_),
    .X(_05017_));
 sky130_fd_sc_hd__a211oi_2 _13073_ (.A1(_04711_),
    .A2(_05017_),
    .B1(_00428_),
    .C1(_01822_),
    .Y(_05018_));
 sky130_fd_sc_hd__a211o_1 _13074_ (.A1(_04711_),
    .A2(_05017_),
    .B1(_00428_),
    .C1(_01822_),
    .X(_05019_));
 sky130_fd_sc_hd__o32a_1 _13075_ (.A1(net144),
    .A2(_02053_),
    .A3(_04918_),
    .B1(_00428_),
    .B2(_01822_),
    .X(_05020_));
 sky130_fd_sc_hd__o32a_2 _13076_ (.A1(_00270_),
    .A2(_00272_),
    .A3(_02053_),
    .B1(_05018_),
    .B2(_05020_),
    .X(_05022_));
 sky130_fd_sc_hd__a2111oi_4 _13077_ (.A1(_00267_),
    .A2(_00269_),
    .B1(_02053_),
    .C1(_05018_),
    .D1(_05020_),
    .Y(_05023_));
 sky130_fd_sc_hd__a32o_1 _13078_ (.A1(_04725_),
    .A2(_04920_),
    .A3(_04921_),
    .B1(_04924_),
    .B2(_04926_),
    .X(_05024_));
 sky130_fd_sc_hd__o21ai_1 _13079_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__or3_1 _13080_ (.A(_05022_),
    .B(_05023_),
    .C(_05024_),
    .X(_05026_));
 sky130_fd_sc_hd__o21ai_1 _13081_ (.A1(_04931_),
    .A2(_04933_),
    .B1(_04932_),
    .Y(_05027_));
 sky130_fd_sc_hd__a21oi_1 _13082_ (.A1(_05025_),
    .A2(_05026_),
    .B1(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__and3_1 _13083_ (.A(_05027_),
    .B(_05026_),
    .C(_05025_),
    .X(_05029_));
 sky130_fd_sc_hd__or2_1 _13084_ (.A(_05028_),
    .B(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__and3_1 _13085_ (.A(_05015_),
    .B(_05016_),
    .C(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__nand3_1 _13086_ (.A(_05015_),
    .B(_05016_),
    .C(_05030_),
    .Y(_05033_));
 sky130_fd_sc_hd__a21o_1 _13087_ (.A1(_05015_),
    .A2(_05016_),
    .B1(_05030_),
    .X(_05034_));
 sky130_fd_sc_hd__nand2_1 _13088_ (.A(_05033_),
    .B(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__a311o_1 _13089_ (.A1(net156),
    .A2(_03445_),
    .A3(_03448_),
    .B1(_03583_),
    .C1(net155),
    .X(_05036_));
 sky130_fd_sc_hd__o31a_1 _13090_ (.A1(_03479_),
    .A2(_03522_),
    .A3(_03912_),
    .B1(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__o21a_1 _13091_ (.A1(_04906_),
    .A2(_04909_),
    .B1(_04907_),
    .X(_05038_));
 sky130_fd_sc_hd__o311a_1 _13092_ (.A1(_03479_),
    .A2(_03522_),
    .A3(_03912_),
    .B1(_05036_),
    .C1(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__nor2_1 _13093_ (.A(_05037_),
    .B(_05038_),
    .Y(_05040_));
 sky130_fd_sc_hd__or2_1 _13094_ (.A(_05039_),
    .B(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__nand2_1 _13095_ (.A(_04913_),
    .B(_04916_),
    .Y(_05042_));
 sky130_fd_sc_hd__a21oi_1 _13096_ (.A1(_04913_),
    .A2(_04916_),
    .B1(_05041_),
    .Y(_05044_));
 sky130_fd_sc_hd__xnor2_2 _13097_ (.A(_05041_),
    .B(_05042_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_1 _13098_ (.A(_05045_),
    .B(_05034_),
    .Y(_05046_));
 sky130_fd_sc_hd__xnor2_1 _13099_ (.A(_05035_),
    .B(_05045_),
    .Y(_05047_));
 sky130_fd_sc_hd__nor2_1 _13100_ (.A(_04986_),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__inv_2 _13101_ (.A(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__a21o_1 _13102_ (.A1(_04986_),
    .A2(_05047_),
    .B1(_04985_),
    .X(_05050_));
 sky130_fd_sc_hd__nand3_1 _13103_ (.A(_04985_),
    .B(_04986_),
    .C(_05047_),
    .Y(_05051_));
 sky130_fd_sc_hd__o21a_1 _13104_ (.A1(_04986_),
    .A2(_05047_),
    .B1(_05050_),
    .X(_05052_));
 sky130_fd_sc_hd__a2bb2o_1 _13105_ (.A1_N(_04985_),
    .A2_N(_05049_),
    .B1(_05051_),
    .B2(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__o32a_2 _13106_ (.A1(_04839_),
    .A2(_04840_),
    .A3(_04863_),
    .B1(_04866_),
    .B2(_04823_),
    .X(_05055_));
 sky130_fd_sc_hd__or3_1 _13107_ (.A(_00532_),
    .B(_01658_),
    .C(_01660_),
    .X(_05056_));
 sky130_fd_sc_hd__o32a_1 _13108_ (.A1(_00532_),
    .A2(_01542_),
    .A3(_04808_),
    .B1(_01662_),
    .B2(_00192_),
    .X(_05057_));
 sky130_fd_sc_hd__o32a_1 _13109_ (.A1(_00532_),
    .A2(_01542_),
    .A3(_04808_),
    .B1(_01882_),
    .B2(_00366_),
    .X(_05058_));
 sky130_fd_sc_hd__o32ai_1 _13110_ (.A1(_00532_),
    .A2(_01542_),
    .A3(_04808_),
    .B1(_01882_),
    .B2(_00366_),
    .Y(_05059_));
 sky130_fd_sc_hd__o31a_1 _13111_ (.A1(_00366_),
    .A2(_01882_),
    .A3(_05057_),
    .B1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__xnor2_1 _13112_ (.A(_05056_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__o21ba_1 _13113_ (.A1(_04814_),
    .A2(_04815_),
    .B1_N(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__or3b_1 _13114_ (.A(_04814_),
    .B(_04815_),
    .C_N(_05061_),
    .X(_05063_));
 sky130_fd_sc_hd__and2b_1 _13115_ (.A_N(_05062_),
    .B(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__o21a_1 _13116_ (.A1(_04819_),
    .A2(_04822_),
    .B1(_04820_),
    .X(_05066_));
 sky130_fd_sc_hd__xor2_2 _13117_ (.A(_05064_),
    .B(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__or4_4 _13118_ (.A(_00188_),
    .B(_00190_),
    .C(_02092_),
    .D(_02094_),
    .X(_05068_));
 sky130_fd_sc_hd__o32a_1 _13119_ (.A1(net149),
    .A2(_02692_),
    .A3(_02694_),
    .B1(net148),
    .B2(_02433_),
    .X(_05069_));
 sky130_fd_sc_hd__a31oi_1 _13120_ (.A1(_00072_),
    .A2(_02697_),
    .A3(_04842_),
    .B1(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__and4_1 _13121_ (.A(_07200_),
    .B(_03087_),
    .C(_03320_),
    .D(_05316_),
    .X(_05071_));
 sky130_fd_sc_hd__o32a_1 _13122_ (.A1(_07189_),
    .A2(net132),
    .A3(net130),
    .B1(_05327_),
    .B2(_03319_),
    .X(_05072_));
 sky130_fd_sc_hd__a32o_1 _13123_ (.A1(_05316_),
    .A2(_03316_),
    .A3(_03318_),
    .B1(_07200_),
    .B2(_03087_),
    .X(_05073_));
 sky130_fd_sc_hd__a2bb2o_1 _13124_ (.A1_N(_05071_),
    .A2_N(_05072_),
    .B1(_07440_),
    .B2(_02926_),
    .X(_05074_));
 sky130_fd_sc_hd__or4bb_1 _13125_ (.A(_05071_),
    .B(_07441_),
    .C_N(_02926_),
    .D_N(_05073_),
    .X(_05075_));
 sky130_fd_sc_hd__a21o_1 _13126_ (.A1(_05074_),
    .A2(_05075_),
    .B1(_05070_),
    .X(_05077_));
 sky130_fd_sc_hd__nand3_1 _13127_ (.A(_05075_),
    .B(_05070_),
    .C(_05074_),
    .Y(_05078_));
 sky130_fd_sc_hd__and3_1 _13128_ (.A(_05077_),
    .B(_05078_),
    .C(_04843_),
    .X(_05079_));
 sky130_fd_sc_hd__a21oi_1 _13129_ (.A1(_05077_),
    .A2(_05078_),
    .B1(_04843_),
    .Y(_05080_));
 sky130_fd_sc_hd__or2_1 _13130_ (.A(_05079_),
    .B(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__or3b_1 _13131_ (.A(net149),
    .B(_02433_),
    .C_N(_04847_),
    .X(_05082_));
 sky130_fd_sc_hd__and3_1 _13132_ (.A(_05081_),
    .B(_05082_),
    .C(_04848_),
    .X(_05083_));
 sky130_fd_sc_hd__a21o_1 _13133_ (.A1(_04848_),
    .A2(_05082_),
    .B1(_05081_),
    .X(_05084_));
 sky130_fd_sc_hd__and2b_1 _13134_ (.A_N(_05083_),
    .B(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__xnor2_1 _13135_ (.A(_05068_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21ai_1 _13136_ (.A1(_04841_),
    .A2(_04852_),
    .B1(_04853_),
    .Y(_05088_));
 sky130_fd_sc_hd__nor2_1 _13137_ (.A(_05086_),
    .B(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__nand2_1 _13138_ (.A(_05086_),
    .B(_05088_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2b_1 _13139_ (.A_N(_05089_),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__a21oi_1 _13140_ (.A1(_04859_),
    .A2(_04862_),
    .B1(_04860_),
    .Y(_05092_));
 sky130_fd_sc_hd__and2b_1 _13141_ (.A_N(_05092_),
    .B(_05091_),
    .X(_05093_));
 sky130_fd_sc_hd__a211oi_2 _13142_ (.A1(_04859_),
    .A2(_04862_),
    .B1(_04860_),
    .C1(_05091_),
    .Y(_05094_));
 sky130_fd_sc_hd__o32a_1 _13143_ (.A1(_04244_),
    .A2(_03652_),
    .A3(_04491_),
    .B1(_03832_),
    .B2(_03906_),
    .X(_05095_));
 sky130_fd_sc_hd__a21oi_1 _13144_ (.A1(_04829_),
    .A2(_04833_),
    .B1(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__and3_1 _13145_ (.A(_04829_),
    .B(_04833_),
    .C(_05095_),
    .X(_05097_));
 sky130_fd_sc_hd__a21boi_2 _13146_ (.A1(_04838_),
    .A2(_04836_),
    .B1_N(_04837_),
    .Y(_05099_));
 sky130_fd_sc_hd__o21ai_2 _13147_ (.A1(_05096_),
    .A2(_05097_),
    .B1(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nor2_1 _13148_ (.A(_05097_),
    .B(_05099_),
    .Y(_05101_));
 sky130_fd_sc_hd__inv_2 _13149_ (.A(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__o221ai_4 _13150_ (.A1(_05099_),
    .A2(_05097_),
    .B1(_05094_),
    .B2(_05093_),
    .C1(_05100_),
    .Y(_05103_));
 sky130_fd_sc_hd__inv_2 _13151_ (.A(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__a211oi_2 _13152_ (.A1(_05100_),
    .A2(_05102_),
    .B1(_05093_),
    .C1(_05094_),
    .Y(_05105_));
 sky130_fd_sc_hd__nor2_1 _13153_ (.A(_05067_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__o21a_1 _13154_ (.A1(_05104_),
    .A2(_05105_),
    .B1(_05067_),
    .X(_05107_));
 sky130_fd_sc_hd__a21o_1 _13155_ (.A1(_05106_),
    .A2(_05103_),
    .B1(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__a211o_1 _13156_ (.A1(_04823_),
    .A2(_04865_),
    .B1(_04866_),
    .C1(_05108_),
    .X(_05110_));
 sky130_fd_sc_hd__xnor2_2 _13157_ (.A(_05055_),
    .B(_05108_),
    .Y(_05111_));
 sky130_fd_sc_hd__a22oi_1 _13158_ (.A1(_04804_),
    .A2(_04870_),
    .B1(_04874_),
    .B2(_04685_),
    .Y(_05112_));
 sky130_fd_sc_hd__a21o_1 _13159_ (.A1(_04875_),
    .A2(_04872_),
    .B1(_04871_),
    .X(_05113_));
 sky130_fd_sc_hd__xnor2_4 _13160_ (.A(_05111_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__a21oi_4 _13161_ (.A1(_04894_),
    .A2(_04895_),
    .B1(_04898_),
    .Y(_05115_));
 sky130_fd_sc_hd__and3_1 _13162_ (.A(net137),
    .B(_00740_),
    .C(_00739_),
    .X(_05116_));
 sky130_fd_sc_hd__a31o_1 _13163_ (.A1(_01034_),
    .A2(_01036_),
    .A3(_01222_),
    .B1(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__nand4_2 _13164_ (.A(_00743_),
    .B(_01038_),
    .C(net137),
    .D(_01222_),
    .Y(_05118_));
 sky130_fd_sc_hd__nand2_1 _13165_ (.A(_05117_),
    .B(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__and3_1 _13166_ (.A(_01059_),
    .B(_01185_),
    .C(_01187_),
    .X(_05121_));
 sky130_fd_sc_hd__a221oi_1 _13167_ (.A1(_00567_),
    .A2(_00568_),
    .B1(_01535_),
    .B2(_01537_),
    .C1(_01540_),
    .Y(_05122_));
 sky130_fd_sc_hd__a32o_1 _13168_ (.A1(_00569_),
    .A2(_01539_),
    .A3(_01541_),
    .B1(_00904_),
    .B2(_01273_),
    .X(_05123_));
 sky130_fd_sc_hd__o21ai_1 _13169_ (.A1(_01542_),
    .A2(_04880_),
    .B1(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__o21ai_1 _13170_ (.A1(_01058_),
    .A2(_01188_),
    .B1(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__o2111ai_1 _13171_ (.A1(_04880_),
    .A2(_01542_),
    .B1(_01189_),
    .C1(_01059_),
    .D1(_05123_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand2_1 _13172_ (.A(_05124_),
    .B(_05121_),
    .Y(_05127_));
 sky130_fd_sc_hd__o221ai_2 _13173_ (.A1(_01058_),
    .A2(_01188_),
    .B1(_01542_),
    .B2(_04880_),
    .C1(_05123_),
    .Y(_05128_));
 sky130_fd_sc_hd__nand4_1 _13174_ (.A(_05117_),
    .B(_05118_),
    .C(_05125_),
    .D(_05126_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand3_1 _13175_ (.A(_05119_),
    .B(_05127_),
    .C(_05128_),
    .Y(_05130_));
 sky130_fd_sc_hd__nand4_1 _13176_ (.A(_05117_),
    .B(_05118_),
    .C(_05127_),
    .D(_05128_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand3_1 _13177_ (.A(_05119_),
    .B(_05125_),
    .C(_05126_),
    .Y(_05133_));
 sky130_fd_sc_hd__o211ai_1 _13178_ (.A1(_01188_),
    .A2(_04880_),
    .B1(_05129_),
    .C1(_05130_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand3b_1 _13179_ (.A_N(_04881_),
    .B(_05132_),
    .C(_05133_),
    .Y(_05135_));
 sky130_fd_sc_hd__o31a_1 _13180_ (.A1(_00744_),
    .A2(_01221_),
    .A3(_04882_),
    .B1(_04884_),
    .X(_05136_));
 sky130_fd_sc_hd__nand3_1 _13181_ (.A(_05134_),
    .B(_05135_),
    .C(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__a21o_2 _13182_ (.A1(_05134_),
    .A2(_05135_),
    .B1(_05136_),
    .X(_05138_));
 sky130_fd_sc_hd__nand4_2 _13183_ (.A(_00581_),
    .B(_01590_),
    .C(_05137_),
    .D(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__a32o_1 _13184_ (.A1(_00581_),
    .A2(_01585_),
    .A3(_01588_),
    .B1(_05137_),
    .B2(_05138_),
    .X(_05140_));
 sky130_fd_sc_hd__nand2_1 _13185_ (.A(_05139_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__o31ai_2 _13186_ (.A1(_00580_),
    .A2(net136),
    .A3(_04887_),
    .B1(_04891_),
    .Y(_05143_));
 sky130_fd_sc_hd__o31a_1 _13187_ (.A1(_00580_),
    .A2(net136),
    .A3(_04887_),
    .B1(_04891_),
    .X(_05144_));
 sky130_fd_sc_hd__nand3_2 _13188_ (.A(_05139_),
    .B(_05140_),
    .C(_05143_),
    .Y(_05145_));
 sky130_fd_sc_hd__a21o_1 _13189_ (.A1(_05139_),
    .A2(_05140_),
    .B1(_05143_),
    .X(_05146_));
 sky130_fd_sc_hd__nand2_2 _13190_ (.A(_05145_),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__xor2_4 _13191_ (.A(_05115_),
    .B(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__and2_2 _13192_ (.A(_05114_),
    .B(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__nor2_2 _13193_ (.A(_05148_),
    .B(_05114_),
    .Y(_05150_));
 sky130_fd_sc_hd__o21ai_1 _13194_ (.A1(_05149_),
    .A2(_05150_),
    .B1(_05053_),
    .Y(_05151_));
 sky130_fd_sc_hd__nor2_2 _13195_ (.A(_05150_),
    .B(_05053_),
    .Y(_05152_));
 sky130_fd_sc_hd__o31ai_4 _13196_ (.A1(_05053_),
    .A2(_05149_),
    .A3(_05150_),
    .B1(_05151_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand2_2 _13197_ (.A(_04984_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__inv_2 _13198_ (.A(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__nor2_1 _13199_ (.A(_04984_),
    .B(_05154_),
    .Y(_05157_));
 sky130_fd_sc_hd__o221ai_1 _13200_ (.A1(_04803_),
    .A2(_04975_),
    .B1(_05156_),
    .B2(_05157_),
    .C1(_04979_),
    .Y(_05158_));
 sky130_fd_sc_hd__a211o_1 _13201_ (.A1(_04976_),
    .A2(_04979_),
    .B1(_05156_),
    .C1(_05157_),
    .X(_05159_));
 sky130_fd_sc_hd__o211ai_4 _13202_ (.A1(_04984_),
    .A2(_05154_),
    .B1(_04976_),
    .C1(_04979_),
    .Y(_05160_));
 sky130_fd_sc_hd__and2_1 _13203_ (.A(_05158_),
    .B(_05159_),
    .X(_05161_));
 sky130_fd_sc_hd__o311a_1 _13204_ (.A1(_04613_),
    .A2(_04797_),
    .A3(_04982_),
    .B1(_05161_),
    .C1(_00845_),
    .X(_05162_));
 sky130_fd_sc_hd__a21oi_1 _13205_ (.A1(_00845_),
    .A2(_04983_),
    .B1(_05161_),
    .Y(_05163_));
 sky130_fd_sc_hd__nor2_1 _13206_ (.A(_05162_),
    .B(_05163_),
    .Y(net95));
 sky130_fd_sc_hd__a21o_1 _13207_ (.A1(_05158_),
    .A2(_05159_),
    .B1(_04983_),
    .X(_05165_));
 sky130_fd_sc_hd__o21ai_2 _13208_ (.A1(_05067_),
    .A2(_05105_),
    .B1(_05103_),
    .Y(_05166_));
 sky130_fd_sc_hd__o32ai_1 _13209_ (.A1(_00366_),
    .A2(_01882_),
    .A3(_05057_),
    .B1(_05058_),
    .B2(_05056_),
    .Y(_05167_));
 sky130_fd_sc_hd__a31o_1 _13210_ (.A1(_00533_),
    .A2(_01879_),
    .A3(net134),
    .B1(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__or3b_2 _13211_ (.A(_00532_),
    .B(_01882_),
    .C_N(_05167_),
    .X(_05169_));
 sky130_fd_sc_hd__o21ai_2 _13212_ (.A1(_05062_),
    .A2(_05066_),
    .B1(_05063_),
    .Y(_05170_));
 sky130_fd_sc_hd__a21o_1 _13213_ (.A1(_05168_),
    .A2(_05169_),
    .B1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nand3_1 _13214_ (.A(_05170_),
    .B(_05169_),
    .C(_05168_),
    .Y(_05172_));
 sky130_fd_sc_hd__and2_1 _13215_ (.A(_05171_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__a2111oi_1 _13216_ (.A1(_04255_),
    .A2(_03831_),
    .B1(_04827_),
    .C1(_05096_),
    .D1(_05101_),
    .Y(_05175_));
 sky130_fd_sc_hd__a2111o_1 _13217_ (.A1(_04255_),
    .A2(_03831_),
    .B1(_04827_),
    .C1(_05096_),
    .D1(_05101_),
    .X(_05176_));
 sky130_fd_sc_hd__a21boi_1 _13218_ (.A1(_05077_),
    .A2(_04843_),
    .B1_N(_05078_),
    .Y(_05177_));
 sky130_fd_sc_hd__a31o_1 _13219_ (.A1(_05073_),
    .A2(_07440_),
    .A3(_02926_),
    .B1(_05071_),
    .X(_05178_));
 sky130_fd_sc_hd__a31oi_1 _13220_ (.A1(_00072_),
    .A2(_02697_),
    .A3(_04842_),
    .B1(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__a31o_1 _13221_ (.A1(_00072_),
    .A2(_02697_),
    .A3(_04842_),
    .B1(_05178_),
    .X(_05180_));
 sky130_fd_sc_hd__and4_1 _13222_ (.A(_04842_),
    .B(_05178_),
    .C(_00072_),
    .D(_02697_),
    .X(_05181_));
 sky130_fd_sc_hd__nor2_1 _13223_ (.A(_05179_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__a32o_1 _13224_ (.A1(_05316_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_07200_),
    .B2(_03320_),
    .X(_05183_));
 sky130_fd_sc_hd__or3_1 _13225_ (.A(_07146_),
    .B(_07168_),
    .C(_03652_),
    .X(_05184_));
 sky130_fd_sc_hd__and4_1 _13226_ (.A(_07200_),
    .B(_03320_),
    .C(_03653_),
    .D(_05316_),
    .X(_05186_));
 sky130_fd_sc_hd__o31ai_1 _13227_ (.A1(_05327_),
    .A2(_03319_),
    .A3(_05184_),
    .B1(_05183_),
    .Y(_05187_));
 sky130_fd_sc_hd__and4b_1 _13228_ (.A_N(_05187_),
    .B(_03087_),
    .C(_07437_),
    .D(net162),
    .X(_05188_));
 sky130_fd_sc_hd__o31a_1 _13229_ (.A1(_07441_),
    .A2(net132),
    .A3(net130),
    .B1(_05187_),
    .X(_05189_));
 sky130_fd_sc_hd__o21ai_1 _13230_ (.A1(_07441_),
    .A2(_03086_),
    .B1(_05187_),
    .Y(_05190_));
 sky130_fd_sc_hd__o32a_1 _13231_ (.A1(net149),
    .A2(_02920_),
    .A3(_02923_),
    .B1(_05188_),
    .B2(_05189_),
    .X(_05191_));
 sky130_fd_sc_hd__a2111oi_1 _13232_ (.A1(_07534_),
    .A2(_07535_),
    .B1(_02925_),
    .C1(_05188_),
    .D1(_05189_),
    .Y(_05192_));
 sky130_fd_sc_hd__nor2_1 _13233_ (.A(_05191_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__xnor2_1 _13234_ (.A(_05182_),
    .B(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__and2_1 _13235_ (.A(_05177_),
    .B(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__nor2_1 _13236_ (.A(_05177_),
    .B(_05194_),
    .Y(_05197_));
 sky130_fd_sc_hd__or4_1 _13237_ (.A(_00361_),
    .B(_00363_),
    .C(net133),
    .D(_02094_),
    .X(_05198_));
 sky130_fd_sc_hd__o32a_1 _13238_ (.A1(net148),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_00192_),
    .B2(_02433_),
    .X(_05199_));
 sky130_fd_sc_hd__or4_1 _13239_ (.A(net148),
    .B(_00192_),
    .C(_02433_),
    .D(_02696_),
    .X(_05200_));
 sky130_fd_sc_hd__nand2b_1 _13240_ (.A_N(_05199_),
    .B(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__xnor2_1 _13241_ (.A(_05198_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__o21bai_1 _13242_ (.A1(_05195_),
    .A2(_05197_),
    .B1_N(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__or3b_1 _13243_ (.A(_05195_),
    .B(_05197_),
    .C_N(_05202_),
    .X(_05204_));
 sky130_fd_sc_hd__o31a_1 _13244_ (.A1(_00192_),
    .A2(_02096_),
    .A3(_05083_),
    .B1(_05084_),
    .X(_05205_));
 sky130_fd_sc_hd__a21oi_1 _13245_ (.A1(_05203_),
    .A2(_05204_),
    .B1(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__o2111ai_2 _13246_ (.A1(_05068_),
    .A2(_05083_),
    .B1(_05084_),
    .C1(_05203_),
    .D1(_05204_),
    .Y(_05208_));
 sky130_fd_sc_hd__nand2b_1 _13247_ (.A_N(_05206_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__o21ai_2 _13248_ (.A1(_05089_),
    .A2(_05092_),
    .B1(_05090_),
    .Y(_05210_));
 sky130_fd_sc_hd__xor2_1 _13249_ (.A(_05209_),
    .B(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__xnor2_1 _13250_ (.A(_05209_),
    .B(_05210_),
    .Y(_05212_));
 sky130_fd_sc_hd__xor2_1 _13251_ (.A(_05176_),
    .B(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__a21oi_1 _13252_ (.A1(_05171_),
    .A2(_05172_),
    .B1(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__o21ai_1 _13253_ (.A1(_05176_),
    .A2(_05212_),
    .B1(_05173_),
    .Y(_05215_));
 sky130_fd_sc_hd__a21oi_1 _13254_ (.A1(_05176_),
    .A2(_05212_),
    .B1(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nor2_1 _13255_ (.A(_05214_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__nor2_1 _13256_ (.A(_05166_),
    .B(_05217_),
    .Y(_05219_));
 sky130_fd_sc_hd__o21ai_1 _13257_ (.A1(_05173_),
    .A2(_05213_),
    .B1(_05166_),
    .Y(_05220_));
 sky130_fd_sc_hd__o21ba_1 _13258_ (.A1(_05216_),
    .A2(_05220_),
    .B1_N(_05219_),
    .X(_05221_));
 sky130_fd_sc_hd__o2bb2ai_1 _13259_ (.A1_N(_05055_),
    .A2_N(_05108_),
    .B1(_05112_),
    .B2(_04871_),
    .Y(_05222_));
 sky130_fd_sc_hd__o21ai_2 _13260_ (.A1(_05055_),
    .A2(_05108_),
    .B1(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__xnor2_4 _13261_ (.A(_05221_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__o2bb2a_1 _13262_ (.A1_N(_05121_),
    .A2_N(_05123_),
    .B1(_01542_),
    .B2(_04880_),
    .X(_05225_));
 sky130_fd_sc_hd__o41a_1 _13263_ (.A1(_00744_),
    .A2(_01037_),
    .A3(_01221_),
    .A4(net136),
    .B1(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__nor2_1 _13264_ (.A(_05118_),
    .B(_05225_),
    .Y(_05227_));
 sky130_fd_sc_hd__o211a_1 _13265_ (.A1(_01181_),
    .A2(_01182_),
    .B1(_01218_),
    .C1(_01220_),
    .X(_05228_));
 sky130_fd_sc_hd__nand3_2 _13266_ (.A(_01659_),
    .B(net140),
    .C(_00569_),
    .Y(_05230_));
 sky130_fd_sc_hd__o21ai_2 _13267_ (.A1(_00903_),
    .A2(_01542_),
    .B1(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__o211ai_4 _13268_ (.A1(_00894_),
    .A2(_00896_),
    .B1(_01659_),
    .C1(net140),
    .Y(_05232_));
 sky130_fd_sc_hd__nand4_2 _13269_ (.A(_01659_),
    .B(_00569_),
    .C(_00904_),
    .D(net140),
    .Y(_05233_));
 sky130_fd_sc_hd__and3_1 _13270_ (.A(_00904_),
    .B(_01664_),
    .C(_05122_),
    .X(_05234_));
 sky130_fd_sc_hd__nand4_1 _13271_ (.A(_05122_),
    .B(net140),
    .C(_01659_),
    .D(_00904_),
    .Y(_05235_));
 sky130_fd_sc_hd__o2111ai_4 _13272_ (.A1(_05233_),
    .A2(_01542_),
    .B1(_01273_),
    .C1(_01059_),
    .D1(_05231_),
    .Y(_05236_));
 sky130_fd_sc_hd__a22oi_1 _13273_ (.A1(_01059_),
    .A2(_01273_),
    .B1(_05231_),
    .B2(_05235_),
    .Y(_05237_));
 sky130_fd_sc_hd__a32o_1 _13274_ (.A1(_01055_),
    .A2(_01057_),
    .A3(_01273_),
    .B1(_05231_),
    .B2(_05235_),
    .X(_05238_));
 sky130_fd_sc_hd__a22o_1 _13275_ (.A1(_01189_),
    .A2(_01222_),
    .B1(_05236_),
    .B2(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__nand4_2 _13276_ (.A(_01189_),
    .B(_01222_),
    .C(_05236_),
    .D(_05238_),
    .Y(_05240_));
 sky130_fd_sc_hd__a211o_1 _13277_ (.A1(_05239_),
    .A2(_05240_),
    .B1(_05226_),
    .C1(_05227_),
    .X(_05241_));
 sky130_fd_sc_hd__o211ai_2 _13278_ (.A1(_05226_),
    .A2(_05227_),
    .B1(_05239_),
    .C1(_05240_),
    .Y(_05242_));
 sky130_fd_sc_hd__a21bo_1 _13279_ (.A1(_04881_),
    .A2(_05129_),
    .B1_N(_05130_),
    .X(_05243_));
 sky130_fd_sc_hd__a21oi_1 _13280_ (.A1(_05241_),
    .A2(_05242_),
    .B1(_05243_),
    .Y(_05244_));
 sky130_fd_sc_hd__a21o_1 _13281_ (.A1(_05241_),
    .A2(_05242_),
    .B1(_05243_),
    .X(_05245_));
 sky130_fd_sc_hd__and3_2 _13282_ (.A(_05241_),
    .B(_05243_),
    .C(_05242_),
    .X(_05246_));
 sky130_fd_sc_hd__nand3_1 _13283_ (.A(_05241_),
    .B(_05242_),
    .C(_05243_),
    .Y(_05247_));
 sky130_fd_sc_hd__and3_1 _13284_ (.A(_00581_),
    .B(_01820_),
    .C(_01821_),
    .X(_05248_));
 sky130_fd_sc_hd__nand4_1 _13285_ (.A(_01038_),
    .B(_01590_),
    .C(net137),
    .D(_00743_),
    .Y(_05249_));
 sky130_fd_sc_hd__o32a_1 _13286_ (.A1(_01584_),
    .A2(_01586_),
    .A3(_00744_),
    .B1(_01037_),
    .B2(net136),
    .X(_05251_));
 sky130_fd_sc_hd__a31o_1 _13287_ (.A1(_05116_),
    .A2(_01590_),
    .A3(_01038_),
    .B1(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__xnor2_1 _13288_ (.A(_05248_),
    .B(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__xor2_1 _13289_ (.A(_05248_),
    .B(_05252_),
    .X(_05254_));
 sky130_fd_sc_hd__nand3_2 _13290_ (.A(_05245_),
    .B(_05247_),
    .C(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__o21ai_2 _13291_ (.A1(_05244_),
    .A2(_05246_),
    .B1(_05253_),
    .Y(_05256_));
 sky130_fd_sc_hd__or3b_2 _13292_ (.A(_00580_),
    .B(_01589_),
    .C_N(_05137_),
    .X(_05257_));
 sky130_fd_sc_hd__a22oi_4 _13293_ (.A1(_05255_),
    .A2(_05256_),
    .B1(_05257_),
    .B2(_05138_),
    .Y(_05258_));
 sky130_fd_sc_hd__and4_1 _13294_ (.A(_05138_),
    .B(_05255_),
    .C(_05256_),
    .D(_05257_),
    .X(_05259_));
 sky130_fd_sc_hd__nand4_1 _13295_ (.A(_05138_),
    .B(_05255_),
    .C(_05256_),
    .D(_05257_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand2_1 _13296_ (.A(_05115_),
    .B(_05145_),
    .Y(_05262_));
 sky130_fd_sc_hd__a21o_1 _13297_ (.A1(_05141_),
    .A2(_05144_),
    .B1(_05115_),
    .X(_05263_));
 sky130_fd_sc_hd__o221a_2 _13298_ (.A1(_05141_),
    .A2(_05144_),
    .B1(_05258_),
    .B2(_05259_),
    .C1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__a211oi_4 _13299_ (.A1(_05145_),
    .A2(_05263_),
    .B1(_05259_),
    .C1(_05258_),
    .Y(_05265_));
 sky130_fd_sc_hd__or2_1 _13300_ (.A(_05264_),
    .B(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__or3_1 _13301_ (.A(_05264_),
    .B(_05265_),
    .C(_05224_),
    .X(_05267_));
 sky130_fd_sc_hd__o21ai_1 _13302_ (.A1(_05264_),
    .A2(_05265_),
    .B1(_05224_),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _13303_ (.A(_05267_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__a2111oi_4 _13304_ (.A1(_04726_),
    .A2(_03911_),
    .B1(_04903_),
    .C1(_05040_),
    .D1(_05044_),
    .Y(_05270_));
 sky130_fd_sc_hd__o31a_1 _13305_ (.A1(_05425_),
    .A2(_03449_),
    .A3(_05005_),
    .B1(_05004_),
    .X(_05271_));
 sky130_fd_sc_hd__a41o_1 _13306_ (.A1(_04939_),
    .A2(_04997_),
    .A3(_07513_),
    .A4(_02356_),
    .B1(_04998_),
    .X(_05273_));
 sky130_fd_sc_hd__o31ai_1 _13307_ (.A1(_07512_),
    .A2(_02632_),
    .A3(_04992_),
    .B1(_04991_),
    .Y(_05274_));
 sky130_fd_sc_hd__or4b_1 _13308_ (.A(net152),
    .B(_03179_),
    .C(_04938_),
    .D_N(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__a41o_1 _13309_ (.A1(_06341_),
    .A2(net151),
    .A3(_02858_),
    .A4(_03180_),
    .B1(_05274_),
    .X(_05276_));
 sky130_fd_sc_hd__or3_1 _13310_ (.A(_07508_),
    .B(_07510_),
    .C(_02857_),
    .X(_05277_));
 sky130_fd_sc_hd__a32o_1 _13311_ (.A1(_00275_),
    .A2(net139),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_00150_),
    .X(_05278_));
 sky130_fd_sc_hd__or4_2 _13312_ (.A(net144),
    .B(_00274_),
    .C(_02241_),
    .D(_02355_),
    .X(_05279_));
 sky130_fd_sc_hd__a22oi_2 _13313_ (.A1(_00010_),
    .A2(_02633_),
    .B1(_05278_),
    .B2(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__and4_1 _13314_ (.A(_00010_),
    .B(_02633_),
    .C(_05278_),
    .D(_05279_),
    .X(_05281_));
 sky130_fd_sc_hd__o21ai_1 _13315_ (.A1(_05280_),
    .A2(_05281_),
    .B1(_05277_),
    .Y(_05282_));
 sky130_fd_sc_hd__or4_1 _13316_ (.A(_07512_),
    .B(_02857_),
    .C(_05280_),
    .D(_05281_),
    .X(_05284_));
 sky130_fd_sc_hd__nand2_1 _13317_ (.A(_05282_),
    .B(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__a21oi_1 _13318_ (.A1(_05275_),
    .A2(_05276_),
    .B1(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__and3_1 _13319_ (.A(_05275_),
    .B(_05276_),
    .C(_05285_),
    .X(_05287_));
 sky130_fd_sc_hd__o21ai_1 _13320_ (.A1(_05286_),
    .A2(_05287_),
    .B1(_05273_),
    .Y(_05288_));
 sky130_fd_sc_hd__or3_1 _13321_ (.A(_05273_),
    .B(_05286_),
    .C(_05287_),
    .X(_05289_));
 sky130_fd_sc_hd__and3_2 _13322_ (.A(_05392_),
    .B(_05414_),
    .C(_03584_),
    .X(_05290_));
 sky130_fd_sc_hd__or3_1 _13323_ (.A(net152),
    .B(_03444_),
    .C(_03447_),
    .X(_05291_));
 sky130_fd_sc_hd__and4_1 _13324_ (.A(_06341_),
    .B(net151),
    .C(_03180_),
    .D(_03450_),
    .X(_05292_));
 sky130_fd_sc_hd__a32o_1 _13325_ (.A1(net151),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_03450_),
    .B2(_06341_),
    .X(_05293_));
 sky130_fd_sc_hd__o31a_1 _13326_ (.A1(_06331_),
    .A2(_03179_),
    .A3(_05291_),
    .B1(_05293_),
    .X(_05295_));
 sky130_fd_sc_hd__xor2_1 _13327_ (.A(_05290_),
    .B(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__a21oi_1 _13328_ (.A1(_05288_),
    .A2(_05289_),
    .B1(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__and3_1 _13329_ (.A(_05288_),
    .B(_05289_),
    .C(_05296_),
    .X(_05298_));
 sky130_fd_sc_hd__or2_1 _13330_ (.A(_05297_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__xor2_1 _13331_ (.A(_05271_),
    .B(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__nand2_1 _13332_ (.A(_05013_),
    .B(_05014_),
    .Y(_05301_));
 sky130_fd_sc_hd__nand2_1 _13333_ (.A(_05012_),
    .B(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__xor2_1 _13334_ (.A(_05300_),
    .B(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__o31a_2 _13335_ (.A1(_00274_),
    .A2(_02053_),
    .A3(_05020_),
    .B1(_05019_),
    .X(_05304_));
 sky130_fd_sc_hd__o31a_1 _13336_ (.A1(net142),
    .A2(_02049_),
    .A3(_02051_),
    .B1(_05304_),
    .X(_05306_));
 sky130_fd_sc_hd__a211oi_4 _13337_ (.A1(_00422_),
    .A2(_00423_),
    .B1(_02053_),
    .C1(_05304_),
    .Y(_05307_));
 sky130_fd_sc_hd__a21bo_1 _13338_ (.A1(_05027_),
    .A2(_05026_),
    .B1_N(_05025_),
    .X(_05308_));
 sky130_fd_sc_hd__nor3_1 _13339_ (.A(_05306_),
    .B(_05307_),
    .C(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__o21a_1 _13340_ (.A1(_05306_),
    .A2(_05307_),
    .B1(_05308_),
    .X(_05310_));
 sky130_fd_sc_hd__o21a_1 _13341_ (.A1(_05309_),
    .A2(_05310_),
    .B1(_05303_),
    .X(_05311_));
 sky130_fd_sc_hd__or3_1 _13342_ (.A(_05303_),
    .B(_05309_),
    .C(_05310_),
    .X(_05312_));
 sky130_fd_sc_hd__o21ai_1 _13343_ (.A1(_05270_),
    .A2(_05311_),
    .B1(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__inv_2 _13344_ (.A(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__a21o_1 _13345_ (.A1(_05270_),
    .A2(_05311_),
    .B1(_05313_),
    .X(_05315_));
 sky130_fd_sc_hd__o41a_1 _13346_ (.A1(_05270_),
    .A2(_05303_),
    .A3(_05309_),
    .A4(_05310_),
    .B1(_05315_),
    .X(_05317_));
 sky130_fd_sc_hd__a21oi_1 _13347_ (.A1(_05033_),
    .A2(_05046_),
    .B1(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand3b_1 _13348_ (.A_N(_05031_),
    .B(_05317_),
    .C(_05046_),
    .Y(_05319_));
 sky130_fd_sc_hd__and2b_1 _13349_ (.A_N(_05318_),
    .B(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__xnor2_1 _13350_ (.A(_05052_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__and2_1 _13351_ (.A(_05269_),
    .B(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__nor2_1 _13352_ (.A(_05269_),
    .B(_05321_),
    .Y(_05323_));
 sky130_fd_sc_hd__nor2_1 _13353_ (.A(_05322_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__a211oi_1 _13354_ (.A1(_05114_),
    .A2(_05148_),
    .B1(_05152_),
    .C1(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__a2bb2o_1 _13355_ (.A1_N(_05149_),
    .A2_N(_05152_),
    .B1(_05269_),
    .B2(_05321_),
    .X(_05326_));
 sky130_fd_sc_hd__o21a_1 _13356_ (.A1(_05149_),
    .A2(_05152_),
    .B1(_05324_),
    .X(_05328_));
 sky130_fd_sc_hd__o2bb2ai_1 _13357_ (.A1_N(_05155_),
    .A2_N(_05160_),
    .B1(_05325_),
    .B2(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__o311ai_4 _13358_ (.A1(_05149_),
    .A2(_05324_),
    .A3(_05152_),
    .B1(_05155_),
    .C1(_05160_),
    .Y(_05330_));
 sky130_fd_sc_hd__o21a_1 _13359_ (.A1(_05328_),
    .A2(_05330_),
    .B1(_05329_),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_1 _13360_ (.A1(_00845_),
    .A2(_05165_),
    .B1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__o221a_1 _13361_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_05161_),
    .B2(_04983_),
    .C1(_05331_),
    .X(_05333_));
 sky130_fd_sc_hd__nor2_1 _13362_ (.A(_05332_),
    .B(_05333_),
    .Y(net96));
 sky130_fd_sc_hd__nor2_1 _13363_ (.A(_05331_),
    .B(_05165_),
    .Y(_05334_));
 sky130_fd_sc_hd__o21ai_1 _13364_ (.A1(_05331_),
    .A2(_05165_),
    .B1(_00845_),
    .Y(_05335_));
 sky130_fd_sc_hd__o21a_1 _13365_ (.A1(_05175_),
    .A2(_05211_),
    .B1(_05215_),
    .X(_05336_));
 sky130_fd_sc_hd__a21oi_1 _13366_ (.A1(_05198_),
    .A2(_05200_),
    .B1(_05199_),
    .Y(_05338_));
 sky130_fd_sc_hd__a31o_1 _13367_ (.A1(_07540_),
    .A2(_02926_),
    .A3(_05190_),
    .B1(_05188_),
    .X(_05339_));
 sky130_fd_sc_hd__nor2_1 _13368_ (.A(_05338_),
    .B(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__a311o_1 _13369_ (.A1(_07540_),
    .A2(_02926_),
    .A3(_05190_),
    .B1(_05338_),
    .C1(_05188_),
    .X(_05341_));
 sky130_fd_sc_hd__nand2_1 _13370_ (.A(_05339_),
    .B(_05338_),
    .Y(_05342_));
 sky130_fd_sc_hd__o32a_1 _13371_ (.A1(net149),
    .A2(net132),
    .A3(net130),
    .B1(net148),
    .B2(_02925_),
    .X(_05343_));
 sky130_fd_sc_hd__and4_1 _13372_ (.A(_07540_),
    .B(_00072_),
    .C(_02926_),
    .D(_03087_),
    .X(_05344_));
 sky130_fd_sc_hd__or4_1 _13373_ (.A(_07189_),
    .B(_07441_),
    .C(_03319_),
    .D(_03652_),
    .X(_05345_));
 sky130_fd_sc_hd__a32o_1 _13374_ (.A1(_07200_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_03320_),
    .B2(_07440_),
    .X(_05346_));
 sky130_fd_sc_hd__o2bb2a_1 _13375_ (.A1_N(_05345_),
    .A2_N(_05346_),
    .B1(_05327_),
    .B2(_03832_),
    .X(_05347_));
 sky130_fd_sc_hd__o21ai_1 _13376_ (.A1(_05343_),
    .A2(_05344_),
    .B1(_05347_),
    .Y(_05349_));
 sky130_fd_sc_hd__or3_1 _13377_ (.A(_05343_),
    .B(_05344_),
    .C(_05347_),
    .X(_05350_));
 sky130_fd_sc_hd__a21oi_1 _13378_ (.A1(_05349_),
    .A2(_05350_),
    .B1(_05186_),
    .Y(_05351_));
 sky130_fd_sc_hd__and3_1 _13379_ (.A(_05350_),
    .B(_05186_),
    .C(_05349_),
    .X(_05352_));
 sky130_fd_sc_hd__or2_1 _13380_ (.A(_05351_),
    .B(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__and3_1 _13381_ (.A(_05341_),
    .B(_05342_),
    .C(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__a21oi_1 _13382_ (.A1(_05341_),
    .A2(_05342_),
    .B1(_05353_),
    .Y(_05355_));
 sky130_fd_sc_hd__or2_1 _13383_ (.A(_05354_),
    .B(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__inv_2 _13384_ (.A(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__a21oi_2 _13385_ (.A1(_05193_),
    .A2(_05180_),
    .B1(_05181_),
    .Y(_05358_));
 sky130_fd_sc_hd__xnor2_1 _13386_ (.A(_05356_),
    .B(_05358_),
    .Y(_05360_));
 sky130_fd_sc_hd__or3_1 _13387_ (.A(_00532_),
    .B(net133),
    .C(_02094_),
    .X(_05361_));
 sky130_fd_sc_hd__o32a_1 _13388_ (.A1(_00192_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_00366_),
    .B2(_02433_),
    .X(_05362_));
 sky130_fd_sc_hd__or4_1 _13389_ (.A(_00192_),
    .B(_00366_),
    .C(_02433_),
    .D(_02696_),
    .X(_05363_));
 sky130_fd_sc_hd__nand2b_1 _13390_ (.A_N(_05362_),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__xnor2_1 _13391_ (.A(_05361_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__xnor2_1 _13392_ (.A(_05360_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__o21bai_1 _13393_ (.A1(_05202_),
    .A2(_05195_),
    .B1_N(_05197_),
    .Y(_05367_));
 sky130_fd_sc_hd__and2_1 _13394_ (.A(_05366_),
    .B(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__nor2_1 _13395_ (.A(_05366_),
    .B(_05367_),
    .Y(_05369_));
 sky130_fd_sc_hd__a21oi_1 _13396_ (.A1(_05210_),
    .A2(_05208_),
    .B1(_05206_),
    .Y(_05371_));
 sky130_fd_sc_hd__o21ai_1 _13397_ (.A1(_05368_),
    .A2(_05369_),
    .B1(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__or3_1 _13398_ (.A(_05371_),
    .B(_05369_),
    .C(_05368_),
    .X(_05373_));
 sky130_fd_sc_hd__nand2_1 _13399_ (.A(_05372_),
    .B(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__a21boi_1 _13400_ (.A1(_05170_),
    .A2(_05168_),
    .B1_N(_05169_),
    .Y(_05375_));
 sky130_fd_sc_hd__xnor2_1 _13401_ (.A(_05374_),
    .B(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__nor2_1 _13402_ (.A(_05336_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__or2_1 _13403_ (.A(_05336_),
    .B(_05376_),
    .X(_05378_));
 sky130_fd_sc_hd__o211a_1 _13404_ (.A1(_05175_),
    .A2(_05211_),
    .B1(_05215_),
    .C1(_05376_),
    .X(_05379_));
 sky130_fd_sc_hd__or2_1 _13405_ (.A(_05377_),
    .B(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__o211ai_1 _13406_ (.A1(_05220_),
    .A2(_05216_),
    .B1(_05110_),
    .C1(_05222_),
    .Y(_05382_));
 sky130_fd_sc_hd__o21ai_2 _13407_ (.A1(_05166_),
    .A2(_05217_),
    .B1(_05382_),
    .Y(_05383_));
 sky130_fd_sc_hd__xnor2_2 _13408_ (.A(_05380_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__or4_2 _13409_ (.A(_00576_),
    .B(_00578_),
    .C(_02049_),
    .D(_02051_),
    .X(_05385_));
 sky130_fd_sc_hd__o32a_1 _13410_ (.A1(_01037_),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(_00744_),
    .X(_05386_));
 sky130_fd_sc_hd__or4_1 _13411_ (.A(_00744_),
    .B(_01037_),
    .C(_01589_),
    .D(_01822_),
    .X(_05387_));
 sky130_fd_sc_hd__nand2b_1 _13412_ (.A_N(_05386_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__xor2_2 _13413_ (.A(_05385_),
    .B(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__a21oi_1 _13414_ (.A1(_05239_),
    .A2(_05240_),
    .B1(_05227_),
    .Y(_05390_));
 sky130_fd_sc_hd__and3b_1 _13415_ (.A_N(_05226_),
    .B(_05239_),
    .C(_05240_),
    .X(_05391_));
 sky130_fd_sc_hd__o31a_1 _13416_ (.A1(_00580_),
    .A2(_01822_),
    .A3(_05251_),
    .B1(_05249_),
    .X(_05393_));
 sky130_fd_sc_hd__o31ai_1 _13417_ (.A1(_00580_),
    .A2(_01822_),
    .A3(_05251_),
    .B1(_05249_),
    .Y(_05394_));
 sky130_fd_sc_hd__o21ai_1 _13418_ (.A1(_01188_),
    .A2(_01221_),
    .B1(_05236_),
    .Y(_05395_));
 sky130_fd_sc_hd__and3_1 _13419_ (.A(_05238_),
    .B(_05394_),
    .C(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__nand3_1 _13420_ (.A(_05238_),
    .B(_05394_),
    .C(_05395_),
    .Y(_05397_));
 sky130_fd_sc_hd__o311ai_2 _13421_ (.A1(_01188_),
    .A2(_01221_),
    .A3(_05237_),
    .B1(_05393_),
    .C1(_05236_),
    .Y(_05398_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(_05397_),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__o32a_1 _13423_ (.A1(_01184_),
    .A2(_01186_),
    .A3(net136),
    .B1(_01272_),
    .B2(_01221_),
    .X(_05400_));
 sky130_fd_sc_hd__nand4_1 _13424_ (.A(_01189_),
    .B(_01222_),
    .C(_01273_),
    .D(net137),
    .Y(_05401_));
 sky130_fd_sc_hd__a31oi_1 _13425_ (.A1(_01273_),
    .A2(net137),
    .A3(_05228_),
    .B1(_05400_),
    .Y(_05402_));
 sky130_fd_sc_hd__a31o_1 _13426_ (.A1(_01273_),
    .A2(net137),
    .A3(_05228_),
    .B1(_05400_),
    .X(_05404_));
 sky130_fd_sc_hd__and3_1 _13427_ (.A(_01059_),
    .B(_01539_),
    .C(_01541_),
    .X(_05405_));
 sky130_fd_sc_hd__nand3_1 _13428_ (.A(net134),
    .B(_00569_),
    .C(_01879_),
    .Y(_05406_));
 sky130_fd_sc_hd__o21ai_2 _13429_ (.A1(_00903_),
    .A2(_01662_),
    .B1(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__o211ai_4 _13430_ (.A1(_00894_),
    .A2(_00896_),
    .B1(_01879_),
    .C1(net134),
    .Y(_05408_));
 sky130_fd_sc_hd__o2bb2ai_1 _13431_ (.A1_N(_05232_),
    .A2_N(_05406_),
    .B1(_05408_),
    .B2(_05230_),
    .Y(_05409_));
 sky130_fd_sc_hd__o21ai_1 _13432_ (.A1(_01058_),
    .A2(_01542_),
    .B1(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__o211ai_1 _13433_ (.A1(_05230_),
    .A2(_05408_),
    .B1(_05405_),
    .C1(_05407_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_1 _13434_ (.A(_05409_),
    .B(_05405_),
    .Y(_05412_));
 sky130_fd_sc_hd__o221ai_2 _13435_ (.A1(_01058_),
    .A2(_01542_),
    .B1(_05230_),
    .B2(_05408_),
    .C1(_05407_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand3_2 _13436_ (.A(_05404_),
    .B(_05412_),
    .C(_05413_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand3_1 _13437_ (.A(_05410_),
    .B(_05411_),
    .C(_05402_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21o_1 _13438_ (.A1(_05415_),
    .A2(_05416_),
    .B1(_05234_),
    .X(_05417_));
 sky130_fd_sc_hd__nand3_1 _13439_ (.A(_05415_),
    .B(_05416_),
    .C(_05234_),
    .Y(_05418_));
 sky130_fd_sc_hd__o21ai_1 _13440_ (.A1(_01542_),
    .A2(_05233_),
    .B1(_05416_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand3_1 _13441_ (.A(_05399_),
    .B(_05417_),
    .C(_05418_),
    .Y(_05420_));
 sky130_fd_sc_hd__a21o_1 _13442_ (.A1(_05417_),
    .A2(_05418_),
    .B1(_05399_),
    .X(_05421_));
 sky130_fd_sc_hd__a2bb2oi_2 _13443_ (.A1_N(_05227_),
    .A2_N(_05391_),
    .B1(_05420_),
    .B2(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__o211ai_2 _13444_ (.A1(_05226_),
    .A2(_05390_),
    .B1(_05420_),
    .C1(_05421_),
    .Y(_05423_));
 sky130_fd_sc_hd__or2_1 _13445_ (.A(_05389_),
    .B(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__a21o_1 _13446_ (.A1(_05423_),
    .A2(_05389_),
    .B1(_05422_),
    .X(_05426_));
 sky130_fd_sc_hd__a21oi_2 _13447_ (.A1(_05423_),
    .A2(_05389_),
    .B1(_05422_),
    .Y(_05427_));
 sky130_fd_sc_hd__a22oi_4 _13448_ (.A1(_05389_),
    .A2(_05422_),
    .B1(_05424_),
    .B2(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__nor2_1 _13449_ (.A(_05244_),
    .B(_05253_),
    .Y(_05429_));
 sky130_fd_sc_hd__a21oi_1 _13450_ (.A1(_05245_),
    .A2(_05254_),
    .B1(_05246_),
    .Y(_05430_));
 sky130_fd_sc_hd__o21a_1 _13451_ (.A1(_05246_),
    .A2(_05429_),
    .B1(_05428_),
    .X(_05431_));
 sky130_fd_sc_hd__xor2_1 _13452_ (.A(_05428_),
    .B(_05430_),
    .X(_05432_));
 sky130_fd_sc_hd__a31oi_4 _13453_ (.A1(_05146_),
    .A2(_05260_),
    .A3(_05262_),
    .B1(_05258_),
    .Y(_05433_));
 sky130_fd_sc_hd__xnor2_2 _13454_ (.A(_05432_),
    .B(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__or2_1 _13455_ (.A(_05434_),
    .B(_05384_),
    .X(_05435_));
 sky130_fd_sc_hd__nand2_1 _13456_ (.A(_05384_),
    .B(_05434_),
    .Y(_05437_));
 sky130_fd_sc_hd__nand2_1 _13457_ (.A(_05435_),
    .B(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__o211a_2 _13458_ (.A1(_00299_),
    .A2(_07366_),
    .B1(_07368_),
    .C1(_03584_),
    .X(_05439_));
 sky130_fd_sc_hd__o32a_1 _13459_ (.A1(_06331_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(net152),
    .B2(_03449_),
    .X(_05440_));
 sky130_fd_sc_hd__a31o_1 _13460_ (.A1(_05439_),
    .A2(_03450_),
    .A3(_06341_),
    .B1(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__o31a_1 _13461_ (.A1(_05381_),
    .A2(_05403_),
    .A3(_03912_),
    .B1(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__o21bai_2 _13462_ (.A1(_05277_),
    .A2(_05280_),
    .B1_N(_05281_),
    .Y(_05443_));
 sky130_fd_sc_hd__a311oi_2 _13463_ (.A1(_05436_),
    .A2(_03584_),
    .A3(_05293_),
    .B1(_05443_),
    .C1(_05292_),
    .Y(_05444_));
 sky130_fd_sc_hd__o211ai_2 _13464_ (.A1(_05290_),
    .A2(_05292_),
    .B1(_05293_),
    .C1(_05443_),
    .Y(_05445_));
 sky130_fd_sc_hd__and2b_1 _13465_ (.A_N(_05444_),
    .B(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__a32o_1 _13466_ (.A1(_07513_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_00010_),
    .B2(_02858_),
    .X(_05448_));
 sky130_fd_sc_hd__or4_1 _13467_ (.A(_07512_),
    .B(_00009_),
    .C(_02857_),
    .D(_03179_),
    .X(_05449_));
 sky130_fd_sc_hd__o31a_1 _13468_ (.A1(_00009_),
    .A2(_03179_),
    .A3(_05277_),
    .B1(_05448_),
    .X(_05450_));
 sky130_fd_sc_hd__o221a_1 _13469_ (.A1(_00299_),
    .A2(_00424_),
    .B1(_02350_),
    .B2(_02351_),
    .C1(_00427_),
    .X(_05451_));
 sky130_fd_sc_hd__or4_1 _13470_ (.A(_00274_),
    .B(net142),
    .C(_02241_),
    .D(_02355_),
    .X(_05452_));
 sky130_fd_sc_hd__o32a_1 _13471_ (.A1(_00274_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(net142),
    .B2(_02241_),
    .X(_05453_));
 sky130_fd_sc_hd__a31o_1 _13472_ (.A1(_02240_),
    .A2(_05451_),
    .A3(_00275_),
    .B1(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__o21ai_1 _13473_ (.A1(net144),
    .A2(_02632_),
    .B1(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__or4_1 _13474_ (.A(_00145_),
    .B(_00147_),
    .C(_02632_),
    .D(_05454_),
    .X(_05456_));
 sky130_fd_sc_hd__and2_1 _13475_ (.A(_05455_),
    .B(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__xnor2_1 _13476_ (.A(_05450_),
    .B(_05457_),
    .Y(_05459_));
 sky130_fd_sc_hd__xnor2_2 _13477_ (.A(_05279_),
    .B(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__xnor2_1 _13478_ (.A(_05446_),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand2_1 _13479_ (.A(_05275_),
    .B(_05285_),
    .Y(_05462_));
 sky130_fd_sc_hd__a21oi_1 _13480_ (.A1(_05276_),
    .A2(_05462_),
    .B1(_05461_),
    .Y(_05463_));
 sky130_fd_sc_hd__nand3_1 _13481_ (.A(_05461_),
    .B(_05462_),
    .C(_05276_),
    .Y(_05464_));
 sky130_fd_sc_hd__nor2_1 _13482_ (.A(_05442_),
    .B(_05463_),
    .Y(_05465_));
 sky130_fd_sc_hd__a31o_1 _13483_ (.A1(_05276_),
    .A2(_05461_),
    .A3(_05462_),
    .B1(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__or2_1 _13484_ (.A(_05463_),
    .B(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__a22oi_1 _13485_ (.A1(_05464_),
    .A2(_05465_),
    .B1(_05467_),
    .B2(_05442_),
    .Y(_05468_));
 sky130_fd_sc_hd__a21bo_1 _13486_ (.A1(_05289_),
    .A2(_05296_),
    .B1_N(_05288_),
    .X(_05470_));
 sky130_fd_sc_hd__nor2_1 _13487_ (.A(_05468_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__nand2_1 _13488_ (.A(_05468_),
    .B(_05470_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2b_1 _13489_ (.A_N(_05471_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__o2bb2a_1 _13490_ (.A1_N(_05012_),
    .A2_N(_05301_),
    .B1(_05299_),
    .B2(_05271_),
    .X(_05474_));
 sky130_fd_sc_hd__a21o_1 _13491_ (.A1(_05271_),
    .A2(_05299_),
    .B1(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__xnor2_1 _13492_ (.A(_05473_),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__o21ba_1 _13493_ (.A1(_05306_),
    .A2(_05308_),
    .B1_N(_05307_),
    .X(_05477_));
 sky130_fd_sc_hd__xnor2_1 _13494_ (.A(_05476_),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__nor2_1 _13495_ (.A(_05314_),
    .B(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_1 _13496_ (.A(_05314_),
    .B(_05478_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand2b_1 _13497_ (.A_N(_05479_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__a31o_1 _13498_ (.A1(_05049_),
    .A2(_05050_),
    .A3(_05319_),
    .B1(_05318_),
    .X(_05483_));
 sky130_fd_sc_hd__xor2_2 _13499_ (.A(_05482_),
    .B(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__xnor2_2 _13500_ (.A(_05438_),
    .B(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__a21oi_1 _13501_ (.A1(_05224_),
    .A2(_05266_),
    .B1(_05321_),
    .Y(_05486_));
 sky130_fd_sc_hd__inv_2 _13502_ (.A(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__a21o_1 _13503_ (.A1(_05267_),
    .A2(_05487_),
    .B1(_05485_),
    .X(_05488_));
 sky130_fd_sc_hd__o211ai_4 _13504_ (.A1(_05224_),
    .A2(_05266_),
    .B1(_05487_),
    .C1(_05485_),
    .Y(_05489_));
 sky130_fd_sc_hd__nand2_1 _13505_ (.A(_05488_),
    .B(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__o21a_1 _13506_ (.A1(_05323_),
    .A2(_05326_),
    .B1(_05330_),
    .X(_05492_));
 sky130_fd_sc_hd__o211ai_4 _13507_ (.A1(_05326_),
    .A2(_05323_),
    .B1(_05488_),
    .C1(_05330_),
    .Y(_05493_));
 sky130_fd_sc_hd__xnor2_2 _13508_ (.A(_05490_),
    .B(_05492_),
    .Y(_05494_));
 sky130_fd_sc_hd__xor2_1 _13509_ (.A(_05335_),
    .B(_05494_),
    .X(net97));
 sky130_fd_sc_hd__a2bb2o_1 _13510_ (.A1_N(_00812_),
    .A2_N(_00823_),
    .B1(_05334_),
    .B2(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__a21boi_2 _13511_ (.A1(_05435_),
    .A2(_05484_),
    .B1_N(_05437_),
    .Y(_05496_));
 sky130_fd_sc_hd__and3_1 _13512_ (.A(_00581_),
    .B(net139),
    .C(_02237_),
    .X(_05497_));
 sky130_fd_sc_hd__a21oi_1 _13513_ (.A1(_05385_),
    .A2(_05387_),
    .B1(_05386_),
    .Y(_05498_));
 sky130_fd_sc_hd__a21oi_1 _13514_ (.A1(_05415_),
    .A2(_05419_),
    .B1(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__a21o_1 _13515_ (.A1(_05415_),
    .A2(_05419_),
    .B1(_05498_),
    .X(_05500_));
 sky130_fd_sc_hd__nand3_1 _13516_ (.A(_05415_),
    .B(_05419_),
    .C(_05498_),
    .Y(_05502_));
 sky130_fd_sc_hd__a32o_1 _13517_ (.A1(net137),
    .A2(_01271_),
    .A3(_01269_),
    .B1(_01189_),
    .B2(_01590_),
    .X(_05503_));
 sky130_fd_sc_hd__nand4_2 _13518_ (.A(net137),
    .B(_01590_),
    .C(_01189_),
    .D(_01273_),
    .Y(_05504_));
 sky130_fd_sc_hd__and2_1 _13519_ (.A(_05503_),
    .B(_05504_),
    .X(_05505_));
 sky130_fd_sc_hd__and3_2 _13520_ (.A(_01222_),
    .B(_01539_),
    .C(_01541_),
    .X(_05506_));
 sky130_fd_sc_hd__o32a_1 _13521_ (.A1(_01058_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_01882_),
    .B2(_00903_),
    .X(_05507_));
 sky130_fd_sc_hd__a32o_2 _13522_ (.A1(_00904_),
    .A2(_01879_),
    .A3(net134),
    .B1(_01059_),
    .B2(_01664_),
    .X(_05508_));
 sky130_fd_sc_hd__o21ai_4 _13523_ (.A1(net48),
    .A2(_01877_),
    .B1(_01059_),
    .Y(_05509_));
 sky130_fd_sc_hd__nor4_2 _13524_ (.A(_00903_),
    .B(_01058_),
    .C(_01662_),
    .D(_01882_),
    .Y(_05510_));
 sky130_fd_sc_hd__o22ai_4 _13525_ (.A1(_01221_),
    .A2(_01542_),
    .B1(_05507_),
    .B2(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__o311ai_4 _13526_ (.A1(_05509_),
    .A2(_01878_),
    .A3(_05232_),
    .B1(_05506_),
    .C1(_05508_),
    .Y(_05513_));
 sky130_fd_sc_hd__and3_1 _13527_ (.A(_05511_),
    .B(_05513_),
    .C(_05505_),
    .X(_05514_));
 sky130_fd_sc_hd__a21oi_1 _13528_ (.A1(_05511_),
    .A2(_05513_),
    .B1(_05505_),
    .Y(_05515_));
 sky130_fd_sc_hd__a22o_1 _13529_ (.A1(_05503_),
    .A2(_05504_),
    .B1(_05511_),
    .B2(_05513_),
    .X(_05516_));
 sky130_fd_sc_hd__o22ai_1 _13530_ (.A1(_01058_),
    .A2(_01542_),
    .B1(_05230_),
    .B2(_05408_),
    .Y(_05517_));
 sky130_fd_sc_hd__and2_1 _13531_ (.A(_05407_),
    .B(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__o21ai_2 _13532_ (.A1(_05514_),
    .A2(_05515_),
    .B1(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__a211o_1 _13533_ (.A1(_05407_),
    .A2(_05517_),
    .B1(_05515_),
    .C1(_05514_),
    .X(_05520_));
 sky130_fd_sc_hd__nand4_1 _13534_ (.A(_05500_),
    .B(_05502_),
    .C(_05519_),
    .D(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__a22o_1 _13535_ (.A1(_05500_),
    .A2(_05502_),
    .B1(_05519_),
    .B2(_05520_),
    .X(_05522_));
 sky130_fd_sc_hd__a31oi_1 _13536_ (.A1(_05398_),
    .A2(_05417_),
    .A3(_05418_),
    .B1(_05396_),
    .Y(_05524_));
 sky130_fd_sc_hd__nand3_1 _13537_ (.A(_05521_),
    .B(_05522_),
    .C(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__a21o_1 _13538_ (.A1(_05521_),
    .A2(_05522_),
    .B1(_05524_),
    .X(_05526_));
 sky130_fd_sc_hd__o21ai_1 _13539_ (.A1(_01037_),
    .A2(_01822_),
    .B1(_05401_),
    .Y(_05527_));
 sky130_fd_sc_hd__and4b_1 _13540_ (.A_N(_05401_),
    .B(_01821_),
    .C(_01820_),
    .D(_01038_),
    .X(_05528_));
 sky130_fd_sc_hd__or4_1 _13541_ (.A(_01033_),
    .B(_01035_),
    .C(_01822_),
    .D(_05401_),
    .X(_05529_));
 sky130_fd_sc_hd__o2bb2a_1 _13542_ (.A1_N(_05527_),
    .A2_N(_05529_),
    .B1(_00744_),
    .B2(_02053_),
    .X(_05530_));
 sky130_fd_sc_hd__and4_1 _13543_ (.A(_02054_),
    .B(_05527_),
    .C(_05529_),
    .D(_00743_),
    .X(_05531_));
 sky130_fd_sc_hd__nor2_1 _13544_ (.A(_05530_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__a21oi_1 _13545_ (.A1(_05525_),
    .A2(_05526_),
    .B1(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__and3_1 _13546_ (.A(_05525_),
    .B(_05526_),
    .C(_05532_),
    .X(_05535_));
 sky130_fd_sc_hd__nor2_1 _13547_ (.A(_05533_),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__xor2_2 _13548_ (.A(_05426_),
    .B(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__o32ai_4 _13549_ (.A1(_05246_),
    .A2(_05428_),
    .A3(_05429_),
    .B1(_05431_),
    .B2(_05433_),
    .Y(_05538_));
 sky130_fd_sc_hd__xnor2_4 _13550_ (.A(_05537_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__and3_1 _13551_ (.A(_02095_),
    .B(_00569_),
    .C(_02093_),
    .X(_05540_));
 sky130_fd_sc_hd__a2111oi_4 _13552_ (.A1(_00567_),
    .A2(_00568_),
    .B1(net133),
    .C1(_02094_),
    .D1(_05539_),
    .Y(_05541_));
 sky130_fd_sc_hd__o21ai_2 _13553_ (.A1(_00570_),
    .A2(_02096_),
    .B1(_05539_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand2b_1 _13554_ (.A_N(_05541_),
    .B(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__xnor2_1 _13555_ (.A(_05497_),
    .B(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__a21o_1 _13556_ (.A1(_05357_),
    .A2(_05358_),
    .B1(_05365_),
    .X(_05546_));
 sky130_fd_sc_hd__o21a_1 _13557_ (.A1(_05357_),
    .A2(_05358_),
    .B1(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__o21a_1 _13558_ (.A1(_05340_),
    .A2(_05353_),
    .B1(_05342_),
    .X(_05548_));
 sky130_fd_sc_hd__a21boi_2 _13559_ (.A1(_05186_),
    .A2(_05349_),
    .B1_N(_05350_),
    .Y(_05549_));
 sky130_fd_sc_hd__a211oi_2 _13560_ (.A1(_05361_),
    .A2(_05363_),
    .B1(_05362_),
    .C1(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__o311a_1 _13561_ (.A1(_00532_),
    .A2(_02096_),
    .A3(_05362_),
    .B1(_05363_),
    .C1(_05549_),
    .X(_05551_));
 sky130_fd_sc_hd__and3_1 _13562_ (.A(_00193_),
    .B(_02922_),
    .C(_02924_),
    .X(_05552_));
 sky130_fd_sc_hd__o32a_1 _13563_ (.A1(net148),
    .A2(net131),
    .A3(net130),
    .B1(_00192_),
    .B2(_02925_),
    .X(_05553_));
 sky130_fd_sc_hd__and3_1 _13564_ (.A(_05552_),
    .B(_03087_),
    .C(_00072_),
    .X(_05554_));
 sky130_fd_sc_hd__and3_1 _13565_ (.A(_07540_),
    .B(_03316_),
    .C(_03318_),
    .X(_05555_));
 sky130_fd_sc_hd__o22a_1 _13566_ (.A1(net149),
    .A2(_03319_),
    .B1(_07441_),
    .B2(_03652_),
    .X(_05557_));
 sky130_fd_sc_hd__and3_1 _13567_ (.A(_07440_),
    .B(_05555_),
    .C(_03653_),
    .X(_05558_));
 sky130_fd_sc_hd__o32a_1 _13568_ (.A1(_07146_),
    .A2(_07168_),
    .A3(_03832_),
    .B1(_05557_),
    .B2(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__or3_1 _13569_ (.A(_05553_),
    .B(_05554_),
    .C(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__o21ai_1 _13570_ (.A1(_05553_),
    .A2(_05554_),
    .B1(_05559_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand2_1 _13571_ (.A(_05560_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__or4b_1 _13572_ (.A(_07441_),
    .B(_03319_),
    .C(_05184_),
    .D_N(_05561_),
    .X(_05563_));
 sky130_fd_sc_hd__xnor2_1 _13573_ (.A(_05345_),
    .B(_05562_),
    .Y(_05564_));
 sky130_fd_sc_hd__o21ai_1 _13574_ (.A1(_05550_),
    .A2(_05551_),
    .B1(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__or3_1 _13575_ (.A(_05550_),
    .B(_05551_),
    .C(_05564_),
    .X(_05566_));
 sky130_fd_sc_hd__and2_1 _13576_ (.A(_05565_),
    .B(_05566_),
    .X(_05568_));
 sky130_fd_sc_hd__and2b_1 _13577_ (.A_N(_05548_),
    .B(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__nand2b_1 _13578_ (.A_N(_05568_),
    .B(_05548_),
    .Y(_05570_));
 sky130_fd_sc_hd__and2b_1 _13579_ (.A_N(_05569_),
    .B(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__a221o_1 _13580_ (.A1(net25),
    .A2(_00530_),
    .B1(_02430_),
    .B2(_02431_),
    .C1(_00527_),
    .X(_05572_));
 sky130_fd_sc_hd__and3_1 _13581_ (.A(_05344_),
    .B(_02697_),
    .C(_00367_),
    .X(_05573_));
 sky130_fd_sc_hd__a21oi_1 _13582_ (.A1(_00367_),
    .A2(_02697_),
    .B1(_05344_),
    .Y(_05574_));
 sky130_fd_sc_hd__o2111ai_1 _13583_ (.A1(_05573_),
    .A2(_05574_),
    .B1(_00528_),
    .C1(_00531_),
    .D1(_02432_),
    .Y(_05575_));
 sky130_fd_sc_hd__a311o_1 _13584_ (.A1(_00528_),
    .A2(_00531_),
    .A3(_02432_),
    .B1(_05573_),
    .C1(_05574_),
    .X(_05576_));
 sky130_fd_sc_hd__nand2_1 _13585_ (.A(_05575_),
    .B(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__xnor2_1 _13586_ (.A(_05571_),
    .B(_05577_),
    .Y(_05579_));
 sky130_fd_sc_hd__xnor2_1 _13587_ (.A(_05547_),
    .B(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21bai_1 _13588_ (.A1(_05369_),
    .A2(_05371_),
    .B1_N(_05368_),
    .Y(_05581_));
 sky130_fd_sc_hd__xnor2_1 _13589_ (.A(_05580_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__inv_2 _13590_ (.A(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__o21a_1 _13591_ (.A1(_05374_),
    .A2(_05375_),
    .B1(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__or3_1 _13592_ (.A(_05374_),
    .B(_05375_),
    .C(_05583_),
    .X(_05585_));
 sky130_fd_sc_hd__nand2b_1 _13593_ (.A_N(_05584_),
    .B(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__o21a_1 _13594_ (.A1(_05379_),
    .A2(_05383_),
    .B1(_05378_),
    .X(_05587_));
 sky130_fd_sc_hd__xor2_2 _13595_ (.A(_05586_),
    .B(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__nor2_1 _13596_ (.A(_05544_),
    .B(_05588_),
    .Y(_05590_));
 sky130_fd_sc_hd__o21a_1 _13597_ (.A1(_05471_),
    .A2(_05475_),
    .B1(_05472_),
    .X(_05591_));
 sky130_fd_sc_hd__or2_1 _13598_ (.A(_05444_),
    .B(_05460_),
    .X(_05592_));
 sky130_fd_sc_hd__a21bo_1 _13599_ (.A1(_05450_),
    .A2(_05457_),
    .B1_N(_05279_),
    .X(_05593_));
 sky130_fd_sc_hd__o21a_1 _13600_ (.A1(_05450_),
    .A2(_05457_),
    .B1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__or4b_1 _13601_ (.A(_06331_),
    .B(_03583_),
    .C(_05291_),
    .D_N(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__a31oi_2 _13602_ (.A1(_06341_),
    .A2(_03450_),
    .A3(_05439_),
    .B1(_05594_),
    .Y(_05596_));
 sky130_fd_sc_hd__inv_2 _13603_ (.A(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__and3_1 _13604_ (.A(_07513_),
    .B(_03445_),
    .C(_03448_),
    .X(_05598_));
 sky130_fd_sc_hd__a31o_1 _13605_ (.A1(_00010_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_05598_),
    .X(_05599_));
 sky130_fd_sc_hd__or4_1 _13606_ (.A(_00005_),
    .B(_00007_),
    .C(_03444_),
    .D(_03447_),
    .X(_05601_));
 sky130_fd_sc_hd__or4_2 _13607_ (.A(_07512_),
    .B(_00009_),
    .C(_03179_),
    .D(_03449_),
    .X(_05602_));
 sky130_fd_sc_hd__and3_1 _13608_ (.A(_05451_),
    .B(_02633_),
    .C(_00275_),
    .X(_05603_));
 sky130_fd_sc_hd__o32a_1 _13609_ (.A1(_00274_),
    .A2(_02628_),
    .A3(_02630_),
    .B1(net142),
    .B2(_02355_),
    .X(_05604_));
 sky130_fd_sc_hd__a31o_1 _13610_ (.A1(_00271_),
    .A2(_00273_),
    .A3(_02633_),
    .B1(_05451_),
    .X(_05605_));
 sky130_fd_sc_hd__o211a_1 _13611_ (.A1(_05603_),
    .A2(_05604_),
    .B1(_00150_),
    .C1(_02858_),
    .X(_05606_));
 sky130_fd_sc_hd__a311oi_2 _13612_ (.A1(_00146_),
    .A2(_00148_),
    .A3(_02858_),
    .B1(_05603_),
    .C1(_05604_),
    .Y(_05607_));
 sky130_fd_sc_hd__a211oi_1 _13613_ (.A1(_05599_),
    .A2(_05602_),
    .B1(_05606_),
    .C1(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__a211o_1 _13614_ (.A1(_05599_),
    .A2(_05602_),
    .B1(_05606_),
    .C1(_05607_),
    .X(_05609_));
 sky130_fd_sc_hd__o211a_1 _13615_ (.A1(_05606_),
    .A2(_05607_),
    .B1(_05599_),
    .C1(_05602_),
    .X(_05610_));
 sky130_fd_sc_hd__o31ai_2 _13616_ (.A1(net144),
    .A2(_02632_),
    .A3(_05453_),
    .B1(_05452_),
    .Y(_05612_));
 sky130_fd_sc_hd__o21a_1 _13617_ (.A1(_05608_),
    .A2(_05610_),
    .B1(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__nor3_1 _13618_ (.A(_05608_),
    .B(_05612_),
    .C(_05610_),
    .Y(_05614_));
 sky130_fd_sc_hd__nor2_1 _13619_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__and3_1 _13620_ (.A(_05595_),
    .B(_05597_),
    .C(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__o2bb2a_1 _13621_ (.A1_N(_05595_),
    .A2_N(_05597_),
    .B1(_05613_),
    .B2(_05614_),
    .X(_05617_));
 sky130_fd_sc_hd__nor2_1 _13622_ (.A(_05616_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__a21o_1 _13623_ (.A1(_05445_),
    .A2(_05592_),
    .B1(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__o211ai_2 _13624_ (.A1(_05444_),
    .A2(_05460_),
    .B1(_05445_),
    .C1(_05618_),
    .Y(_05620_));
 sky130_fd_sc_hd__or4_1 _13625_ (.A(net152),
    .B(_03581_),
    .C(_03582_),
    .D(_05449_),
    .X(_05621_));
 sky130_fd_sc_hd__o21ai_1 _13626_ (.A1(net152),
    .A2(_03583_),
    .B1(_05449_),
    .Y(_05623_));
 sky130_fd_sc_hd__and3_1 _13627_ (.A(_03911_),
    .B(_06320_),
    .C(_06309_),
    .X(_05624_));
 sky130_fd_sc_hd__a21o_1 _13628_ (.A1(_05621_),
    .A2(_05623_),
    .B1(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__and3_1 _13629_ (.A(_05619_),
    .B(_05620_),
    .C(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a21oi_1 _13630_ (.A1(_05619_),
    .A2(_05620_),
    .B1(_05625_),
    .Y(_05627_));
 sky130_fd_sc_hd__nor2_1 _13631_ (.A(_05626_),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_1 _13632_ (.A(_05466_),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__nor3b_1 _13633_ (.A(_05466_),
    .B(_05628_),
    .C_N(_05591_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_1 _13634_ (.A(_05591_),
    .B(_05629_),
    .Y(_05631_));
 sky130_fd_sc_hd__o21a_1 _13635_ (.A1(_05466_),
    .A2(_05628_),
    .B1(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__o22ai_1 _13636_ (.A1(_05591_),
    .A2(_05629_),
    .B1(_05632_),
    .B2(_05630_),
    .Y(_05634_));
 sky130_fd_sc_hd__o21ba_1 _13637_ (.A1(_05476_),
    .A2(_05477_),
    .B1_N(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__or3b_1 _13638_ (.A(_05476_),
    .B(_05477_),
    .C_N(_05634_),
    .X(_05636_));
 sky130_fd_sc_hd__o21ai_2 _13639_ (.A1(_05479_),
    .A2(_05483_),
    .B1(_05481_),
    .Y(_05637_));
 sky130_fd_sc_hd__o21ai_2 _13640_ (.A1(_05635_),
    .A2(_05637_),
    .B1(_05636_),
    .Y(_05638_));
 sky130_fd_sc_hd__a21o_1 _13641_ (.A1(_05635_),
    .A2(_05637_),
    .B1(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__o21a_1 _13642_ (.A1(_05636_),
    .A2(_05637_),
    .B1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__and2_1 _13643_ (.A(_05544_),
    .B(_05588_),
    .X(_05641_));
 sky130_fd_sc_hd__o21ba_1 _13644_ (.A1(_05590_),
    .A2(_05640_),
    .B1_N(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__nor3_2 _13645_ (.A(_05590_),
    .B(_05640_),
    .C(_05641_),
    .Y(_05643_));
 sky130_fd_sc_hd__o21ai_1 _13646_ (.A1(_05590_),
    .A2(_05641_),
    .B1(_05640_),
    .Y(_05645_));
 sky130_fd_sc_hd__and2b_1 _13647_ (.A_N(_05643_),
    .B(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__or2_1 _13648_ (.A(_05496_),
    .B(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nand2_1 _13649_ (.A(_05496_),
    .B(_05645_),
    .Y(_05648_));
 sky130_fd_sc_hd__or2_1 _13650_ (.A(_05643_),
    .B(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__o2111ai_1 _13651_ (.A1(_05643_),
    .A2(_05648_),
    .B1(_05647_),
    .C1(_05489_),
    .D1(_05493_),
    .Y(_05650_));
 sky130_fd_sc_hd__a22o_1 _13652_ (.A1(_05489_),
    .A2(_05493_),
    .B1(_05647_),
    .B2(_05649_),
    .X(_05651_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(_05650_),
    .B(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__xor2_1 _13654_ (.A(_05495_),
    .B(_05652_),
    .X(net99));
 sky130_fd_sc_hd__and3_1 _13655_ (.A(_05334_),
    .B(_05494_),
    .C(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__nand2_1 _13656_ (.A(_05620_),
    .B(_05625_),
    .Y(_05655_));
 sky130_fd_sc_hd__o32a_1 _13657_ (.A1(_07512_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(_00009_),
    .B2(_03449_),
    .X(_05656_));
 sky130_fd_sc_hd__a31o_1 _13658_ (.A1(_00010_),
    .A2(_03584_),
    .A3(_05598_),
    .B1(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__o41a_1 _13659_ (.A1(_00321_),
    .A2(net24),
    .A3(_07369_),
    .A4(_03580_),
    .B1(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__o21a_1 _13660_ (.A1(_05596_),
    .A2(_05615_),
    .B1(_05595_),
    .X(_05659_));
 sky130_fd_sc_hd__a21oi_1 _13661_ (.A1(_05609_),
    .A2(_05612_),
    .B1(_05610_),
    .Y(_05660_));
 sky130_fd_sc_hd__or4_1 _13662_ (.A(net152),
    .B(_03583_),
    .C(_05449_),
    .D(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__nand2_1 _13663_ (.A(_05621_),
    .B(_05660_),
    .Y(_05662_));
 sky130_fd_sc_hd__o32a_1 _13664_ (.A1(net142),
    .A2(_02628_),
    .A3(_02630_),
    .B1(_02857_),
    .B2(_00274_),
    .X(_05663_));
 sky130_fd_sc_hd__and4_1 _13665_ (.A(_00275_),
    .B(_00429_),
    .C(_02633_),
    .D(_02858_),
    .X(_05664_));
 sky130_fd_sc_hd__o22ai_1 _13666_ (.A1(net144),
    .A2(_03179_),
    .B1(_05663_),
    .B2(_05664_),
    .Y(_05666_));
 sky130_fd_sc_hd__or4_1 _13667_ (.A(net144),
    .B(_03179_),
    .C(_05663_),
    .D(_05664_),
    .X(_05667_));
 sky130_fd_sc_hd__a31o_1 _13668_ (.A1(_00146_),
    .A2(_00148_),
    .A3(_02858_),
    .B1(_05603_),
    .X(_05668_));
 sky130_fd_sc_hd__a22oi_2 _13669_ (.A1(_05666_),
    .A2(_05667_),
    .B1(_05668_),
    .B2(_05605_),
    .Y(_05669_));
 sky130_fd_sc_hd__and4_1 _13670_ (.A(_05605_),
    .B(_05666_),
    .C(_05667_),
    .D(_05668_),
    .X(_05670_));
 sky130_fd_sc_hd__o21ai_1 _13671_ (.A1(_05669_),
    .A2(_05670_),
    .B1(_05602_),
    .Y(_05671_));
 sky130_fd_sc_hd__or3_1 _13672_ (.A(_05602_),
    .B(_05669_),
    .C(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__and2_1 _13673_ (.A(_05671_),
    .B(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__and3_1 _13674_ (.A(_05673_),
    .B(_05662_),
    .C(_05661_),
    .X(_05674_));
 sky130_fd_sc_hd__a21oi_1 _13675_ (.A1(_05661_),
    .A2(_05662_),
    .B1(_05673_),
    .Y(_05675_));
 sky130_fd_sc_hd__or2_1 _13676_ (.A(_05674_),
    .B(_05675_),
    .X(_05677_));
 sky130_fd_sc_hd__xor2_1 _13677_ (.A(_05659_),
    .B(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__xor2_1 _13678_ (.A(_05658_),
    .B(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__a21oi_1 _13679_ (.A1(_05619_),
    .A2(_05655_),
    .B1(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__nand3_1 _13680_ (.A(_05679_),
    .B(_05655_),
    .C(_05619_),
    .Y(_05681_));
 sky130_fd_sc_hd__or2_1 _13681_ (.A(_05632_),
    .B(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__a21oi_1 _13682_ (.A1(_05632_),
    .A2(_05681_),
    .B1(_05680_),
    .Y(_05683_));
 sky130_fd_sc_hd__a22o_1 _13683_ (.A1(_05632_),
    .A2(_05680_),
    .B1(_05682_),
    .B2(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__xnor2_1 _13684_ (.A(_05638_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__o21ai_2 _13685_ (.A1(_05584_),
    .A2(_05587_),
    .B1(_05585_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21ai_1 _13686_ (.A1(_05569_),
    .A2(_05577_),
    .B1(_05570_),
    .Y(_05688_));
 sky130_fd_sc_hd__nor2_1 _13687_ (.A(_05551_),
    .B(_05564_),
    .Y(_05689_));
 sky130_fd_sc_hd__o21ba_1 _13688_ (.A1(_05572_),
    .A2(_05574_),
    .B1_N(_05573_),
    .X(_05690_));
 sky130_fd_sc_hd__a21oi_1 _13689_ (.A1(_05560_),
    .A2(_05563_),
    .B1(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__a21o_1 _13690_ (.A1(_05560_),
    .A2(_05563_),
    .B1(_05690_),
    .X(_05692_));
 sky130_fd_sc_hd__and3_1 _13691_ (.A(_05560_),
    .B(_05563_),
    .C(_05690_),
    .X(_05693_));
 sky130_fd_sc_hd__a32o_1 _13692_ (.A1(_07540_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_00072_),
    .B2(_03320_),
    .X(_05694_));
 sky130_fd_sc_hd__or4_2 _13693_ (.A(net149),
    .B(net148),
    .C(_03319_),
    .D(_03652_),
    .X(_05695_));
 sky130_fd_sc_hd__o2bb2a_1 _13694_ (.A1_N(_05694_),
    .A2_N(_05695_),
    .B1(_07441_),
    .B2(_03832_),
    .X(_05696_));
 sky130_fd_sc_hd__o41a_1 _13695_ (.A1(_07441_),
    .A2(net149),
    .A3(_03319_),
    .A4(_03652_),
    .B1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__or4b_1 _13696_ (.A(_07441_),
    .B(_03652_),
    .C(_05696_),
    .D_N(_05555_),
    .X(_05699_));
 sky130_fd_sc_hd__and2b_1 _13697_ (.A_N(_05697_),
    .B(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__xnor2_1 _13698_ (.A(_05554_),
    .B(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__o21ai_1 _13699_ (.A1(_05691_),
    .A2(_05693_),
    .B1(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__or3_1 _13700_ (.A(_05691_),
    .B(_05693_),
    .C(_05701_),
    .X(_05703_));
 sky130_fd_sc_hd__nand2_1 _13701_ (.A(_05702_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21ba_1 _13702_ (.A1(_05550_),
    .A2(_05689_),
    .B1_N(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__or3b_1 _13703_ (.A(_05550_),
    .B(_05689_),
    .C_N(_05704_),
    .X(_05706_));
 sky130_fd_sc_hd__and2b_1 _13704_ (.A_N(_05705_),
    .B(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__or3_2 _13705_ (.A(_00532_),
    .B(_02692_),
    .C(_02694_),
    .X(_05708_));
 sky130_fd_sc_hd__o32a_1 _13706_ (.A1(_00192_),
    .A2(net131),
    .A3(net130),
    .B1(_00366_),
    .B2(_02925_),
    .X(_05710_));
 sky130_fd_sc_hd__a31o_1 _13707_ (.A1(_00367_),
    .A2(_03087_),
    .A3(_05552_),
    .B1(_05710_),
    .X(_05711_));
 sky130_fd_sc_hd__xor2_2 _13708_ (.A(_05708_),
    .B(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__xnor2_1 _13709_ (.A(_05707_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__or2_1 _13710_ (.A(_05688_),
    .B(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__nand2_1 _13711_ (.A(_05688_),
    .B(_05713_),
    .Y(_05715_));
 sky130_fd_sc_hd__o21ba_1 _13712_ (.A1(_05547_),
    .A2(_05579_),
    .B1_N(_05581_),
    .X(_05716_));
 sky130_fd_sc_hd__a21o_1 _13713_ (.A1(_05547_),
    .A2(_05579_),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__a21oi_1 _13714_ (.A1(_05714_),
    .A2(_05715_),
    .B1(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__and3_1 _13715_ (.A(_05714_),
    .B(_05715_),
    .C(_05717_),
    .X(_05719_));
 sky130_fd_sc_hd__or2_1 _13716_ (.A(_05718_),
    .B(_05719_),
    .X(_05721_));
 sky130_fd_sc_hd__nor2_1 _13717_ (.A(_05686_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__and2_1 _13718_ (.A(_05686_),
    .B(_05721_),
    .X(_05723_));
 sky130_fd_sc_hd__and3_1 _13719_ (.A(_00743_),
    .B(_05497_),
    .C(_02356_),
    .X(_05724_));
 sky130_fd_sc_hd__or4_1 _13720_ (.A(_00580_),
    .B(_00744_),
    .C(_02241_),
    .D(_02355_),
    .X(_05725_));
 sky130_fd_sc_hd__o32a_1 _13721_ (.A1(_00580_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_00744_),
    .B2(_02241_),
    .X(_05726_));
 sky130_fd_sc_hd__a31o_1 _13722_ (.A1(_00743_),
    .A2(_02356_),
    .A3(_05497_),
    .B1(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__and3_1 _13723_ (.A(_05540_),
    .B(_00904_),
    .C(_02432_),
    .X(_05728_));
 sky130_fd_sc_hd__o32a_1 _13724_ (.A1(_00903_),
    .A2(net133),
    .A3(_02094_),
    .B1(_02433_),
    .B2(_00570_),
    .X(_05729_));
 sky130_fd_sc_hd__a31oi_2 _13725_ (.A1(_05502_),
    .A2(_05519_),
    .A3(_05520_),
    .B1(_05499_),
    .Y(_05730_));
 sky130_fd_sc_hd__a31o_1 _13726_ (.A1(_00743_),
    .A2(_02054_),
    .A3(_05527_),
    .B1(_05528_),
    .X(_05732_));
 sky130_fd_sc_hd__a31oi_1 _13727_ (.A1(_05505_),
    .A2(_05511_),
    .A3(_05513_),
    .B1(_05518_),
    .Y(_05733_));
 sky130_fd_sc_hd__a31o_1 _13728_ (.A1(_05505_),
    .A2(_05511_),
    .A3(_05513_),
    .B1(_05518_),
    .X(_05734_));
 sky130_fd_sc_hd__nand3_1 _13729_ (.A(_05516_),
    .B(_05734_),
    .C(_05732_),
    .Y(_05735_));
 sky130_fd_sc_hd__a21oi_1 _13730_ (.A1(_05516_),
    .A2(_05734_),
    .B1(_05732_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21bai_1 _13731_ (.A1(_05515_),
    .A2(_05733_),
    .B1_N(_05732_),
    .Y(_05737_));
 sky130_fd_sc_hd__o32a_1 _13732_ (.A1(_01058_),
    .A2(_01662_),
    .A3(_05408_),
    .B1(_01221_),
    .B2(_01542_),
    .X(_05738_));
 sky130_fd_sc_hd__and3_1 _13733_ (.A(net137),
    .B(_01539_),
    .C(_01541_),
    .X(_05739_));
 sky130_fd_sc_hd__o22ai_4 _13734_ (.A1(_01878_),
    .A2(_05509_),
    .B1(_01221_),
    .B2(_01662_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand4b_2 _13735_ (.A_N(_05509_),
    .B(_01879_),
    .C(_01664_),
    .D(_01222_),
    .Y(_05741_));
 sky130_fd_sc_hd__o2bb2ai_2 _13736_ (.A1_N(_05740_),
    .A2_N(_05741_),
    .B1(net136),
    .B2(_01542_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand4_2 _13737_ (.A(_01544_),
    .B(_05740_),
    .C(_05741_),
    .D(net137),
    .Y(_05744_));
 sky130_fd_sc_hd__a2bb2o_1 _13738_ (.A1_N(_05507_),
    .A2_N(_05738_),
    .B1(_05743_),
    .B2(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__o2111ai_4 _13739_ (.A1(_05506_),
    .A2(_05510_),
    .B1(_05743_),
    .C1(_05744_),
    .D1(_05508_),
    .Y(_05746_));
 sky130_fd_sc_hd__nand2_1 _13740_ (.A(_05745_),
    .B(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__nand3b_1 _13741_ (.A_N(_05504_),
    .B(_05745_),
    .C(_05746_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand2_1 _13742_ (.A(_05504_),
    .B(_05747_),
    .Y(_05749_));
 sky130_fd_sc_hd__a41o_1 _13743_ (.A1(_01189_),
    .A2(_01273_),
    .A3(net137),
    .A4(_01590_),
    .B1(_05747_),
    .X(_05750_));
 sky130_fd_sc_hd__a21o_1 _13744_ (.A1(_05745_),
    .A2(_05746_),
    .B1(_05504_),
    .X(_05751_));
 sky130_fd_sc_hd__nand4_1 _13745_ (.A(_05735_),
    .B(_05737_),
    .C(_05748_),
    .D(_05749_),
    .Y(_05752_));
 sky130_fd_sc_hd__a22o_1 _13746_ (.A1(_05735_),
    .A2(_05737_),
    .B1(_05748_),
    .B2(_05749_),
    .X(_05754_));
 sky130_fd_sc_hd__a21o_1 _13747_ (.A1(_05752_),
    .A2(_05754_),
    .B1(_05730_),
    .X(_05755_));
 sky130_fd_sc_hd__nand3_1 _13748_ (.A(_05754_),
    .B(_05730_),
    .C(_05752_),
    .Y(_05756_));
 sky130_fd_sc_hd__nand2_1 _13749_ (.A(_05755_),
    .B(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__or4_1 _13750_ (.A(_01033_),
    .B(_01035_),
    .C(_02049_),
    .D(_02051_),
    .X(_05758_));
 sky130_fd_sc_hd__o32a_1 _13751_ (.A1(_01272_),
    .A2(_01584_),
    .A3(_01586_),
    .B1(_01822_),
    .B2(_01188_),
    .X(_05759_));
 sky130_fd_sc_hd__and4_1 _13752_ (.A(_01189_),
    .B(_01273_),
    .C(_01590_),
    .D(_01823_),
    .X(_05760_));
 sky130_fd_sc_hd__nor2_1 _13753_ (.A(_05759_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__xnor2_1 _13754_ (.A(_05758_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__xor2_1 _13755_ (.A(_05757_),
    .B(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__a21boi_1 _13756_ (.A1(_05525_),
    .A2(_05532_),
    .B1_N(_05526_),
    .Y(_05765_));
 sky130_fd_sc_hd__and2_1 _13757_ (.A(_05763_),
    .B(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__nor2_1 _13758_ (.A(_05763_),
    .B(_05765_),
    .Y(_05767_));
 sky130_fd_sc_hd__o21ai_1 _13759_ (.A1(_05426_),
    .A2(_05536_),
    .B1(_05538_),
    .Y(_05768_));
 sky130_fd_sc_hd__o31a_1 _13760_ (.A1(_05427_),
    .A2(_05533_),
    .A3(_05535_),
    .B1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__or3_1 _13761_ (.A(_05766_),
    .B(_05767_),
    .C(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__o21ai_1 _13762_ (.A1(_05766_),
    .A2(_05767_),
    .B1(_05769_),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _13763_ (.A(_05770_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__a311o_1 _13764_ (.A1(_00904_),
    .A2(_02432_),
    .A3(_05540_),
    .B1(_05729_),
    .C1(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__o21a_1 _13765_ (.A1(_05728_),
    .A2(_05729_),
    .B1(_05772_),
    .X(_05774_));
 sky130_fd_sc_hd__inv_2 _13766_ (.A(_05774_),
    .Y(_05776_));
 sky130_fd_sc_hd__a21oi_1 _13767_ (.A1(_05773_),
    .A2(_05776_),
    .B1(_05727_),
    .Y(_05777_));
 sky130_fd_sc_hd__and3_1 _13768_ (.A(_05727_),
    .B(_05773_),
    .C(_05776_),
    .X(_05778_));
 sky130_fd_sc_hd__nor2_1 _13769_ (.A(_05777_),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__inv_2 _13770_ (.A(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__o211ai_2 _13771_ (.A1(_05497_),
    .A2(_05541_),
    .B1(_05542_),
    .C1(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a311o_1 _13772_ (.A1(_00581_),
    .A2(_02240_),
    .A3(_05542_),
    .B1(_05541_),
    .C1(_05780_),
    .X(_05782_));
 sky130_fd_sc_hd__nand2_1 _13773_ (.A(_05781_),
    .B(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21ai_2 _13774_ (.A1(_05722_),
    .A2(_05723_),
    .B1(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__or3_1 _13775_ (.A(_05722_),
    .B(_05783_),
    .C(_05723_),
    .X(_05785_));
 sky130_fd_sc_hd__nand2_1 _13776_ (.A(_05784_),
    .B(_05785_),
    .Y(_05787_));
 sky130_fd_sc_hd__xor2_1 _13777_ (.A(_05685_),
    .B(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__inv_2 _13778_ (.A(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__or2_1 _13779_ (.A(_05642_),
    .B(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__nand2_2 _13780_ (.A(_05642_),
    .B(_05789_),
    .Y(_05791_));
 sky130_fd_sc_hd__nand2_1 _13781_ (.A(_05790_),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__o211ai_4 _13782_ (.A1(_05496_),
    .A2(_05646_),
    .B1(_05489_),
    .C1(_05493_),
    .Y(_05793_));
 sky130_fd_sc_hd__and3_1 _13783_ (.A(_05649_),
    .B(_05792_),
    .C(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__a21oi_1 _13784_ (.A1(_05649_),
    .A2(_05793_),
    .B1(_05792_),
    .Y(_05795_));
 sky130_fd_sc_hd__or2_1 _13785_ (.A(_05794_),
    .B(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__o21ai_1 _13786_ (.A1(_00834_),
    .A2(_05653_),
    .B1(_05796_),
    .Y(_05798_));
 sky130_fd_sc_hd__or4_1 _13787_ (.A(_00834_),
    .B(_05653_),
    .C(_05794_),
    .D(_05795_),
    .X(_05799_));
 sky130_fd_sc_hd__and2_1 _13788_ (.A(_05798_),
    .B(_05799_),
    .X(net100));
 sky130_fd_sc_hd__o2111a_1 _13789_ (.A1(_05794_),
    .A2(_05795_),
    .B1(_05652_),
    .C1(_05494_),
    .D1(_05334_),
    .X(_05800_));
 sky130_fd_sc_hd__o2bb2a_1 _13790_ (.A1_N(_05796_),
    .A2_N(_05653_),
    .B1(_00823_),
    .B2(_00812_),
    .X(_05801_));
 sky130_fd_sc_hd__nand2_1 _13791_ (.A(_05685_),
    .B(_05785_),
    .Y(_05802_));
 sky130_fd_sc_hd__nand2_2 _13792_ (.A(_05784_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__inv_2 _13793_ (.A(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__a21o_1 _13794_ (.A1(_05701_),
    .A2(_05692_),
    .B1(_05693_),
    .X(_05805_));
 sky130_fd_sc_hd__o41a_1 _13795_ (.A1(_00192_),
    .A2(_00366_),
    .A3(_02925_),
    .A4(_03086_),
    .B1(_05708_),
    .X(_05806_));
 sky130_fd_sc_hd__o41a_1 _13796_ (.A1(net148),
    .A2(_00192_),
    .A3(_02925_),
    .A4(_03086_),
    .B1(_05699_),
    .X(_05808_));
 sky130_fd_sc_hd__o22a_1 _13797_ (.A1(_05710_),
    .A2(_05806_),
    .B1(_05808_),
    .B2(_05697_),
    .X(_05809_));
 sky130_fd_sc_hd__nor4_1 _13798_ (.A(_05697_),
    .B(_05710_),
    .C(_05806_),
    .D(_05808_),
    .Y(_05810_));
 sky130_fd_sc_hd__nor2_1 _13799_ (.A(_05809_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__o32a_1 _13800_ (.A1(net148),
    .A2(_03652_),
    .A3(_05555_),
    .B1(_03832_),
    .B2(net149),
    .X(_05812_));
 sky130_fd_sc_hd__xor2_2 _13801_ (.A(_05811_),
    .B(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__nand2_1 _13802_ (.A(_05805_),
    .B(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__a211o_1 _13803_ (.A1(_05701_),
    .A2(_05692_),
    .B1(_05693_),
    .C1(_05813_),
    .X(_05815_));
 sky130_fd_sc_hd__or3_1 _13804_ (.A(_00532_),
    .B(_02920_),
    .C(_02923_),
    .X(_05816_));
 sky130_fd_sc_hd__and3_1 _13805_ (.A(_00367_),
    .B(_03316_),
    .C(_03318_),
    .X(_05817_));
 sky130_fd_sc_hd__or3_1 _13806_ (.A(_00361_),
    .B(_00363_),
    .C(_03319_),
    .X(_05819_));
 sky130_fd_sc_hd__o32a_1 _13807_ (.A1(_00366_),
    .A2(net132),
    .A3(net130),
    .B1(_03319_),
    .B2(_00192_),
    .X(_05820_));
 sky130_fd_sc_hd__a31o_1 _13808_ (.A1(_00193_),
    .A2(_03087_),
    .A3(_05817_),
    .B1(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__xnor2_1 _13809_ (.A(_05816_),
    .B(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__a21oi_1 _13810_ (.A1(_05814_),
    .A2(_05815_),
    .B1(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__and3_1 _13811_ (.A(_05814_),
    .B(_05815_),
    .C(_05822_),
    .X(_05824_));
 sky130_fd_sc_hd__a21oi_1 _13812_ (.A1(_05706_),
    .A2(_05712_),
    .B1(_05705_),
    .Y(_05825_));
 sky130_fd_sc_hd__o21ba_1 _13813_ (.A1(_05823_),
    .A2(_05824_),
    .B1_N(_05825_),
    .X(_05826_));
 sky130_fd_sc_hd__o21bai_1 _13814_ (.A1(_05823_),
    .A2(_05824_),
    .B1_N(_05825_),
    .Y(_05827_));
 sky130_fd_sc_hd__a2111oi_2 _13815_ (.A1(_05706_),
    .A2(_05712_),
    .B1(_05823_),
    .C1(_05824_),
    .D1(_05705_),
    .Y(_05828_));
 sky130_fd_sc_hd__nor2_1 _13816_ (.A(_05826_),
    .B(_05828_),
    .Y(_05830_));
 sky130_fd_sc_hd__a21bo_1 _13817_ (.A1(_05714_),
    .A2(_05717_),
    .B1_N(_05715_),
    .X(_05831_));
 sky130_fd_sc_hd__xnor2_2 _13818_ (.A(_05830_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__a21o_1 _13819_ (.A1(_05686_),
    .A2(_05721_),
    .B1(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__nand2_2 _13820_ (.A(_05723_),
    .B(_05832_),
    .Y(_05834_));
 sky130_fd_sc_hd__a31o_1 _13821_ (.A1(_05754_),
    .A2(_05730_),
    .A3(_05752_),
    .B1(_05762_),
    .X(_05835_));
 sky130_fd_sc_hd__nand2_1 _13822_ (.A(_05755_),
    .B(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__a31o_1 _13823_ (.A1(_05735_),
    .A2(_05750_),
    .A3(_05751_),
    .B1(_05736_),
    .X(_05837_));
 sky130_fd_sc_hd__nor2_1 _13824_ (.A(_05759_),
    .B(_05758_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_1 _13825_ (.A(_05504_),
    .B(_05746_),
    .Y(_05839_));
 sky130_fd_sc_hd__o211ai_2 _13826_ (.A1(_05760_),
    .A2(_05838_),
    .B1(_05839_),
    .C1(_05745_),
    .Y(_05841_));
 sky130_fd_sc_hd__a211o_1 _13827_ (.A1(_05745_),
    .A2(_05839_),
    .B1(_05838_),
    .C1(_05760_),
    .X(_05842_));
 sky130_fd_sc_hd__or4_1 _13828_ (.A(_01399_),
    .B(_01404_),
    .C(_01658_),
    .D(_01660_),
    .X(_05843_));
 sky130_fd_sc_hd__a22oi_1 _13829_ (.A1(_01059_),
    .A2(_01664_),
    .B1(_05740_),
    .B2(_05739_),
    .Y(_05844_));
 sky130_fd_sc_hd__a211oi_1 _13830_ (.A1(_01214_),
    .A2(_01215_),
    .B1(_01882_),
    .C1(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__a32o_1 _13831_ (.A1(_01222_),
    .A2(_01879_),
    .A3(net134),
    .B1(_05740_),
    .B2(_05739_),
    .X(_05846_));
 sky130_fd_sc_hd__o31ai_1 _13832_ (.A1(_01221_),
    .A2(_01882_),
    .A3(_05844_),
    .B1(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__xnor2_1 _13833_ (.A(_05843_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__a21boi_1 _13834_ (.A1(_05841_),
    .A2(_05842_),
    .B1_N(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__and3b_1 _13835_ (.A_N(_05848_),
    .B(_05842_),
    .C(_05841_),
    .X(_05850_));
 sky130_fd_sc_hd__o21a_1 _13836_ (.A1(_05849_),
    .A2(_05850_),
    .B1(_05837_),
    .X(_05852_));
 sky130_fd_sc_hd__or3_1 _13837_ (.A(_05837_),
    .B(_05849_),
    .C(_05850_),
    .X(_05853_));
 sky130_fd_sc_hd__nand2b_1 _13838_ (.A_N(_05852_),
    .B(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__and4_1 _13839_ (.A(_01273_),
    .B(_01544_),
    .C(_01590_),
    .D(_01823_),
    .X(_05855_));
 sky130_fd_sc_hd__or4_1 _13840_ (.A(_01272_),
    .B(_01542_),
    .C(_01589_),
    .D(_01822_),
    .X(_05856_));
 sky130_fd_sc_hd__a32o_1 _13841_ (.A1(_01273_),
    .A2(_01820_),
    .A3(_01821_),
    .B1(_01544_),
    .B2(_01590_),
    .X(_05857_));
 sky130_fd_sc_hd__a2111oi_1 _13842_ (.A1(_05856_),
    .A2(_05857_),
    .B1(_01184_),
    .C1(_01186_),
    .D1(_02053_),
    .Y(_05858_));
 sky130_fd_sc_hd__o311a_1 _13843_ (.A1(_01184_),
    .A2(_01186_),
    .A3(_02053_),
    .B1(_05856_),
    .C1(_05857_),
    .X(_05859_));
 sky130_fd_sc_hd__nor2_1 _13844_ (.A(_05858_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__and2_1 _13845_ (.A(_05854_),
    .B(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__nor2_1 _13846_ (.A(_05854_),
    .B(_05860_),
    .Y(_05863_));
 sky130_fd_sc_hd__o2bb2a_1 _13847_ (.A1_N(_05755_),
    .A2_N(_05835_),
    .B1(_05861_),
    .B2(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__nor3_1 _13848_ (.A(_05863_),
    .B(_05836_),
    .C(_05861_),
    .Y(_05865_));
 sky130_fd_sc_hd__nor2_1 _13849_ (.A(_05864_),
    .B(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__o21ba_1 _13850_ (.A1(_05766_),
    .A2(_05769_),
    .B1_N(_05767_),
    .X(_05867_));
 sky130_fd_sc_hd__xor2_2 _13851_ (.A(_05866_),
    .B(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__or3_1 _13852_ (.A(_00570_),
    .B(_02692_),
    .C(_02694_),
    .X(_05869_));
 sky130_fd_sc_hd__o32a_1 _13853_ (.A1(_00570_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_00903_),
    .B2(_02433_),
    .X(_05870_));
 sky130_fd_sc_hd__and4_1 _13854_ (.A(_00569_),
    .B(_02432_),
    .C(_02697_),
    .D(_00904_),
    .X(_05871_));
 sky130_fd_sc_hd__or4_1 _13855_ (.A(_01058_),
    .B(_02096_),
    .C(_05870_),
    .D(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__o22ai_1 _13856_ (.A1(_01058_),
    .A2(_02096_),
    .B1(_05870_),
    .B2(_05871_),
    .Y(_05874_));
 sky130_fd_sc_hd__a21oi_1 _13857_ (.A1(_05872_),
    .A2(_05874_),
    .B1(_05728_),
    .Y(_05875_));
 sky130_fd_sc_hd__and3_1 _13858_ (.A(_05872_),
    .B(_05874_),
    .C(_05728_),
    .X(_05876_));
 sky130_fd_sc_hd__or2_1 _13859_ (.A(_05875_),
    .B(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__xor2_1 _13860_ (.A(_05868_),
    .B(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__o32a_1 _13861_ (.A1(_00744_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_01037_),
    .B2(_02241_),
    .X(_05879_));
 sky130_fd_sc_hd__and4_1 _13862_ (.A(_00743_),
    .B(_02240_),
    .C(_02356_),
    .D(_01038_),
    .X(_05880_));
 sky130_fd_sc_hd__or4_1 _13863_ (.A(_00744_),
    .B(_01037_),
    .C(_02241_),
    .D(_02355_),
    .X(_05881_));
 sky130_fd_sc_hd__o32a_1 _13864_ (.A1(_00576_),
    .A2(_00578_),
    .A3(_02632_),
    .B1(_05879_),
    .B2(_05880_),
    .X(_05882_));
 sky130_fd_sc_hd__or4_1 _13865_ (.A(_00580_),
    .B(_02632_),
    .C(_05879_),
    .D(_05880_),
    .X(_05883_));
 sky130_fd_sc_hd__and2b_1 _13866_ (.A_N(_05882_),
    .B(_05883_),
    .X(_05885_));
 sky130_fd_sc_hd__xor2_1 _13867_ (.A(_05724_),
    .B(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__xnor2_1 _13868_ (.A(_05878_),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__o311a_1 _13869_ (.A1(_05724_),
    .A2(_05726_),
    .A3(_05774_),
    .B1(_05887_),
    .C1(_05773_),
    .X(_05888_));
 sky130_fd_sc_hd__a211o_1 _13870_ (.A1(_05727_),
    .A2(_05773_),
    .B1(_05774_),
    .C1(_05887_),
    .X(_05889_));
 sky130_fd_sc_hd__nand2b_1 _13871_ (.A_N(_05888_),
    .B(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__nand2_1 _13872_ (.A(_05781_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__or3b_1 _13873_ (.A(_05781_),
    .B(_05888_),
    .C_N(_05889_),
    .X(_05892_));
 sky130_fd_sc_hd__nand4_1 _13874_ (.A(_05833_),
    .B(_05834_),
    .C(_05891_),
    .D(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__a22oi_2 _13875_ (.A1(_05833_),
    .A2(_05834_),
    .B1(_05891_),
    .B2(_05892_),
    .Y(_05894_));
 sky130_fd_sc_hd__inv_2 _13876_ (.A(_05894_),
    .Y(_05896_));
 sky130_fd_sc_hd__nand2_1 _13877_ (.A(_05893_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__and3_1 _13878_ (.A(_00146_),
    .B(_00148_),
    .C(_03584_),
    .X(_05898_));
 sky130_fd_sc_hd__o32a_1 _13879_ (.A1(_00009_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(net144),
    .B2(_03449_),
    .X(_05899_));
 sky130_fd_sc_hd__a31o_1 _13880_ (.A1(_05898_),
    .A2(_03450_),
    .A3(_00010_),
    .B1(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__o31a_1 _13881_ (.A1(_07508_),
    .A2(_07510_),
    .A3(_03912_),
    .B1(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__and3_2 _13882_ (.A(_00275_),
    .B(_03176_),
    .C(_03178_),
    .X(_05902_));
 sky130_fd_sc_hd__o32a_1 _13883_ (.A1(net144),
    .A2(_03179_),
    .A3(_05663_),
    .B1(_00274_),
    .B2(_02632_),
    .X(_05903_));
 sky130_fd_sc_hd__or3_1 _13884_ (.A(net142),
    .B(_02857_),
    .C(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__o32ai_2 _13885_ (.A1(net144),
    .A2(_03179_),
    .A3(_05663_),
    .B1(net142),
    .B2(_02857_),
    .Y(_05905_));
 sky130_fd_sc_hd__a21oi_1 _13886_ (.A1(_05904_),
    .A2(_05905_),
    .B1(_05902_),
    .Y(_05907_));
 sky130_fd_sc_hd__o311a_1 _13887_ (.A1(net142),
    .A2(_02857_),
    .A3(_05903_),
    .B1(_05905_),
    .C1(_05902_),
    .X(_05908_));
 sky130_fd_sc_hd__nor2_1 _13888_ (.A(_05907_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__o21ba_1 _13889_ (.A1(_05602_),
    .A2(_05669_),
    .B1_N(_05670_),
    .X(_05910_));
 sky130_fd_sc_hd__and4b_1 _13890_ (.A_N(_05910_),
    .B(_03584_),
    .C(_00010_),
    .D(_05598_),
    .X(_05911_));
 sky130_fd_sc_hd__o31ai_1 _13891_ (.A1(_07512_),
    .A2(_03583_),
    .A3(_05601_),
    .B1(_05910_),
    .Y(_05912_));
 sky130_fd_sc_hd__and2b_1 _13892_ (.A_N(_05911_),
    .B(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__xor2_1 _13893_ (.A(_05909_),
    .B(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__a21bo_1 _13894_ (.A1(_05673_),
    .A2(_05662_),
    .B1_N(_05661_),
    .X(_05915_));
 sky130_fd_sc_hd__nor2_2 _13895_ (.A(_05914_),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_1 _13896_ (.A(_05914_),
    .B(_05915_),
    .Y(_05918_));
 sky130_fd_sc_hd__nor2_1 _13897_ (.A(_05901_),
    .B(_05916_),
    .Y(_05919_));
 sky130_fd_sc_hd__o311a_2 _13898_ (.A1(_07508_),
    .A2(_07510_),
    .A3(_03912_),
    .B1(_05900_),
    .C1(_05918_),
    .X(_05920_));
 sky130_fd_sc_hd__o21ai_1 _13899_ (.A1(_05914_),
    .A2(_05915_),
    .B1(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__a22o_1 _13900_ (.A1(_05918_),
    .A2(_05919_),
    .B1(_05921_),
    .B2(_05901_),
    .X(_05922_));
 sky130_fd_sc_hd__o21a_1 _13901_ (.A1(_05659_),
    .A2(_05677_),
    .B1(_05658_),
    .X(_05923_));
 sky130_fd_sc_hd__a21oi_1 _13902_ (.A1(_05659_),
    .A2(_05677_),
    .B1(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__and2b_1 _13903_ (.A_N(_05924_),
    .B(_05922_),
    .X(_05925_));
 sky130_fd_sc_hd__nand2b_1 _13904_ (.A_N(_05922_),
    .B(_05924_),
    .Y(_05926_));
 sky130_fd_sc_hd__nand2b_1 _13905_ (.A_N(_05925_),
    .B(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__xnor2_1 _13906_ (.A(_05683_),
    .B(_05927_),
    .Y(_05929_));
 sky130_fd_sc_hd__inv_2 _13907_ (.A(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand3_2 _13908_ (.A(_05638_),
    .B(_05684_),
    .C(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__a21o_1 _13909_ (.A1(_05638_),
    .A2(_05684_),
    .B1(_05930_),
    .X(_05932_));
 sky130_fd_sc_hd__nand2_1 _13910_ (.A(_05931_),
    .B(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__xnor2_2 _13911_ (.A(_05897_),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__inv_2 _13912_ (.A(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__or2_1 _13913_ (.A(_05803_),
    .B(_05934_),
    .X(_05936_));
 sky130_fd_sc_hd__a21o_1 _13914_ (.A1(_05784_),
    .A2(_05802_),
    .B1(_05935_),
    .X(_05937_));
 sky130_fd_sc_hd__o211ai_4 _13915_ (.A1(_05643_),
    .A2(_05648_),
    .B1(_05790_),
    .C1(_05793_),
    .Y(_05938_));
 sky130_fd_sc_hd__o211ai_4 _13916_ (.A1(_05935_),
    .A2(_05804_),
    .B1(_05791_),
    .C1(_05938_),
    .Y(_05940_));
 sky130_fd_sc_hd__and4_1 _13917_ (.A(_05791_),
    .B(_05936_),
    .C(_05937_),
    .D(_05938_),
    .X(_05941_));
 sky130_fd_sc_hd__a22oi_2 _13918_ (.A1(_05936_),
    .A2(_05937_),
    .B1(_05938_),
    .B2(_05791_),
    .Y(_05942_));
 sky130_fd_sc_hd__or2_1 _13919_ (.A(_05941_),
    .B(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__xnor2_1 _13920_ (.A(_05801_),
    .B(_05943_),
    .Y(net101));
 sky130_fd_sc_hd__o221a_1 _13921_ (.A1(_05794_),
    .A2(_05795_),
    .B1(_05941_),
    .B2(_05942_),
    .C1(_05653_),
    .X(_05944_));
 sky130_fd_sc_hd__o21a_1 _13922_ (.A1(_05805_),
    .A2(_05813_),
    .B1(_05822_),
    .X(_05945_));
 sky130_fd_sc_hd__a21o_1 _13923_ (.A1(_05805_),
    .A2(_05813_),
    .B1(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__a31o_1 _13924_ (.A1(_00193_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_05817_),
    .X(_05947_));
 sky130_fd_sc_hd__or4_2 _13925_ (.A(_00192_),
    .B(_00366_),
    .C(_03319_),
    .D(_03652_),
    .X(_05948_));
 sky130_fd_sc_hd__o2bb2a_1 _13926_ (.A1_N(_05947_),
    .A2_N(_05948_),
    .B1(net148),
    .B2(_03832_),
    .X(_05950_));
 sky130_fd_sc_hd__o32a_1 _13927_ (.A1(_00192_),
    .A2(_03086_),
    .A3(_05819_),
    .B1(_05820_),
    .B2(_05816_),
    .X(_05951_));
 sky130_fd_sc_hd__o21a_1 _13928_ (.A1(_05695_),
    .A2(_05951_),
    .B1(_05950_),
    .X(_05952_));
 sky130_fd_sc_hd__a21oi_2 _13929_ (.A1(_05695_),
    .A2(_05951_),
    .B1(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__a31o_1 _13930_ (.A1(_05695_),
    .A2(_05950_),
    .A3(_05951_),
    .B1(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__o31a_1 _13931_ (.A1(_05695_),
    .A2(_05950_),
    .A3(_05951_),
    .B1(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__o21ba_1 _13932_ (.A1(_05809_),
    .A2(_05812_),
    .B1_N(_05810_),
    .X(_05956_));
 sky130_fd_sc_hd__nand2_1 _13933_ (.A(_05956_),
    .B(_05955_),
    .Y(_05957_));
 sky130_fd_sc_hd__or2_1 _13934_ (.A(_05955_),
    .B(_05956_),
    .X(_05958_));
 sky130_fd_sc_hd__o311a_1 _13935_ (.A1(_00532_),
    .A2(net131),
    .A3(net130),
    .B1(_05957_),
    .C1(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__a2111oi_1 _13936_ (.A1(_05957_),
    .A2(_05958_),
    .B1(_00532_),
    .C1(net131),
    .D1(net130),
    .Y(_05961_));
 sky130_fd_sc_hd__nor2_2 _13937_ (.A(_05959_),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__xnor2_2 _13938_ (.A(_05946_),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a21oi_2 _13939_ (.A1(_05831_),
    .A2(_05827_),
    .B1(_05828_),
    .Y(_05964_));
 sky130_fd_sc_hd__xor2_4 _13940_ (.A(_05963_),
    .B(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__xnor2_1 _13941_ (.A(_05834_),
    .B(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__o21ba_1 _13942_ (.A1(_05877_),
    .A2(_05868_),
    .B1_N(_05886_),
    .X(_05967_));
 sky130_fd_sc_hd__a21oi_1 _13943_ (.A1(_05868_),
    .A2(_05877_),
    .B1(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__o32a_1 _13944_ (.A1(_01037_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_01188_),
    .B2(_02241_),
    .X(_05969_));
 sky130_fd_sc_hd__and4_1 _13945_ (.A(_02240_),
    .B(_02356_),
    .C(_01038_),
    .D(_01189_),
    .X(_05970_));
 sky130_fd_sc_hd__or4_1 _13946_ (.A(_01037_),
    .B(_01188_),
    .C(_02241_),
    .D(_02355_),
    .X(_05972_));
 sky130_fd_sc_hd__o32a_1 _13947_ (.A1(_00744_),
    .A2(_02628_),
    .A3(_02630_),
    .B1(_05969_),
    .B2(_05970_),
    .X(_05973_));
 sky130_fd_sc_hd__or4_1 _13948_ (.A(_00744_),
    .B(_02632_),
    .C(_05969_),
    .D(_05970_),
    .X(_05974_));
 sky130_fd_sc_hd__and2b_1 _13949_ (.A_N(_05973_),
    .B(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__a21oi_1 _13950_ (.A1(_00581_),
    .A2(_02858_),
    .B1(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__and3_1 _13951_ (.A(_05975_),
    .B(_02858_),
    .C(_00581_),
    .X(_05977_));
 sky130_fd_sc_hd__o21ai_1 _13952_ (.A1(_05976_),
    .A2(_05977_),
    .B1(_05881_),
    .Y(_05978_));
 sky130_fd_sc_hd__or3_1 _13953_ (.A(_05881_),
    .B(_05976_),
    .C(_05977_),
    .X(_05979_));
 sky130_fd_sc_hd__o21a_1 _13954_ (.A1(_05725_),
    .A2(_05882_),
    .B1(_05883_),
    .X(_05980_));
 sky130_fd_sc_hd__a21oi_1 _13955_ (.A1(_05978_),
    .A2(_05979_),
    .B1(_05980_),
    .Y(_05981_));
 sky130_fd_sc_hd__and3_1 _13956_ (.A(_05978_),
    .B(_05979_),
    .C(_05980_),
    .X(_05983_));
 sky130_fd_sc_hd__nor2_1 _13957_ (.A(_05981_),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__o21a_1 _13958_ (.A1(_05852_),
    .A2(_05860_),
    .B1(_05853_),
    .X(_05985_));
 sky130_fd_sc_hd__inv_2 _13959_ (.A(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__or3_1 _13960_ (.A(_01272_),
    .B(_02049_),
    .C(_02051_),
    .X(_05987_));
 sky130_fd_sc_hd__nand2_1 _13961_ (.A(_05841_),
    .B(_05848_),
    .Y(_05988_));
 sky130_fd_sc_hd__and3_1 _13962_ (.A(_05846_),
    .B(net137),
    .C(_01664_),
    .X(_05989_));
 sky130_fd_sc_hd__a31o_1 _13963_ (.A1(_01189_),
    .A2(_02054_),
    .A3(_05857_),
    .B1(_05855_),
    .X(_05990_));
 sky130_fd_sc_hd__o21a_1 _13964_ (.A1(_05845_),
    .A2(_05989_),
    .B1(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__a311oi_1 _13965_ (.A1(net137),
    .A2(_01664_),
    .A3(_05846_),
    .B1(_05990_),
    .C1(_05845_),
    .Y(_05992_));
 sky130_fd_sc_hd__or4_2 _13966_ (.A(net136),
    .B(_01589_),
    .C(_01662_),
    .D(_01882_),
    .X(_05994_));
 sky130_fd_sc_hd__o32a_1 _13967_ (.A1(_01589_),
    .A2(_01658_),
    .A3(_01660_),
    .B1(_01882_),
    .B2(net136),
    .X(_05995_));
 sky130_fd_sc_hd__a32o_1 _13968_ (.A1(net137),
    .A2(_01879_),
    .A3(net134),
    .B1(_01590_),
    .B2(_01664_),
    .X(_05996_));
 sky130_fd_sc_hd__a211o_1 _13969_ (.A1(_05994_),
    .A2(_05996_),
    .B1(_01542_),
    .C1(_01822_),
    .X(_05997_));
 sky130_fd_sc_hd__o211ai_1 _13970_ (.A1(_01542_),
    .A2(_01822_),
    .B1(_05994_),
    .C1(_05996_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand2_1 _13971_ (.A(_05997_),
    .B(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__or3_1 _13972_ (.A(_05991_),
    .B(_05992_),
    .C(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__a2bb2o_1 _13973_ (.A1_N(_05991_),
    .A2_N(_05992_),
    .B1(_05997_),
    .B2(_05998_),
    .X(_06001_));
 sky130_fd_sc_hd__nand2_1 _13974_ (.A(_06000_),
    .B(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__a21oi_1 _13975_ (.A1(_05842_),
    .A2(_05988_),
    .B1(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand3_1 _13976_ (.A(_05842_),
    .B(_05988_),
    .C(_06002_),
    .Y(_06005_));
 sky130_fd_sc_hd__and2b_1 _13977_ (.A_N(_06003_),
    .B(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__xnor2_1 _13978_ (.A(_05987_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__nor2_1 _13979_ (.A(_05986_),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_1 _13980_ (.A(_05986_),
    .B(_06007_),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2b_1 _13981_ (.A_N(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__o21ba_1 _13982_ (.A1(_05864_),
    .A2(_05867_),
    .B1_N(_05865_),
    .X(_06011_));
 sky130_fd_sc_hd__xnor2_2 _13983_ (.A(_06010_),
    .B(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__and3_1 _13984_ (.A(_02922_),
    .B(_02924_),
    .C(_00569_),
    .X(_06013_));
 sky130_fd_sc_hd__a31o_1 _13985_ (.A1(_00904_),
    .A2(_02693_),
    .A3(_02695_),
    .B1(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__o31ai_2 _13986_ (.A1(_00903_),
    .A2(_02925_),
    .A3(_05869_),
    .B1(_06014_),
    .Y(_06016_));
 sky130_fd_sc_hd__o31a_1 _13987_ (.A1(_01054_),
    .A2(_01056_),
    .A3(_02433_),
    .B1(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__or4_1 _13988_ (.A(_01054_),
    .B(_01056_),
    .C(_02433_),
    .D(_06016_),
    .X(_06018_));
 sky130_fd_sc_hd__nand2b_1 _13989_ (.A_N(_06017_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__a31o_1 _13990_ (.A1(_01222_),
    .A2(_02093_),
    .A3(_02095_),
    .B1(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__or4b_1 _13991_ (.A(_01221_),
    .B(net133),
    .C(_02094_),
    .D_N(_06019_),
    .X(_06021_));
 sky130_fd_sc_hd__nand2_1 _13992_ (.A(_06020_),
    .B(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__a41o_1 _13993_ (.A1(_00569_),
    .A2(_00904_),
    .A3(_02432_),
    .A4(_02697_),
    .B1(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__or4b_1 _13994_ (.A(_00903_),
    .B(_02433_),
    .C(_05869_),
    .D_N(_06022_),
    .X(_06024_));
 sky130_fd_sc_hd__a21boi_1 _13995_ (.A1(_05728_),
    .A2(_05874_),
    .B1_N(_05872_),
    .Y(_06025_));
 sky130_fd_sc_hd__a21oi_1 _13996_ (.A1(_06023_),
    .A2(_06024_),
    .B1(_06025_),
    .Y(_06027_));
 sky130_fd_sc_hd__and3_1 _13997_ (.A(_06023_),
    .B(_06024_),
    .C(_06025_),
    .X(_06028_));
 sky130_fd_sc_hd__nor2_1 _13998_ (.A(_06027_),
    .B(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__and3_1 _13999_ (.A(_05984_),
    .B(_06012_),
    .C(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__or2_1 _14000_ (.A(_06012_),
    .B(_06029_),
    .X(_06031_));
 sky130_fd_sc_hd__a2bb2o_1 _14001_ (.A1_N(_05981_),
    .A2_N(_05983_),
    .B1(_06012_),
    .B2(_06029_),
    .X(_06032_));
 sky130_fd_sc_hd__o21ai_2 _14002_ (.A1(_06012_),
    .A2(_06029_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__o22a_1 _14003_ (.A1(_05984_),
    .A2(_06031_),
    .B1(_06030_),
    .B2(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__nand2b_1 _14004_ (.A_N(_05968_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__nand2b_1 _14005_ (.A_N(_06034_),
    .B(_05968_),
    .Y(_06036_));
 sky130_fd_sc_hd__o21a_1 _14006_ (.A1(_05781_),
    .A2(_05888_),
    .B1(_05889_),
    .X(_06038_));
 sky130_fd_sc_hd__a21oi_1 _14007_ (.A1(_06035_),
    .A2(_06036_),
    .B1(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__and3_1 _14008_ (.A(_06035_),
    .B(_06036_),
    .C(_06038_),
    .X(_06040_));
 sky130_fd_sc_hd__nor2_1 _14009_ (.A(_06039_),
    .B(_06040_),
    .Y(_06041_));
 sky130_fd_sc_hd__nand2_1 _14010_ (.A(_05966_),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__inv_2 _14011_ (.A(_06042_),
    .Y(_06043_));
 sky130_fd_sc_hd__or2_1 _14012_ (.A(_05966_),
    .B(_06041_),
    .X(_06044_));
 sky130_fd_sc_hd__o21a_1 _14013_ (.A1(_05925_),
    .A2(_05683_),
    .B1(_05926_),
    .X(_06045_));
 sky130_fd_sc_hd__o21a_1 _14014_ (.A1(_05909_),
    .A2(_05911_),
    .B1(_05912_),
    .X(_06046_));
 sky130_fd_sc_hd__o32a_1 _14015_ (.A1(_00274_),
    .A2(_03444_),
    .A3(_03447_),
    .B1(net142),
    .B2(_03179_),
    .X(_06047_));
 sky130_fd_sc_hd__a32o_1 _14016_ (.A1(_00429_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_03450_),
    .B2(_00275_),
    .X(_06049_));
 sky130_fd_sc_hd__a31o_1 _14017_ (.A1(_00429_),
    .A2(_03450_),
    .A3(_05902_),
    .B1(_06047_),
    .X(_06050_));
 sky130_fd_sc_hd__xnor2_1 _14018_ (.A(_05898_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__a21boi_1 _14019_ (.A1(_05902_),
    .A2(_05905_),
    .B1_N(_05904_),
    .Y(_06052_));
 sky130_fd_sc_hd__o31a_1 _14020_ (.A1(net144),
    .A2(_03583_),
    .A3(_05601_),
    .B1(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__or4_1 _14021_ (.A(net144),
    .B(_03583_),
    .C(_05601_),
    .D(_06052_),
    .X(_06054_));
 sky130_fd_sc_hd__and2b_1 _14022_ (.A_N(_06053_),
    .B(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__and2b_1 _14023_ (.A_N(_06051_),
    .B(_06054_),
    .X(_06056_));
 sky130_fd_sc_hd__xor2_1 _14024_ (.A(_06051_),
    .B(_06055_),
    .X(_06057_));
 sky130_fd_sc_hd__or2_1 _14025_ (.A(_06046_),
    .B(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__nand2_1 _14026_ (.A(_06057_),
    .B(_06046_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _14027_ (.A(_06058_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__o31a_1 _14028_ (.A1(_00005_),
    .A2(_00007_),
    .A3(_03912_),
    .B1(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__o21a_1 _14029_ (.A1(_05916_),
    .A2(_05920_),
    .B1(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__o32ai_4 _14030_ (.A1(_05916_),
    .A2(_05920_),
    .A3(_06062_),
    .B1(_06063_),
    .B2(_06045_),
    .Y(_06064_));
 sky130_fd_sc_hd__o41a_1 _14031_ (.A1(_05916_),
    .A2(_05920_),
    .A3(_06062_),
    .A4(_06045_),
    .B1(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__a21o_1 _14032_ (.A1(_06045_),
    .A2(_06063_),
    .B1(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__a211o_1 _14033_ (.A1(_06045_),
    .A2(_06063_),
    .B1(_06065_),
    .C1(_05931_),
    .X(_06067_));
 sky130_fd_sc_hd__nand2_1 _14034_ (.A(_05931_),
    .B(_06066_),
    .Y(_06068_));
 sky130_fd_sc_hd__nand2_1 _14035_ (.A(_06067_),
    .B(_06068_),
    .Y(_06069_));
 sky130_fd_sc_hd__a21boi_1 _14036_ (.A1(_06042_),
    .A2(_06044_),
    .B1_N(_06069_),
    .Y(_06071_));
 sky130_fd_sc_hd__and3b_1 _14037_ (.A_N(_06069_),
    .B(_06044_),
    .C(_06042_),
    .X(_06072_));
 sky130_fd_sc_hd__nor2_1 _14038_ (.A(_06071_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__o21ai_1 _14039_ (.A1(_05894_),
    .A2(_05933_),
    .B1(_05893_),
    .Y(_06074_));
 sky130_fd_sc_hd__nor2_1 _14040_ (.A(_06073_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__inv_2 _14041_ (.A(_06075_),
    .Y(_06076_));
 sky130_fd_sc_hd__nand2_1 _14042_ (.A(_06073_),
    .B(_06074_),
    .Y(_06077_));
 sky130_fd_sc_hd__o2111ai_2 _14043_ (.A1(_05803_),
    .A2(_05934_),
    .B1(_05940_),
    .C1(_06076_),
    .D1(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__a22o_1 _14044_ (.A1(_05936_),
    .A2(_05940_),
    .B1(_06076_),
    .B2(_06077_),
    .X(_06079_));
 sky130_fd_sc_hd__and2_1 _14045_ (.A(_06078_),
    .B(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__o21ai_1 _14046_ (.A1(_00834_),
    .A2(_05944_),
    .B1(_06080_),
    .Y(_06082_));
 sky130_fd_sc_hd__a221o_1 _14047_ (.A1(_06078_),
    .A2(_06079_),
    .B1(_05800_),
    .B2(_05943_),
    .C1(_00834_),
    .X(_06083_));
 sky130_fd_sc_hd__and2_1 _14048_ (.A(_06082_),
    .B(_06083_),
    .X(net102));
 sky130_fd_sc_hd__o2111a_1 _14049_ (.A1(_05941_),
    .A2(_05942_),
    .B1(_06078_),
    .C1(_06079_),
    .D1(_05800_),
    .X(_06084_));
 sky130_fd_sc_hd__a31o_1 _14050_ (.A1(_06080_),
    .A2(_05943_),
    .A3(_05800_),
    .B1(_00834_),
    .X(_06085_));
 sky130_fd_sc_hd__o21ai_2 _14051_ (.A1(_06043_),
    .A2(_06069_),
    .B1(_06044_),
    .Y(_06086_));
 sky130_fd_sc_hd__a32o_1 _14052_ (.A1(_00367_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_00533_),
    .B2(_03320_),
    .X(_06087_));
 sky130_fd_sc_hd__or4_1 _14053_ (.A(_00366_),
    .B(_00532_),
    .C(_03319_),
    .D(_03652_),
    .X(_06088_));
 sky130_fd_sc_hd__o31a_1 _14054_ (.A1(_00532_),
    .A2(_03652_),
    .A3(_05819_),
    .B1(_06087_),
    .X(_06089_));
 sky130_fd_sc_hd__and3_1 _14055_ (.A(_03831_),
    .B(_00191_),
    .C(_00189_),
    .X(_06090_));
 sky130_fd_sc_hd__o21a_1 _14056_ (.A1(_06089_),
    .A2(_06090_),
    .B1(_05953_),
    .X(_06092_));
 sky130_fd_sc_hd__a311oi_4 _14057_ (.A1(_00189_),
    .A2(_03831_),
    .A3(_00191_),
    .B1(_06089_),
    .C1(_05953_),
    .Y(_06093_));
 sky130_fd_sc_hd__o21ai_1 _14058_ (.A1(_06092_),
    .A2(_06093_),
    .B1(_05948_),
    .Y(_06094_));
 sky130_fd_sc_hd__or3_1 _14059_ (.A(_05948_),
    .B(_06092_),
    .C(_06093_),
    .X(_06095_));
 sky130_fd_sc_hd__a2bb2o_1 _14060_ (.A1_N(_05955_),
    .A2_N(_05956_),
    .B1(_00533_),
    .B2(_03087_),
    .X(_06096_));
 sky130_fd_sc_hd__a22o_1 _14061_ (.A1(_06094_),
    .A2(_06095_),
    .B1(_06096_),
    .B2(_05957_),
    .X(_06097_));
 sky130_fd_sc_hd__and4_1 _14062_ (.A(_05957_),
    .B(_06094_),
    .C(_06095_),
    .D(_06096_),
    .X(_06098_));
 sky130_fd_sc_hd__nand4_1 _14063_ (.A(_05957_),
    .B(_06094_),
    .C(_06095_),
    .D(_06096_),
    .Y(_06099_));
 sky130_fd_sc_hd__and2_1 _14064_ (.A(_06097_),
    .B(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__a221o_1 _14065_ (.A1(_05946_),
    .A2(_05962_),
    .B1(_05831_),
    .B2(_05827_),
    .C1(_05828_),
    .X(_06101_));
 sky130_fd_sc_hd__o21ai_2 _14066_ (.A1(_05946_),
    .A2(_05962_),
    .B1(_06101_),
    .Y(_06103_));
 sky130_fd_sc_hd__xor2_2 _14067_ (.A(_06100_),
    .B(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__o21ba_1 _14068_ (.A1(_05834_),
    .A2(_05965_),
    .B1_N(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__nor3b_2 _14069_ (.A(_05834_),
    .B(_05965_),
    .C_N(_06104_),
    .Y(_06106_));
 sky130_fd_sc_hd__o31a_1 _14070_ (.A1(_01272_),
    .A2(_02053_),
    .A3(_06003_),
    .B1(_06005_),
    .X(_06107_));
 sky130_fd_sc_hd__and3_1 _14071_ (.A(_01544_),
    .B(_02050_),
    .C(_02052_),
    .X(_06108_));
 sky130_fd_sc_hd__o32a_1 _14072_ (.A1(_01658_),
    .A2(_01660_),
    .A3(_01822_),
    .B1(_01882_),
    .B2(_01589_),
    .X(_06109_));
 sky130_fd_sc_hd__and4_1 _14073_ (.A(_01590_),
    .B(_01664_),
    .C(_01823_),
    .D(_01883_),
    .X(_06110_));
 sky130_fd_sc_hd__nor2_1 _14074_ (.A(_06109_),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__xnor2_1 _14075_ (.A(_06108_),
    .B(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__o21bai_1 _14076_ (.A1(_05991_),
    .A2(_05999_),
    .B1_N(_05992_),
    .Y(_06114_));
 sky130_fd_sc_hd__and2_1 _14077_ (.A(_06114_),
    .B(_06112_),
    .X(_06115_));
 sky130_fd_sc_hd__nor2_1 _14078_ (.A(_06112_),
    .B(_06114_),
    .Y(_06116_));
 sky130_fd_sc_hd__or2_1 _14079_ (.A(_06115_),
    .B(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__o31a_1 _14080_ (.A1(_01542_),
    .A2(_01822_),
    .A3(_05995_),
    .B1(_05994_),
    .X(_06118_));
 sky130_fd_sc_hd__o311a_1 _14081_ (.A1(_01542_),
    .A2(_01822_),
    .A3(_05995_),
    .B1(_06117_),
    .C1(_05994_),
    .X(_06119_));
 sky130_fd_sc_hd__nor2_1 _14082_ (.A(_06117_),
    .B(_06118_),
    .Y(_06120_));
 sky130_fd_sc_hd__or3_1 _14083_ (.A(_06119_),
    .B(_06120_),
    .C(_06107_),
    .X(_06121_));
 sky130_fd_sc_hd__o221a_1 _14084_ (.A1(_06003_),
    .A2(_05987_),
    .B1(_06120_),
    .B2(_06119_),
    .C1(_06005_),
    .X(_06122_));
 sky130_fd_sc_hd__o21ai_1 _14085_ (.A1(_06119_),
    .A2(_06120_),
    .B1(_06107_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _14086_ (.A(_06121_),
    .B(_06123_),
    .Y(_06125_));
 sky130_fd_sc_hd__o21a_1 _14087_ (.A1(_06008_),
    .A2(_06011_),
    .B1(_06009_),
    .X(_06126_));
 sky130_fd_sc_hd__xnor2_2 _14088_ (.A(_06125_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__or4_1 _14089_ (.A(_01399_),
    .B(_01404_),
    .C(net133),
    .D(_02094_),
    .X(_06128_));
 sky130_fd_sc_hd__and3_1 _14090_ (.A(_01222_),
    .B(_02427_),
    .C(_02428_),
    .X(_06129_));
 sky130_fd_sc_hd__or4_1 _14091_ (.A(_00570_),
    .B(_00903_),
    .C(_02925_),
    .D(_03086_),
    .X(_06130_));
 sky130_fd_sc_hd__o32a_1 _14092_ (.A1(_00570_),
    .A2(net131),
    .A3(net130),
    .B1(_00903_),
    .B2(_02925_),
    .X(_06131_));
 sky130_fd_sc_hd__a31o_1 _14093_ (.A1(_00904_),
    .A2(_03087_),
    .A3(_06013_),
    .B1(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__o31a_1 _14094_ (.A1(_01058_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__o21ai_1 _14095_ (.A1(_01058_),
    .A2(_02696_),
    .B1(_06132_),
    .Y(_06134_));
 sky130_fd_sc_hd__and4b_1 _14096_ (.A_N(_06132_),
    .B(_02695_),
    .C(_02693_),
    .D(_01059_),
    .X(_06136_));
 sky130_fd_sc_hd__o21ai_1 _14097_ (.A1(_06133_),
    .A2(_06136_),
    .B1(_06129_),
    .Y(_06137_));
 sky130_fd_sc_hd__a311o_1 _14098_ (.A1(_01218_),
    .A2(_01220_),
    .A3(_02432_),
    .B1(_06133_),
    .C1(_06136_),
    .X(_06138_));
 sky130_fd_sc_hd__nand2_1 _14099_ (.A(_06137_),
    .B(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__a31oi_2 _14100_ (.A1(_00904_),
    .A2(_02697_),
    .A3(_06013_),
    .B1(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__or4b_1 _14101_ (.A(_00903_),
    .B(_02925_),
    .C(_05869_),
    .D_N(_06139_),
    .X(_06141_));
 sky130_fd_sc_hd__and2b_1 _14102_ (.A_N(_06140_),
    .B(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__xor2_1 _14103_ (.A(_06128_),
    .B(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__o32a_1 _14104_ (.A1(_01058_),
    .A2(_02433_),
    .A3(_06016_),
    .B1(_01221_),
    .B2(_02096_),
    .X(_06144_));
 sky130_fd_sc_hd__o21ai_1 _14105_ (.A1(_06017_),
    .A2(_06144_),
    .B1(_06143_),
    .Y(_06145_));
 sky130_fd_sc_hd__or3_1 _14106_ (.A(_06017_),
    .B(_06144_),
    .C(_06143_),
    .X(_06147_));
 sky130_fd_sc_hd__a21boi_1 _14107_ (.A1(_06024_),
    .A2(_06025_),
    .B1_N(_06023_),
    .Y(_06148_));
 sky130_fd_sc_hd__a21oi_1 _14108_ (.A1(_06145_),
    .A2(_06147_),
    .B1(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__and3_1 _14109_ (.A(_06145_),
    .B(_06147_),
    .C(_06148_),
    .X(_06150_));
 sky130_fd_sc_hd__or2_1 _14110_ (.A(_06149_),
    .B(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__nor2_1 _14111_ (.A(_06127_),
    .B(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2_1 _14112_ (.A(_06127_),
    .B(_06151_),
    .Y(_06153_));
 sky130_fd_sc_hd__nand2b_1 _14113_ (.A_N(_06152_),
    .B(_06153_),
    .Y(_06154_));
 sky130_fd_sc_hd__o31a_1 _14114_ (.A1(_00580_),
    .A2(_02857_),
    .A3(_05973_),
    .B1(_05974_),
    .X(_06155_));
 sky130_fd_sc_hd__a22o_1 _14115_ (.A1(_00741_),
    .A2(_00742_),
    .B1(_02852_),
    .B2(_02853_),
    .X(_06156_));
 sky130_fd_sc_hd__a32o_1 _14116_ (.A1(_01273_),
    .A2(_02236_),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_01189_),
    .X(_06158_));
 sky130_fd_sc_hd__or4_1 _14117_ (.A(_01188_),
    .B(_01272_),
    .C(_02241_),
    .D(_02355_),
    .X(_06159_));
 sky130_fd_sc_hd__nand2_1 _14118_ (.A(_06158_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__o31a_1 _14119_ (.A1(_01033_),
    .A2(_01035_),
    .A3(_02632_),
    .B1(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__or4_1 _14120_ (.A(_01033_),
    .B(_01035_),
    .C(_02632_),
    .D(_06160_),
    .X(_06162_));
 sky130_fd_sc_hd__and2b_1 _14121_ (.A_N(_06161_),
    .B(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__xor2_1 _14122_ (.A(_06156_),
    .B(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__o41a_1 _14123_ (.A1(_01037_),
    .A2(_01188_),
    .A3(_02241_),
    .A4(_02355_),
    .B1(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__or2_1 _14124_ (.A(_05972_),
    .B(_06164_),
    .X(_06166_));
 sky130_fd_sc_hd__nand2b_1 _14125_ (.A_N(_06165_),
    .B(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__o31a_1 _14126_ (.A1(_00580_),
    .A2(_03175_),
    .A3(_03177_),
    .B1(_06167_),
    .X(_06169_));
 sky130_fd_sc_hd__or4_1 _14127_ (.A(_00580_),
    .B(_03175_),
    .C(_03177_),
    .D(_06167_),
    .X(_06170_));
 sky130_fd_sc_hd__nand2b_1 _14128_ (.A_N(_06169_),
    .B(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__or2_1 _14129_ (.A(_06155_),
    .B(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__o311a_1 _14130_ (.A1(_00580_),
    .A2(_02857_),
    .A3(_05973_),
    .B1(_05974_),
    .C1(_06171_),
    .X(_06173_));
 sky130_fd_sc_hd__nand2_1 _14131_ (.A(_06155_),
    .B(_06171_),
    .Y(_06174_));
 sky130_fd_sc_hd__and2_1 _14132_ (.A(_06172_),
    .B(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__nand2_1 _14133_ (.A(_05979_),
    .B(_05980_),
    .Y(_06176_));
 sky130_fd_sc_hd__nand2_1 _14134_ (.A(_05978_),
    .B(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__xnor2_1 _14135_ (.A(_06175_),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__xnor2_1 _14136_ (.A(_06154_),
    .B(_06178_),
    .Y(_06180_));
 sky130_fd_sc_hd__and2_1 _14137_ (.A(_06033_),
    .B(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__nand2_1 _14138_ (.A(_06033_),
    .B(_06180_),
    .Y(_06182_));
 sky130_fd_sc_hd__or2_1 _14139_ (.A(_06033_),
    .B(_06180_),
    .X(_06183_));
 sky130_fd_sc_hd__a21boi_1 _14140_ (.A1(_06036_),
    .A2(_06038_),
    .B1_N(_06035_),
    .Y(_06184_));
 sky130_fd_sc_hd__or3b_1 _14141_ (.A(_06181_),
    .B(_06184_),
    .C_N(_06183_),
    .X(_06185_));
 sky130_fd_sc_hd__a21bo_1 _14142_ (.A1(_06182_),
    .A2(_06183_),
    .B1_N(_06184_),
    .X(_06186_));
 sky130_fd_sc_hd__a211oi_1 _14143_ (.A1(_06185_),
    .A2(_06186_),
    .B1(_06105_),
    .C1(_06106_),
    .Y(_06187_));
 sky130_fd_sc_hd__a211o_1 _14144_ (.A1(_06185_),
    .A2(_06186_),
    .B1(_06105_),
    .C1(_06106_),
    .X(_06188_));
 sky130_fd_sc_hd__o211a_1 _14145_ (.A1(_06105_),
    .A2(_06106_),
    .B1(_06185_),
    .C1(_06186_),
    .X(_06189_));
 sky130_fd_sc_hd__or2_1 _14146_ (.A(_06187_),
    .B(_06189_),
    .X(_06191_));
 sky130_fd_sc_hd__and4_1 _14147_ (.A(_00275_),
    .B(_00429_),
    .C(_03450_),
    .D(_03584_),
    .X(_06192_));
 sky130_fd_sc_hd__o32a_1 _14148_ (.A1(_00274_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(net142),
    .B2(_03449_),
    .X(_06193_));
 sky130_fd_sc_hd__o22a_1 _14149_ (.A1(_03912_),
    .A2(net144),
    .B1(_06193_),
    .B2(_06192_),
    .X(_06194_));
 sky130_fd_sc_hd__or3_1 _14150_ (.A(_06053_),
    .B(_06056_),
    .C(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__o21ai_1 _14151_ (.A1(_06053_),
    .A2(_06056_),
    .B1(_06194_),
    .Y(_06196_));
 sky130_fd_sc_hd__a32oi_4 _14152_ (.A1(_00429_),
    .A2(_03450_),
    .A3(_05902_),
    .B1(_05898_),
    .B2(_06049_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand3_1 _14153_ (.A(_06195_),
    .B(_06196_),
    .C(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__a21o_1 _14154_ (.A1(_06195_),
    .A2(_06196_),
    .B1(_06197_),
    .X(_06199_));
 sky130_fd_sc_hd__a21oi_1 _14155_ (.A1(_06198_),
    .A2(_06199_),
    .B1(_06060_),
    .Y(_06200_));
 sky130_fd_sc_hd__a21o_1 _14156_ (.A1(_06198_),
    .A2(_06199_),
    .B1(_06060_),
    .X(_06202_));
 sky130_fd_sc_hd__nand3_1 _14157_ (.A(_06060_),
    .B(_06198_),
    .C(_06199_),
    .Y(_06203_));
 sky130_fd_sc_hd__a21oi_1 _14158_ (.A1(_06202_),
    .A2(_06203_),
    .B1(_06064_),
    .Y(_06204_));
 sky130_fd_sc_hd__a21o_1 _14159_ (.A1(_06064_),
    .A2(_06203_),
    .B1(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__xnor2_1 _14160_ (.A(_06067_),
    .B(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__nor2_1 _14161_ (.A(_06191_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__and2_1 _14162_ (.A(_06191_),
    .B(_06206_),
    .X(_06208_));
 sky130_fd_sc_hd__nor2_1 _14163_ (.A(_06207_),
    .B(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__and2_1 _14164_ (.A(_06209_),
    .B(_06086_),
    .X(_06210_));
 sky130_fd_sc_hd__o221a_1 _14165_ (.A1(_06043_),
    .A2(_06069_),
    .B1(_06207_),
    .B2(_06208_),
    .C1(_06044_),
    .X(_06211_));
 sky130_fd_sc_hd__inv_2 _14166_ (.A(_06211_),
    .Y(_06213_));
 sky130_fd_sc_hd__o211ai_2 _14167_ (.A1(_05934_),
    .A2(_05803_),
    .B1(_06077_),
    .C1(_05940_),
    .Y(_06214_));
 sky130_fd_sc_hd__a31oi_1 _14168_ (.A1(_05936_),
    .A2(_05940_),
    .A3(_06077_),
    .B1(_06075_),
    .Y(_06215_));
 sky130_fd_sc_hd__o221a_1 _14169_ (.A1(_06073_),
    .A2(_06074_),
    .B1(_06210_),
    .B2(_06211_),
    .C1(_06214_),
    .X(_06216_));
 sky130_fd_sc_hd__a22oi_4 _14170_ (.A1(_06086_),
    .A2(_06209_),
    .B1(_06214_),
    .B2(_06076_),
    .Y(_06217_));
 sky130_fd_sc_hd__a21oi_2 _14171_ (.A1(_06217_),
    .A2(_06213_),
    .B1(_06216_),
    .Y(_06218_));
 sky130_fd_sc_hd__xor2_1 _14172_ (.A(_06085_),
    .B(_06218_),
    .X(net103));
 sky130_fd_sc_hd__and3_1 _14173_ (.A(_06218_),
    .B(_05944_),
    .C(_06080_),
    .X(_06219_));
 sky130_fd_sc_hd__inv_2 _14174_ (.A(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__a31o_1 _14175_ (.A1(_06218_),
    .A2(_05944_),
    .A3(_06080_),
    .B1(_00834_),
    .X(_06221_));
 sky130_fd_sc_hd__o21ai_2 _14176_ (.A1(_06189_),
    .A2(_06206_),
    .B1(_06188_),
    .Y(_06222_));
 sky130_fd_sc_hd__inv_2 _14177_ (.A(_06222_),
    .Y(_06223_));
 sky130_fd_sc_hd__and3_1 _14178_ (.A(_03831_),
    .B(_00364_),
    .C(_00362_),
    .X(_06224_));
 sky130_fd_sc_hd__a31o_1 _14179_ (.A1(_00533_),
    .A2(_03653_),
    .A3(_05819_),
    .B1(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__o21bai_2 _14180_ (.A1(_05948_),
    .A2(_06093_),
    .B1_N(_06092_),
    .Y(_06226_));
 sky130_fd_sc_hd__or2_1 _14181_ (.A(_06225_),
    .B(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__nand2_1 _14182_ (.A(_06226_),
    .B(_06225_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21o_1 _14183_ (.A1(_06103_),
    .A2(_06097_),
    .B1(_06098_),
    .X(_06229_));
 sky130_fd_sc_hd__a21oi_1 _14184_ (.A1(_06227_),
    .A2(_06228_),
    .B1(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__o21a_1 _14185_ (.A1(_06225_),
    .A2(_06226_),
    .B1(_06229_),
    .X(_06231_));
 sky130_fd_sc_hd__nor2_1 _14186_ (.A(_06230_),
    .B(_06231_),
    .Y(_06233_));
 sky130_fd_sc_hd__or2_1 _14187_ (.A(_06106_),
    .B(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__nand2_1 _14188_ (.A(_06106_),
    .B(_06233_),
    .Y(_06235_));
 sky130_fd_sc_hd__o21a_1 _14189_ (.A1(_06178_),
    .A2(_06152_),
    .B1(_06153_),
    .X(_06236_));
 sky130_fd_sc_hd__o32a_1 _14190_ (.A1(_01542_),
    .A2(_02053_),
    .A3(_06109_),
    .B1(_01589_),
    .B2(_01662_),
    .X(_06237_));
 sky130_fd_sc_hd__or3_1 _14191_ (.A(_01822_),
    .B(_01882_),
    .C(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__o32a_1 _14192_ (.A1(_01542_),
    .A2(_02053_),
    .A3(_06109_),
    .B1(_01822_),
    .B2(_01882_),
    .X(_06239_));
 sky130_fd_sc_hd__o31ai_2 _14193_ (.A1(_01662_),
    .A2(_02053_),
    .A3(_06239_),
    .B1(_06238_),
    .Y(_06240_));
 sky130_fd_sc_hd__o31a_1 _14194_ (.A1(_01658_),
    .A2(_01660_),
    .A3(_02053_),
    .B1(_06239_),
    .X(_06241_));
 sky130_fd_sc_hd__o32a_1 _14195_ (.A1(_01662_),
    .A2(_02053_),
    .A3(_06238_),
    .B1(_06241_),
    .B2(_06240_),
    .X(_06242_));
 sky130_fd_sc_hd__o21ba_1 _14196_ (.A1(_06118_),
    .A2(_06115_),
    .B1_N(_06116_),
    .X(_06244_));
 sky130_fd_sc_hd__and2_1 _14197_ (.A(_06242_),
    .B(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__nor2_1 _14198_ (.A(_06242_),
    .B(_06244_),
    .Y(_06246_));
 sky130_fd_sc_hd__o21a_1 _14199_ (.A1(_06122_),
    .A2(_06126_),
    .B1(_06121_),
    .X(_06247_));
 sky130_fd_sc_hd__o221a_1 _14200_ (.A1(_06245_),
    .A2(_06246_),
    .B1(_06122_),
    .B2(_06126_),
    .C1(_06121_),
    .X(_06248_));
 sky130_fd_sc_hd__nor3_2 _14201_ (.A(_06245_),
    .B(_06246_),
    .C(_06247_),
    .Y(_06249_));
 sky130_fd_sc_hd__o32a_1 _14202_ (.A1(_01221_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(net136),
    .B2(_02433_),
    .X(_06250_));
 sky130_fd_sc_hd__a31o_1 _14203_ (.A1(net137),
    .A2(_02697_),
    .A3(_06129_),
    .B1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__and4_1 _14204_ (.A(_00904_),
    .B(_03087_),
    .C(_03320_),
    .D(_00569_),
    .X(_06252_));
 sky130_fd_sc_hd__o32a_1 _14205_ (.A1(_00903_),
    .A2(net131),
    .A3(net130),
    .B1(_00570_),
    .B2(_03319_),
    .X(_06253_));
 sky130_fd_sc_hd__a32o_1 _14206_ (.A1(_00569_),
    .A2(_03316_),
    .A3(_03318_),
    .B1(_00904_),
    .B2(_03087_),
    .X(_06255_));
 sky130_fd_sc_hd__o32a_1 _14207_ (.A1(_01054_),
    .A2(_01056_),
    .A3(_02925_),
    .B1(_06252_),
    .B2(_06253_),
    .X(_06256_));
 sky130_fd_sc_hd__nor4_1 _14208_ (.A(_01058_),
    .B(_02925_),
    .C(_06252_),
    .D(_06253_),
    .Y(_06257_));
 sky130_fd_sc_hd__o21a_1 _14209_ (.A1(_06256_),
    .A2(_06257_),
    .B1(_06251_),
    .X(_06258_));
 sky130_fd_sc_hd__or3_1 _14210_ (.A(_06251_),
    .B(_06256_),
    .C(_06257_),
    .X(_06259_));
 sky130_fd_sc_hd__nand2b_1 _14211_ (.A_N(_06258_),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__xor2_1 _14212_ (.A(_06130_),
    .B(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__a31o_1 _14213_ (.A1(_01222_),
    .A2(_02432_),
    .A3(_06134_),
    .B1(_06136_),
    .X(_06262_));
 sky130_fd_sc_hd__a311o_1 _14214_ (.A1(_01222_),
    .A2(_02432_),
    .A3(_06134_),
    .B1(_06136_),
    .C1(_06261_),
    .X(_06263_));
 sky130_fd_sc_hd__nand2_1 _14215_ (.A(_06261_),
    .B(_06262_),
    .Y(_06264_));
 sky130_fd_sc_hd__a22oi_1 _14216_ (.A1(_01590_),
    .A2(_02097_),
    .B1(_06263_),
    .B2(_06264_),
    .Y(_06266_));
 sky130_fd_sc_hd__and4_1 _14217_ (.A(_01590_),
    .B(_02097_),
    .C(_06263_),
    .D(_06264_),
    .X(_06267_));
 sky130_fd_sc_hd__or2_1 _14218_ (.A(_06266_),
    .B(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__or4_1 _14219_ (.A(_01399_),
    .B(_01404_),
    .C(_02096_),
    .D(_06140_),
    .X(_06269_));
 sky130_fd_sc_hd__o311a_1 _14220_ (.A1(net136),
    .A2(_02096_),
    .A3(_06140_),
    .B1(_06141_),
    .C1(_06268_),
    .X(_06270_));
 sky130_fd_sc_hd__a21o_1 _14221_ (.A1(_06141_),
    .A2(_06269_),
    .B1(_06268_),
    .X(_06271_));
 sky130_fd_sc_hd__and2b_1 _14222_ (.A_N(_06270_),
    .B(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__a21boi_1 _14223_ (.A1(_06145_),
    .A2(_06148_),
    .B1_N(_06147_),
    .Y(_06273_));
 sky130_fd_sc_hd__xor2_1 _14224_ (.A(_06272_),
    .B(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__or3_1 _14225_ (.A(_06248_),
    .B(_06249_),
    .C(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__o21ai_1 _14226_ (.A1(_06248_),
    .A2(_06249_),
    .B1(_06274_),
    .Y(_06277_));
 sky130_fd_sc_hd__nand2_1 _14227_ (.A(_06275_),
    .B(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__a32o_1 _14228_ (.A1(_03176_),
    .A2(_03178_),
    .A3(_00743_),
    .B1(_01038_),
    .B2(_02858_),
    .X(_06279_));
 sky130_fd_sc_hd__o31a_1 _14229_ (.A1(_01037_),
    .A2(_03179_),
    .A3(_06156_),
    .B1(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__or4_1 _14230_ (.A(_01272_),
    .B(_01542_),
    .C(_02241_),
    .D(_02355_),
    .X(_06281_));
 sky130_fd_sc_hd__o32a_1 _14231_ (.A1(_01272_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_01542_),
    .B2(_02241_),
    .X(_06282_));
 sky130_fd_sc_hd__a32o_1 _14232_ (.A1(_01544_),
    .A2(_02236_),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_01273_),
    .X(_06283_));
 sky130_fd_sc_hd__a2111oi_1 _14233_ (.A1(_06281_),
    .A2(_06283_),
    .B1(_01184_),
    .C1(_01186_),
    .D1(_02632_),
    .Y(_06284_));
 sky130_fd_sc_hd__o311a_1 _14234_ (.A1(_01184_),
    .A2(_01186_),
    .A3(_02632_),
    .B1(_06281_),
    .C1(_06283_),
    .X(_06285_));
 sky130_fd_sc_hd__or3_2 _14235_ (.A(_06280_),
    .B(_06284_),
    .C(_06285_),
    .X(_06286_));
 sky130_fd_sc_hd__o21ai_1 _14236_ (.A1(_06284_),
    .A2(_06285_),
    .B1(_06280_),
    .Y(_06288_));
 sky130_fd_sc_hd__and3_1 _14237_ (.A(_06159_),
    .B(_06286_),
    .C(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__a21oi_1 _14238_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_06159_),
    .Y(_06290_));
 sky130_fd_sc_hd__nor2_1 _14239_ (.A(_06289_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__o31a_1 _14240_ (.A1(_00744_),
    .A2(_02857_),
    .A3(_06161_),
    .B1(_06162_),
    .X(_06292_));
 sky130_fd_sc_hd__nor2_1 _14241_ (.A(_06292_),
    .B(_06291_),
    .Y(_06293_));
 sky130_fd_sc_hd__o311a_1 _14242_ (.A1(_00744_),
    .A2(_02857_),
    .A3(_06161_),
    .B1(_06162_),
    .C1(_06291_),
    .X(_06294_));
 sky130_fd_sc_hd__or4_1 _14243_ (.A(_00580_),
    .B(_03449_),
    .C(_06293_),
    .D(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__o22ai_1 _14244_ (.A1(_00580_),
    .A2(_03449_),
    .B1(_06293_),
    .B2(_06294_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand2_1 _14245_ (.A(_06295_),
    .B(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__o31a_1 _14246_ (.A1(_00580_),
    .A2(_03179_),
    .A3(_06165_),
    .B1(_06166_),
    .X(_06299_));
 sky130_fd_sc_hd__xor2_1 _14247_ (.A(_06297_),
    .B(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__o21a_1 _14248_ (.A1(_06173_),
    .A2(_06177_),
    .B1(_06172_),
    .X(_06301_));
 sky130_fd_sc_hd__xor2_1 _14249_ (.A(_06300_),
    .B(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__xor2_1 _14250_ (.A(_06278_),
    .B(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__nor2_1 _14251_ (.A(_06236_),
    .B(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__nand2_1 _14252_ (.A(_06236_),
    .B(_06303_),
    .Y(_06305_));
 sky130_fd_sc_hd__nand2b_1 _14253_ (.A_N(_06304_),
    .B(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__o21ai_1 _14254_ (.A1(_06181_),
    .A2(_06184_),
    .B1(_06183_),
    .Y(_06307_));
 sky130_fd_sc_hd__or3b_1 _14255_ (.A(_06304_),
    .B(_06307_),
    .C_N(_06305_),
    .X(_06308_));
 sky130_fd_sc_hd__nand2_1 _14256_ (.A(_06306_),
    .B(_06307_),
    .Y(_06310_));
 sky130_fd_sc_hd__nand4_1 _14257_ (.A(_06234_),
    .B(_06235_),
    .C(_06308_),
    .D(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__a22oi_2 _14258_ (.A1(_06234_),
    .A2(_06235_),
    .B1(_06308_),
    .B2(_06310_),
    .Y(_06312_));
 sky130_fd_sc_hd__inv_2 _14259_ (.A(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__nand2_1 _14260_ (.A(_06311_),
    .B(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__o311a_1 _14261_ (.A1(_00274_),
    .A2(_03444_),
    .A3(_03447_),
    .B1(_03584_),
    .C1(_00429_),
    .X(_06315_));
 sky130_fd_sc_hd__a31o_1 _14262_ (.A1(_00271_),
    .A2(_00273_),
    .A3(_03911_),
    .B1(_06315_),
    .X(_06316_));
 sky130_fd_sc_hd__nand2_1 _14263_ (.A(_06195_),
    .B(_06197_),
    .Y(_06317_));
 sky130_fd_sc_hd__and3_1 _14264_ (.A(_06196_),
    .B(_06316_),
    .C(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__a21oi_1 _14265_ (.A1(_06196_),
    .A2(_06317_),
    .B1(_06316_),
    .Y(_06319_));
 sky130_fd_sc_hd__a21oi_1 _14266_ (.A1(_06064_),
    .A2(_06203_),
    .B1(_06200_),
    .Y(_06321_));
 sky130_fd_sc_hd__o21ai_1 _14267_ (.A1(_06318_),
    .A2(_06319_),
    .B1(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__o21ai_1 _14268_ (.A1(_06319_),
    .A2(_06321_),
    .B1(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__nor4_2 _14269_ (.A(_05931_),
    .B(_06066_),
    .C(_06205_),
    .D(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__o21ai_1 _14270_ (.A1(_06067_),
    .A2(_06205_),
    .B1(_06323_),
    .Y(_06325_));
 sky130_fd_sc_hd__nand2b_1 _14271_ (.A_N(_06324_),
    .B(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__xor2_2 _14272_ (.A(_06314_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__inv_2 _14273_ (.A(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__nand2_1 _14274_ (.A(_06327_),
    .B(_06222_),
    .Y(_06329_));
 sky130_fd_sc_hd__or2_1 _14275_ (.A(_06222_),
    .B(_06327_),
    .X(_06330_));
 sky130_fd_sc_hd__nand2_1 _14276_ (.A(_06329_),
    .B(_06330_),
    .Y(_06332_));
 sky130_fd_sc_hd__o21bai_1 _14277_ (.A1(_06211_),
    .A2(_06217_),
    .B1_N(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__o211ai_1 _14278_ (.A1(_06210_),
    .A2(_06215_),
    .B1(_06332_),
    .C1(_06213_),
    .Y(_06334_));
 sky130_fd_sc_hd__nand2_1 _14279_ (.A(_06333_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__xnor2_1 _14280_ (.A(_06221_),
    .B(_06335_),
    .Y(net104));
 sky130_fd_sc_hd__nand4_1 _14281_ (.A(_06084_),
    .B(_06218_),
    .C(_06333_),
    .D(_06334_),
    .Y(_06336_));
 sky130_fd_sc_hd__o21ai_2 _14282_ (.A1(_06312_),
    .A2(_06326_),
    .B1(_06311_),
    .Y(_06337_));
 sky130_fd_sc_hd__o21bai_1 _14283_ (.A1(_06319_),
    .A2(_06321_),
    .B1_N(_06318_),
    .Y(_06338_));
 sky130_fd_sc_hd__a2111oi_4 _14284_ (.A1(_00429_),
    .A2(net129),
    .B1(_06192_),
    .C1(_06324_),
    .D1(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__inv_2 _14285_ (.A(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__a21oi_1 _14286_ (.A1(_06225_),
    .A2(_06226_),
    .B1(_06231_),
    .Y(_06342_));
 sky130_fd_sc_hd__o2111a_1 _14287_ (.A1(_00532_),
    .A2(_03832_),
    .B1(_06088_),
    .C1(_06235_),
    .D1(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__a31o_2 _14288_ (.A1(_01879_),
    .A2(net134),
    .A3(_02054_),
    .B1(_06240_),
    .X(_06344_));
 sky130_fd_sc_hd__or4b_2 _14289_ (.A(_01882_),
    .B(_02049_),
    .C(_02051_),
    .D_N(_06240_),
    .X(_06345_));
 sky130_fd_sc_hd__o21ba_1 _14290_ (.A1(_06245_),
    .A2(_06247_),
    .B1_N(_06246_),
    .X(_06346_));
 sky130_fd_sc_hd__and3_1 _14291_ (.A(_06344_),
    .B(_06345_),
    .C(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__a21oi_1 _14292_ (.A1(_06344_),
    .A2(_06345_),
    .B1(_06346_),
    .Y(_06348_));
 sky130_fd_sc_hd__o21ai_1 _14293_ (.A1(_06130_),
    .A2(_06258_),
    .B1(_06259_),
    .Y(_06349_));
 sky130_fd_sc_hd__a31o_1 _14294_ (.A1(_01059_),
    .A2(_02926_),
    .A3(_06255_),
    .B1(_06252_),
    .X(_06350_));
 sky130_fd_sc_hd__a31oi_1 _14295_ (.A1(net137),
    .A2(_02697_),
    .A3(_06129_),
    .B1(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__nand4_1 _14296_ (.A(_02697_),
    .B(_06350_),
    .C(_06129_),
    .D(net137),
    .Y(_06353_));
 sky130_fd_sc_hd__and2b_1 _14297_ (.A_N(_06351_),
    .B(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__and3_1 _14298_ (.A(_01222_),
    .B(_02922_),
    .C(_02924_),
    .X(_06355_));
 sky130_fd_sc_hd__a32o_1 _14299_ (.A1(_00569_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_00904_),
    .B2(_03320_),
    .X(_06356_));
 sky130_fd_sc_hd__or3_1 _14300_ (.A(_00898_),
    .B(_00901_),
    .C(_03652_),
    .X(_06357_));
 sky130_fd_sc_hd__and4_1 _14301_ (.A(_00904_),
    .B(_03320_),
    .C(_03653_),
    .D(_00569_),
    .X(_06358_));
 sky130_fd_sc_hd__o31ai_1 _14302_ (.A1(_00570_),
    .A2(_03319_),
    .A3(_06357_),
    .B1(_06356_),
    .Y(_06359_));
 sky130_fd_sc_hd__and4b_1 _14303_ (.A_N(_06359_),
    .B(_03084_),
    .C(_03082_),
    .D(_01059_),
    .X(_06360_));
 sky130_fd_sc_hd__or4_1 _14304_ (.A(_01058_),
    .B(net131),
    .C(net130),
    .D(_06359_),
    .X(_06361_));
 sky130_fd_sc_hd__o21ai_1 _14305_ (.A1(_01058_),
    .A2(_03086_),
    .B1(_06359_),
    .Y(_06362_));
 sky130_fd_sc_hd__a32o_1 _14306_ (.A1(_01222_),
    .A2(_02922_),
    .A3(_02924_),
    .B1(_06361_),
    .B2(_06362_),
    .X(_06364_));
 sky130_fd_sc_hd__or4b_1 _14307_ (.A(_01221_),
    .B(_02925_),
    .C(_06360_),
    .D_N(_06362_),
    .X(_06365_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(_06364_),
    .B(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__xnor2_1 _14309_ (.A(_06354_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__or2_1 _14310_ (.A(_06349_),
    .B(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__nand2_1 _14311_ (.A(_06349_),
    .B(_06367_),
    .Y(_06369_));
 sky130_fd_sc_hd__or3_1 _14312_ (.A(_01822_),
    .B(net133),
    .C(_02094_),
    .X(_06370_));
 sky130_fd_sc_hd__o32a_1 _14313_ (.A1(net136),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_01589_),
    .B2(_02433_),
    .X(_06371_));
 sky130_fd_sc_hd__or4_1 _14314_ (.A(net136),
    .B(_01589_),
    .C(_02433_),
    .D(_02696_),
    .X(_06372_));
 sky130_fd_sc_hd__nand2b_1 _14315_ (.A_N(_06371_),
    .B(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__xnor2_1 _14316_ (.A(_06370_),
    .B(_06373_),
    .Y(_06375_));
 sky130_fd_sc_hd__a21o_1 _14317_ (.A1(_06368_),
    .A2(_06369_),
    .B1(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__nand3_1 _14318_ (.A(_06368_),
    .B(_06369_),
    .C(_06375_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand2_1 _14319_ (.A(_06376_),
    .B(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__or4b_1 _14320_ (.A(_01584_),
    .B(_01586_),
    .C(_02096_),
    .D_N(_06263_),
    .X(_06379_));
 sky130_fd_sc_hd__a21boi_1 _14321_ (.A1(_06264_),
    .A2(_06379_),
    .B1_N(_06378_),
    .Y(_06380_));
 sky130_fd_sc_hd__nand3b_1 _14322_ (.A_N(_06378_),
    .B(_06379_),
    .C(_06264_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2b_1 _14323_ (.A_N(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__o21ai_1 _14324_ (.A1(_06270_),
    .A2(_06273_),
    .B1(_06271_),
    .Y(_06383_));
 sky130_fd_sc_hd__and2_1 _14325_ (.A(_06383_),
    .B(_06382_),
    .X(_06384_));
 sky130_fd_sc_hd__nor2_1 _14326_ (.A(_06382_),
    .B(_06383_),
    .Y(_06386_));
 sky130_fd_sc_hd__o22a_1 _14327_ (.A1(_06347_),
    .A2(_06348_),
    .B1(_06384_),
    .B2(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__or4_2 _14328_ (.A(_06347_),
    .B(_06348_),
    .C(_06384_),
    .D(_06386_),
    .X(_06388_));
 sky130_fd_sc_hd__and2b_1 _14329_ (.A_N(_06387_),
    .B(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nand2_1 _14330_ (.A(_06159_),
    .B(_06288_),
    .Y(_06390_));
 sky130_fd_sc_hd__o31ai_1 _14331_ (.A1(_01188_),
    .A2(_02632_),
    .A3(_06282_),
    .B1(_06281_),
    .Y(_06391_));
 sky130_fd_sc_hd__or4b_1 _14332_ (.A(_01037_),
    .B(_03179_),
    .C(_06156_),
    .D_N(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__a41o_1 _14333_ (.A1(_00743_),
    .A2(_01038_),
    .A3(_02858_),
    .A4(_03180_),
    .B1(_06391_),
    .X(_06393_));
 sky130_fd_sc_hd__and3_1 _14334_ (.A(_01189_),
    .B(_02854_),
    .C(_02856_),
    .X(_06394_));
 sky130_fd_sc_hd__o32a_1 _14335_ (.A1(_01542_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_01662_),
    .B2(_02241_),
    .X(_06395_));
 sky130_fd_sc_hd__and4_2 _14336_ (.A(_02240_),
    .B(_02356_),
    .C(_01544_),
    .D(_01664_),
    .X(_06397_));
 sky130_fd_sc_hd__o22ai_2 _14337_ (.A1(_01272_),
    .A2(_02632_),
    .B1(_06395_),
    .B2(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__a2111oi_1 _14338_ (.A1(_01266_),
    .A2(_01267_),
    .B1(_02632_),
    .C1(_06395_),
    .D1(_06397_),
    .Y(_06399_));
 sky130_fd_sc_hd__or4_1 _14339_ (.A(_01272_),
    .B(_02632_),
    .C(_06395_),
    .D(_06397_),
    .X(_06400_));
 sky130_fd_sc_hd__o311a_1 _14340_ (.A1(_01184_),
    .A2(_01186_),
    .A3(_02857_),
    .B1(_06398_),
    .C1(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__a221oi_1 _14341_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_06398_),
    .B2(_06400_),
    .C1(_01188_),
    .Y(_06402_));
 sky130_fd_sc_hd__nor2_1 _14342_ (.A(_06401_),
    .B(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__inv_2 _14343_ (.A(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__a21oi_1 _14344_ (.A1(_06392_),
    .A2(_06393_),
    .B1(_06403_),
    .Y(_06405_));
 sky130_fd_sc_hd__and3_1 _14345_ (.A(_06392_),
    .B(_06393_),
    .C(_06403_),
    .X(_06406_));
 sky130_fd_sc_hd__o211ai_2 _14346_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06286_),
    .C1(_06390_),
    .Y(_06408_));
 sky130_fd_sc_hd__inv_2 _14347_ (.A(_06408_),
    .Y(_06409_));
 sky130_fd_sc_hd__a211o_1 _14348_ (.A1(_06286_),
    .A2(_06390_),
    .B1(_06405_),
    .C1(_06406_),
    .X(_06410_));
 sky130_fd_sc_hd__nand2_1 _14349_ (.A(_06408_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__and3_1 _14350_ (.A(_03448_),
    .B(_00743_),
    .C(_03445_),
    .X(_06412_));
 sky130_fd_sc_hd__and3_1 _14351_ (.A(_06412_),
    .B(_03180_),
    .C(_01038_),
    .X(_06413_));
 sky130_fd_sc_hd__o32a_1 _14352_ (.A1(_00744_),
    .A2(_03444_),
    .A3(_03447_),
    .B1(_01037_),
    .B2(_03179_),
    .X(_06414_));
 sky130_fd_sc_hd__a31o_1 _14353_ (.A1(_01038_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_06412_),
    .X(_06415_));
 sky130_fd_sc_hd__o211a_1 _14354_ (.A1(_06413_),
    .A2(_06414_),
    .B1(_00581_),
    .C1(_03584_),
    .X(_06416_));
 sky130_fd_sc_hd__a211o_1 _14355_ (.A1(_00581_),
    .A2(_03584_),
    .B1(_06413_),
    .C1(_06414_),
    .X(_06417_));
 sky130_fd_sc_hd__nand2b_1 _14356_ (.A_N(_06416_),
    .B(_06417_),
    .Y(_06419_));
 sky130_fd_sc_hd__xnor2_1 _14357_ (.A(_06411_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__a211oi_1 _14358_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_00580_),
    .C1(_03449_),
    .Y(_06421_));
 sky130_fd_sc_hd__o21a_1 _14359_ (.A1(_06293_),
    .A2(_06421_),
    .B1(_06420_),
    .X(_06422_));
 sky130_fd_sc_hd__nor3_1 _14360_ (.A(_06293_),
    .B(_06421_),
    .C(_06420_),
    .Y(_06423_));
 sky130_fd_sc_hd__o221a_1 _14361_ (.A1(_06297_),
    .A2(_06299_),
    .B1(_06177_),
    .B2(_06173_),
    .C1(_06172_),
    .X(_06424_));
 sky130_fd_sc_hd__a21o_1 _14362_ (.A1(_06297_),
    .A2(_06299_),
    .B1(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__o21ai_1 _14363_ (.A1(_06422_),
    .A2(_06423_),
    .B1(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__or3_1 _14364_ (.A(_06422_),
    .B(_06423_),
    .C(_06425_),
    .X(_06427_));
 sky130_fd_sc_hd__nand2_1 _14365_ (.A(_06426_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__inv_2 _14366_ (.A(_06428_),
    .Y(_06430_));
 sky130_fd_sc_hd__xnor2_1 _14367_ (.A(_06389_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__nand2b_1 _14368_ (.A_N(_06302_),
    .B(_06277_),
    .Y(_06432_));
 sky130_fd_sc_hd__o311a_1 _14369_ (.A1(_06248_),
    .A2(_06249_),
    .A3(_06274_),
    .B1(_06432_),
    .C1(_06431_),
    .X(_06433_));
 sky130_fd_sc_hd__a21oi_1 _14370_ (.A1(_06275_),
    .A2(_06432_),
    .B1(_06431_),
    .Y(_06434_));
 sky130_fd_sc_hd__o21a_1 _14371_ (.A1(_06304_),
    .A2(_06307_),
    .B1(_06305_),
    .X(_06435_));
 sky130_fd_sc_hd__o21ai_1 _14372_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__or3_1 _14373_ (.A(_06433_),
    .B(_06434_),
    .C(_06435_),
    .X(_06437_));
 sky130_fd_sc_hd__and3b_1 _14374_ (.A_N(_06343_),
    .B(_06436_),
    .C(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__a21bo_1 _14375_ (.A1(_06436_),
    .A2(_06437_),
    .B1_N(_06343_),
    .X(_06439_));
 sky130_fd_sc_hd__nand2b_1 _14376_ (.A_N(_06438_),
    .B(_06439_),
    .Y(_06441_));
 sky130_fd_sc_hd__xor2_2 _14377_ (.A(_06339_),
    .B(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__and2_1 _14378_ (.A(_06442_),
    .B(_06337_),
    .X(_06443_));
 sky130_fd_sc_hd__inv_2 _14379_ (.A(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__or2_2 _14380_ (.A(_06337_),
    .B(_06442_),
    .X(_06445_));
 sky130_fd_sc_hd__inv_2 _14381_ (.A(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__o21ai_2 _14382_ (.A1(_06222_),
    .A2(_06327_),
    .B1(_06213_),
    .Y(_06447_));
 sky130_fd_sc_hd__o21ai_1 _14383_ (.A1(_06447_),
    .A2(_06217_),
    .B1(_06329_),
    .Y(_06448_));
 sky130_fd_sc_hd__o221ai_2 _14384_ (.A1(_06447_),
    .A2(_06217_),
    .B1(_06443_),
    .B2(_06446_),
    .C1(_06329_),
    .Y(_06449_));
 sky130_fd_sc_hd__nand3_1 _14385_ (.A(_06448_),
    .B(_06445_),
    .C(_06444_),
    .Y(_06450_));
 sky130_fd_sc_hd__and2_1 _14386_ (.A(_06449_),
    .B(_06450_),
    .X(_06452_));
 sky130_fd_sc_hd__o221a_1 _14387_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_06335_),
    .B2(_06220_),
    .C1(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__a21oi_1 _14388_ (.A1(_00845_),
    .A2(_06336_),
    .B1(_06452_),
    .Y(_06454_));
 sky130_fd_sc_hd__nor2_1 _14389_ (.A(_06453_),
    .B(_06454_),
    .Y(net105));
 sky130_fd_sc_hd__a21oi_1 _14390_ (.A1(_06449_),
    .A2(_06450_),
    .B1(_06336_),
    .Y(_06455_));
 sky130_fd_sc_hd__o32a_1 _14391_ (.A1(_06335_),
    .A2(_06452_),
    .A3(_06220_),
    .B1(_00823_),
    .B2(_00812_),
    .X(_06456_));
 sky130_fd_sc_hd__a21oi_4 _14392_ (.A1(_06340_),
    .A2(_06439_),
    .B1(_06438_),
    .Y(_06457_));
 sky130_fd_sc_hd__a21oi_1 _14393_ (.A1(_06388_),
    .A2(_06430_),
    .B1(_06387_),
    .Y(_06458_));
 sky130_fd_sc_hd__a21boi_1 _14394_ (.A1(_06369_),
    .A2(_06375_),
    .B1_N(_06368_),
    .Y(_06459_));
 sky130_fd_sc_hd__a21o_1 _14395_ (.A1(_06353_),
    .A2(_06366_),
    .B1(_06351_),
    .X(_06460_));
 sky130_fd_sc_hd__a21oi_1 _14396_ (.A1(_06370_),
    .A2(_06372_),
    .B1(_06371_),
    .Y(_06462_));
 sky130_fd_sc_hd__a31o_1 _14397_ (.A1(_01222_),
    .A2(_02926_),
    .A3(_06362_),
    .B1(_06360_),
    .X(_06463_));
 sky130_fd_sc_hd__nand2_1 _14398_ (.A(_06463_),
    .B(_06462_),
    .Y(_06464_));
 sky130_fd_sc_hd__a311o_1 _14399_ (.A1(_01222_),
    .A2(_02926_),
    .A3(_06362_),
    .B1(_06462_),
    .C1(_06360_),
    .X(_06465_));
 sky130_fd_sc_hd__and3_1 _14400_ (.A(net137),
    .B(_06355_),
    .C(_03087_),
    .X(_06466_));
 sky130_fd_sc_hd__o32a_1 _14401_ (.A1(_01221_),
    .A2(net131),
    .A3(net130),
    .B1(net136),
    .B2(_02925_),
    .X(_06467_));
 sky130_fd_sc_hd__a32o_1 _14402_ (.A1(_00904_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_01059_),
    .B2(_03320_),
    .X(_06468_));
 sky130_fd_sc_hd__or4_1 _14403_ (.A(_00903_),
    .B(_01058_),
    .C(_03319_),
    .D(_03652_),
    .X(_06469_));
 sky130_fd_sc_hd__o2bb2a_1 _14404_ (.A1_N(_06468_),
    .A2_N(_06469_),
    .B1(_00570_),
    .B2(_03832_),
    .X(_06470_));
 sky130_fd_sc_hd__o21ai_1 _14405_ (.A1(_06466_),
    .A2(_06467_),
    .B1(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__a311o_1 _14406_ (.A1(net137),
    .A2(_03087_),
    .A3(_06355_),
    .B1(_06467_),
    .C1(_06470_),
    .X(_06473_));
 sky130_fd_sc_hd__a21oi_1 _14407_ (.A1(_06471_),
    .A2(_06473_),
    .B1(_06358_),
    .Y(_06474_));
 sky130_fd_sc_hd__and3_1 _14408_ (.A(_06473_),
    .B(_06358_),
    .C(_06471_),
    .X(_06475_));
 sky130_fd_sc_hd__or2_1 _14409_ (.A(_06474_),
    .B(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__and3_1 _14410_ (.A(_06464_),
    .B(_06465_),
    .C(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__a21oi_1 _14411_ (.A1(_06464_),
    .A2(_06465_),
    .B1(_06476_),
    .Y(_06478_));
 sky130_fd_sc_hd__nor2_1 _14412_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__xnor2_1 _14413_ (.A(_06460_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__or4_1 _14414_ (.A(_02049_),
    .B(_02051_),
    .C(net133),
    .D(_02094_),
    .X(_06481_));
 sky130_fd_sc_hd__o32a_1 _14415_ (.A1(_01589_),
    .A2(_02692_),
    .A3(_02694_),
    .B1(_01822_),
    .B2(_02433_),
    .X(_06482_));
 sky130_fd_sc_hd__or4_1 _14416_ (.A(_01589_),
    .B(_01822_),
    .C(_02433_),
    .D(_02696_),
    .X(_06484_));
 sky130_fd_sc_hd__nand2b_1 _14417_ (.A_N(_06482_),
    .B(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__xor2_1 _14418_ (.A(_06481_),
    .B(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__xnor2_1 _14419_ (.A(_06480_),
    .B(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nor2_1 _14420_ (.A(_06459_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand2_1 _14421_ (.A(_06487_),
    .B(_06459_),
    .Y(_06489_));
 sky130_fd_sc_hd__and2b_1 _14422_ (.A_N(_06488_),
    .B(_06489_),
    .X(_06490_));
 sky130_fd_sc_hd__a21oi_1 _14423_ (.A1(_06383_),
    .A2(_06381_),
    .B1(_06380_),
    .Y(_06491_));
 sky130_fd_sc_hd__xor2_1 _14424_ (.A(_06490_),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__nand2_1 _14425_ (.A(_06345_),
    .B(_06346_),
    .Y(_06493_));
 sky130_fd_sc_hd__a21boi_1 _14426_ (.A1(_06344_),
    .A2(_06493_),
    .B1_N(_06492_),
    .Y(_06495_));
 sky130_fd_sc_hd__and3b_1 _14427_ (.A_N(_06492_),
    .B(_06493_),
    .C(_06344_),
    .X(_06496_));
 sky130_fd_sc_hd__nor2_1 _14428_ (.A(_06495_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__or3_1 _14429_ (.A(_03582_),
    .B(_00744_),
    .C(_03581_),
    .X(_06498_));
 sky130_fd_sc_hd__o32a_1 _14430_ (.A1(_03582_),
    .A2(_00744_),
    .A3(_03581_),
    .B1(_01037_),
    .B2(_03449_),
    .X(_06499_));
 sky130_fd_sc_hd__a31o_1 _14431_ (.A1(_01038_),
    .A2(_03584_),
    .A3(_06412_),
    .B1(_06499_),
    .X(_06500_));
 sky130_fd_sc_hd__o21ai_2 _14432_ (.A1(_00580_),
    .A2(_03912_),
    .B1(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__a31o_1 _14433_ (.A1(_00581_),
    .A2(_03584_),
    .A3(_06415_),
    .B1(_06413_),
    .X(_06502_));
 sky130_fd_sc_hd__a31o_1 _14434_ (.A1(_01189_),
    .A2(_02858_),
    .A3(_06398_),
    .B1(_06399_),
    .X(_06503_));
 sky130_fd_sc_hd__nor2_1 _14435_ (.A(_06502_),
    .B(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__nand2_1 _14436_ (.A(_06503_),
    .B(_06502_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand2b_2 _14437_ (.A_N(_06504_),
    .B(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__o32a_1 _14438_ (.A1(_01188_),
    .A2(_03175_),
    .A3(_03177_),
    .B1(_01272_),
    .B2(_02857_),
    .X(_06508_));
 sky130_fd_sc_hd__and3_1 _14439_ (.A(_06394_),
    .B(_03180_),
    .C(_01273_),
    .X(_06509_));
 sky130_fd_sc_hd__or4_1 _14440_ (.A(_01188_),
    .B(_01272_),
    .C(_02857_),
    .D(_03179_),
    .X(_06510_));
 sky130_fd_sc_hd__nor2_1 _14441_ (.A(_06508_),
    .B(_06509_),
    .Y(_06511_));
 sky130_fd_sc_hd__and3_1 _14442_ (.A(_01879_),
    .B(net134),
    .C(_02356_),
    .X(_06512_));
 sky130_fd_sc_hd__or4_1 _14443_ (.A(_01662_),
    .B(_01882_),
    .C(_02241_),
    .D(_02355_),
    .X(_06513_));
 sky130_fd_sc_hd__o32a_1 _14444_ (.A1(_01662_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_01882_),
    .B2(_02241_),
    .X(_06514_));
 sky130_fd_sc_hd__a32o_1 _14445_ (.A1(_01883_),
    .A2(_02236_),
    .A3(_02237_),
    .B1(_02356_),
    .B2(_01664_),
    .X(_06515_));
 sky130_fd_sc_hd__a22oi_1 _14446_ (.A1(_01544_),
    .A2(_02633_),
    .B1(_06513_),
    .B2(_06515_),
    .Y(_06517_));
 sky130_fd_sc_hd__and4_1 _14447_ (.A(_01544_),
    .B(_02633_),
    .C(_06513_),
    .D(_06515_),
    .X(_06518_));
 sky130_fd_sc_hd__nor2_1 _14448_ (.A(_06517_),
    .B(_06518_),
    .Y(_06519_));
 sky130_fd_sc_hd__xor2_2 _14449_ (.A(_06511_),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__xnor2_4 _14450_ (.A(_06397_),
    .B(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__xor2_4 _14451_ (.A(_06507_),
    .B(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__a21bo_2 _14452_ (.A1(_06404_),
    .A2(_06393_),
    .B1_N(_06392_),
    .X(_06523_));
 sky130_fd_sc_hd__a21o_1 _14453_ (.A1(_06522_),
    .A2(_06523_),
    .B1(_06501_),
    .X(_06524_));
 sky130_fd_sc_hd__o21a_1 _14454_ (.A1(_06522_),
    .A2(_06523_),
    .B1(_06501_),
    .X(_06525_));
 sky130_fd_sc_hd__o21ai_1 _14455_ (.A1(_06522_),
    .A2(_06523_),
    .B1(_06524_),
    .Y(_06526_));
 sky130_fd_sc_hd__o31a_1 _14456_ (.A1(_06501_),
    .A2(_06522_),
    .A3(_06523_),
    .B1(_06526_),
    .X(_06528_));
 sky130_fd_sc_hd__a31oi_2 _14457_ (.A1(_06501_),
    .A2(_06522_),
    .A3(_06523_),
    .B1(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__o21ai_2 _14458_ (.A1(_06409_),
    .A2(_06419_),
    .B1(_06410_),
    .Y(_06530_));
 sky130_fd_sc_hd__xor2_1 _14459_ (.A(_06529_),
    .B(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__o21ba_1 _14460_ (.A1(_06423_),
    .A2(_06425_),
    .B1_N(_06422_),
    .X(_06532_));
 sky130_fd_sc_hd__xor2_2 _14461_ (.A(_06531_),
    .B(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__and2_1 _14462_ (.A(_06497_),
    .B(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__nor2_1 _14463_ (.A(_06533_),
    .B(_06497_),
    .Y(_06535_));
 sky130_fd_sc_hd__a2111oi_4 _14464_ (.A1(_06388_),
    .A2(_06430_),
    .B1(_06534_),
    .C1(_06535_),
    .D1(_06387_),
    .Y(_06536_));
 sky130_fd_sc_hd__o21ba_1 _14465_ (.A1(_06534_),
    .A2(_06535_),
    .B1_N(_06458_),
    .X(_06537_));
 sky130_fd_sc_hd__inv_2 _14466_ (.A(_06537_),
    .Y(_06539_));
 sky130_fd_sc_hd__nor2_2 _14467_ (.A(_06536_),
    .B(_06537_),
    .Y(_06540_));
 sky130_fd_sc_hd__o21ba_4 _14468_ (.A1(_06433_),
    .A2(_06435_),
    .B1_N(_06434_),
    .X(_06541_));
 sky130_fd_sc_hd__xor2_4 _14469_ (.A(_06540_),
    .B(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__nand2_4 _14470_ (.A(_06457_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__or2_2 _14471_ (.A(_06457_),
    .B(_06542_),
    .X(_06544_));
 sky130_fd_sc_hd__inv_2 _14472_ (.A(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__o221ai_4 _14473_ (.A1(_06223_),
    .A2(_06328_),
    .B1(_06447_),
    .B2(_06217_),
    .C1(_06444_),
    .Y(_06546_));
 sky130_fd_sc_hd__a22o_1 _14474_ (.A1(_06543_),
    .A2(_06544_),
    .B1(_06546_),
    .B2(_06445_),
    .X(_06547_));
 sky130_fd_sc_hd__o2111ai_2 _14475_ (.A1(_06337_),
    .A2(_06442_),
    .B1(_06543_),
    .C1(_06544_),
    .D1(_06546_),
    .Y(_06548_));
 sky130_fd_sc_hd__nand2_1 _14476_ (.A(_06547_),
    .B(_06548_),
    .Y(_06550_));
 sky130_fd_sc_hd__xnor2_1 _14477_ (.A(_06456_),
    .B(_06550_),
    .Y(net106));
 sky130_fd_sc_hd__a2111oi_1 _14478_ (.A1(_06547_),
    .A2(_06548_),
    .B1(_06335_),
    .C1(_06452_),
    .D1(_06220_),
    .Y(_06551_));
 sky130_fd_sc_hd__a2bb2o_1 _14479_ (.A1_N(_00812_),
    .A2_N(_00823_),
    .B1(_06455_),
    .B2(_06550_),
    .X(_06552_));
 sky130_fd_sc_hd__a21oi_2 _14480_ (.A1(_06539_),
    .A2(_06541_),
    .B1(_06536_),
    .Y(_06553_));
 sky130_fd_sc_hd__o21a_1 _14481_ (.A1(_06511_),
    .A2(_06519_),
    .B1(_06397_),
    .X(_06554_));
 sky130_fd_sc_hd__a21oi_1 _14482_ (.A1(_06511_),
    .A2(_06519_),
    .B1(_06554_),
    .Y(_06555_));
 sky130_fd_sc_hd__nor2_1 _14483_ (.A(_06498_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__or4_1 _14484_ (.A(_01037_),
    .B(_03449_),
    .C(_06498_),
    .D(_06555_),
    .X(_06557_));
 sky130_fd_sc_hd__o31a_1 _14485_ (.A1(_01037_),
    .A2(_03449_),
    .A3(_06498_),
    .B1(_06555_),
    .X(_06558_));
 sky130_fd_sc_hd__a31o_1 _14486_ (.A1(_06556_),
    .A2(_03450_),
    .A3(_01038_),
    .B1(_06558_),
    .X(_06560_));
 sky130_fd_sc_hd__a32o_1 _14487_ (.A1(_01273_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_03450_),
    .B2(_01189_),
    .X(_06561_));
 sky130_fd_sc_hd__or4_1 _14488_ (.A(_01188_),
    .B(_01272_),
    .C(_03179_),
    .D(_03449_),
    .X(_06562_));
 sky130_fd_sc_hd__nand2_1 _14489_ (.A(_06561_),
    .B(_06562_),
    .Y(_06563_));
 sky130_fd_sc_hd__and3_1 _14490_ (.A(_06512_),
    .B(_02633_),
    .C(_01664_),
    .X(_06564_));
 sky130_fd_sc_hd__o32a_1 _14491_ (.A1(_01662_),
    .A2(_02628_),
    .A3(_02630_),
    .B1(_01882_),
    .B2(_02355_),
    .X(_06565_));
 sky130_fd_sc_hd__a31o_1 _14492_ (.A1(_01659_),
    .A2(net140),
    .A3(_02633_),
    .B1(_06512_),
    .X(_06566_));
 sky130_fd_sc_hd__o32a_1 _14493_ (.A1(_01538_),
    .A2(_01540_),
    .A3(_02857_),
    .B1(_06564_),
    .B2(_06565_),
    .X(_06567_));
 sky130_fd_sc_hd__nor4_1 _14494_ (.A(_01542_),
    .B(_02857_),
    .C(_06564_),
    .D(_06565_),
    .Y(_06568_));
 sky130_fd_sc_hd__o21ai_1 _14495_ (.A1(_06567_),
    .A2(_06568_),
    .B1(_06563_),
    .Y(_06569_));
 sky130_fd_sc_hd__or3_1 _14496_ (.A(_06563_),
    .B(_06567_),
    .C(_06568_),
    .X(_06571_));
 sky130_fd_sc_hd__o31ai_2 _14497_ (.A1(_01542_),
    .A2(_02632_),
    .A3(_06514_),
    .B1(_06513_),
    .Y(_06572_));
 sky130_fd_sc_hd__a21oi_1 _14498_ (.A1(_06569_),
    .A2(_06571_),
    .B1(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__and3_1 _14499_ (.A(_06569_),
    .B(_06571_),
    .C(_06572_),
    .X(_06574_));
 sky130_fd_sc_hd__or2_1 _14500_ (.A(_06573_),
    .B(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__and2_1 _14501_ (.A(_06560_),
    .B(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__nor2_1 _14502_ (.A(_06560_),
    .B(_06575_),
    .Y(_06577_));
 sky130_fd_sc_hd__or2_1 _14503_ (.A(_06504_),
    .B(_06521_),
    .X(_06578_));
 sky130_fd_sc_hd__a211oi_1 _14504_ (.A1(_06506_),
    .A2(_06578_),
    .B1(_06577_),
    .C1(_06576_),
    .Y(_06579_));
 sky130_fd_sc_hd__a211o_1 _14505_ (.A1(_06506_),
    .A2(_06578_),
    .B1(_06577_),
    .C1(_06576_),
    .X(_06580_));
 sky130_fd_sc_hd__o221a_1 _14506_ (.A1(_06504_),
    .A2(_06521_),
    .B1(_06576_),
    .B2(_06577_),
    .C1(_06506_),
    .X(_06582_));
 sky130_fd_sc_hd__or4_2 _14507_ (.A(_01037_),
    .B(_03581_),
    .C(_03582_),
    .D(_06510_),
    .X(_06583_));
 sky130_fd_sc_hd__a31o_1 _14508_ (.A1(_01034_),
    .A2(_01036_),
    .A3(_03584_),
    .B1(_06509_),
    .X(_06584_));
 sky130_fd_sc_hd__o2bb2a_1 _14509_ (.A1_N(_06583_),
    .A2_N(_06584_),
    .B1(_00744_),
    .B2(_03912_),
    .X(_06585_));
 sky130_fd_sc_hd__a221o_1 _14510_ (.A1(_00743_),
    .A2(net129),
    .B1(_06583_),
    .B2(_06584_),
    .C1(_06579_),
    .X(_06586_));
 sky130_fd_sc_hd__o21bai_1 _14511_ (.A1(_06579_),
    .A2(_06582_),
    .B1_N(_06585_),
    .Y(_06587_));
 sky130_fd_sc_hd__o21ai_1 _14512_ (.A1(_06582_),
    .A2(_06586_),
    .B1(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__a211o_1 _14513_ (.A1(_06522_),
    .A2(_06523_),
    .B1(_06525_),
    .C1(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__o211a_1 _14514_ (.A1(_06522_),
    .A2(_06523_),
    .B1(_06524_),
    .C1(_06588_),
    .X(_06590_));
 sky130_fd_sc_hd__o211ai_1 _14515_ (.A1(_06522_),
    .A2(_06523_),
    .B1(_06524_),
    .C1(_06588_),
    .Y(_06591_));
 sky130_fd_sc_hd__nand2_1 _14516_ (.A(_06589_),
    .B(_06591_),
    .Y(_06593_));
 sky130_fd_sc_hd__a21o_1 _14517_ (.A1(_06529_),
    .A2(_06530_),
    .B1(_06532_),
    .X(_06594_));
 sky130_fd_sc_hd__o21ai_2 _14518_ (.A1(_06529_),
    .A2(_06530_),
    .B1(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__xor2_2 _14519_ (.A(_06593_),
    .B(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__a21bo_1 _14520_ (.A1(_06479_),
    .A2(_06460_),
    .B1_N(_06486_),
    .X(_06597_));
 sky130_fd_sc_hd__o21a_1 _14521_ (.A1(_06460_),
    .A2(_06479_),
    .B1(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__a21boi_1 _14522_ (.A1(_06358_),
    .A2(_06471_),
    .B1_N(_06473_),
    .Y(_06599_));
 sky130_fd_sc_hd__o311a_1 _14523_ (.A1(_02053_),
    .A2(_02096_),
    .A3(_06482_),
    .B1(_06484_),
    .C1(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__a211oi_1 _14524_ (.A1(_06481_),
    .A2(_06484_),
    .B1(_06482_),
    .C1(_06599_),
    .Y(_06601_));
 sky130_fd_sc_hd__and3_1 _14525_ (.A(_01590_),
    .B(_02922_),
    .C(_02924_),
    .X(_06602_));
 sky130_fd_sc_hd__and3_1 _14526_ (.A(net137),
    .B(_06602_),
    .C(_03087_),
    .X(_06604_));
 sky130_fd_sc_hd__o32a_1 _14527_ (.A1(net136),
    .A2(net131),
    .A3(net130),
    .B1(_01589_),
    .B2(_02925_),
    .X(_06605_));
 sky130_fd_sc_hd__and3_1 _14528_ (.A(_01222_),
    .B(_03316_),
    .C(_03318_),
    .X(_06606_));
 sky130_fd_sc_hd__a31o_1 _14529_ (.A1(_01059_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__or3_1 _14530_ (.A(_01217_),
    .B(_01219_),
    .C(_03652_),
    .X(_06608_));
 sky130_fd_sc_hd__or4_1 _14531_ (.A(_01058_),
    .B(_01221_),
    .C(_03319_),
    .D(_03652_),
    .X(_06609_));
 sky130_fd_sc_hd__nand2_1 _14532_ (.A(_06607_),
    .B(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__o31a_1 _14533_ (.A1(_00898_),
    .A2(_00901_),
    .A3(_03832_),
    .B1(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__or3_1 _14534_ (.A(_06604_),
    .B(_06605_),
    .C(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__o221a_1 _14535_ (.A1(_00903_),
    .A2(_03834_),
    .B1(_06604_),
    .B2(_06605_),
    .C1(_06610_),
    .X(_06613_));
 sky130_fd_sc_hd__o21ai_1 _14536_ (.A1(_06604_),
    .A2(_06605_),
    .B1(_06611_),
    .Y(_06615_));
 sky130_fd_sc_hd__a21bo_1 _14537_ (.A1(_06612_),
    .A2(_06615_),
    .B1_N(_06469_),
    .X(_06616_));
 sky130_fd_sc_hd__or3b_1 _14538_ (.A(_06613_),
    .B(_06469_),
    .C_N(_06612_),
    .X(_06617_));
 sky130_fd_sc_hd__nand2_1 _14539_ (.A(_06616_),
    .B(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__o21bai_1 _14540_ (.A1(_06600_),
    .A2(_06601_),
    .B1_N(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__or3b_1 _14541_ (.A(_06600_),
    .B(_06601_),
    .C_N(_06618_),
    .X(_06620_));
 sky130_fd_sc_hd__nand2_1 _14542_ (.A(_06619_),
    .B(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__nand2_1 _14543_ (.A(_06464_),
    .B(_06476_),
    .Y(_06622_));
 sky130_fd_sc_hd__and3_1 _14544_ (.A(_06465_),
    .B(_06621_),
    .C(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__a21o_1 _14545_ (.A1(_06465_),
    .A2(_06622_),
    .B1(_06621_),
    .X(_06624_));
 sky130_fd_sc_hd__and2b_1 _14546_ (.A_N(_06623_),
    .B(_06624_),
    .X(_06626_));
 sky130_fd_sc_hd__or3_1 _14547_ (.A(_02049_),
    .B(_02051_),
    .C(_02433_),
    .X(_06627_));
 sky130_fd_sc_hd__and3_1 _14548_ (.A(_06466_),
    .B(_02697_),
    .C(_01823_),
    .X(_06628_));
 sky130_fd_sc_hd__a21oi_1 _14549_ (.A1(_01823_),
    .A2(_02697_),
    .B1(_06466_),
    .Y(_06629_));
 sky130_fd_sc_hd__a311o_1 _14550_ (.A1(_02050_),
    .A2(_02432_),
    .A3(_02052_),
    .B1(_06629_),
    .C1(_06628_),
    .X(_06630_));
 sky130_fd_sc_hd__o2111ai_1 _14551_ (.A1(_06628_),
    .A2(_06629_),
    .B1(_02050_),
    .C1(_02052_),
    .D1(_02432_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_1 _14552_ (.A(_06630_),
    .B(_06631_),
    .Y(_06632_));
 sky130_fd_sc_hd__xnor2_1 _14553_ (.A(_06626_),
    .B(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__xor2_1 _14554_ (.A(_06598_),
    .B(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__o21ai_1 _14555_ (.A1(_06488_),
    .A2(_06491_),
    .B1(_06489_),
    .Y(_06635_));
 sky130_fd_sc_hd__xnor2_1 _14556_ (.A(_06634_),
    .B(_06635_),
    .Y(_06637_));
 sky130_fd_sc_hd__or4_1 _14557_ (.A(net133),
    .B(_02094_),
    .C(_02241_),
    .D(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__o31a_1 _14558_ (.A1(net133),
    .A2(_02094_),
    .A3(_02241_),
    .B1(_06637_),
    .X(_06639_));
 sky130_fd_sc_hd__nand2_1 _14559_ (.A(_06596_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__o21a_1 _14560_ (.A1(_06596_),
    .A2(_06639_),
    .B1(_06638_),
    .X(_06641_));
 sky130_fd_sc_hd__o2bb2a_1 _14561_ (.A1_N(_06640_),
    .A2_N(_06641_),
    .B1(_06596_),
    .B2(_06638_),
    .X(_06642_));
 sky130_fd_sc_hd__o21ba_1 _14562_ (.A1(_06495_),
    .A2(_06533_),
    .B1_N(_06496_),
    .X(_06643_));
 sky130_fd_sc_hd__nor2_1 _14563_ (.A(_06643_),
    .B(_06642_),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_1 _14564_ (.A(_06642_),
    .B(_06643_),
    .Y(_06645_));
 sky130_fd_sc_hd__nand2b_1 _14565_ (.A_N(_06644_),
    .B(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__and2b_1 _14566_ (.A_N(_06553_),
    .B(_06646_),
    .X(_06648_));
 sky130_fd_sc_hd__a211oi_1 _14567_ (.A1(_06539_),
    .A2(_06541_),
    .B1(_06646_),
    .C1(_06536_),
    .Y(_06649_));
 sky130_fd_sc_hd__a2111oi_4 _14568_ (.A1(_06539_),
    .A2(_06541_),
    .B1(_06642_),
    .C1(_06643_),
    .D1(_06536_),
    .Y(_06650_));
 sky130_fd_sc_hd__a21oi_1 _14569_ (.A1(_06553_),
    .A2(_06645_),
    .B1(_06644_),
    .Y(_06651_));
 sky130_fd_sc_hd__o21a_1 _14570_ (.A1(_06553_),
    .A2(_06645_),
    .B1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__a21o_2 _14571_ (.A1(_06553_),
    .A2(_06644_),
    .B1(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__inv_2 _14572_ (.A(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__o2bb2ai_4 _14573_ (.A1_N(_06445_),
    .A2_N(_06546_),
    .B1(_06542_),
    .B2(_06457_),
    .Y(_06655_));
 sky130_fd_sc_hd__o211ai_2 _14574_ (.A1(_06337_),
    .A2(_06442_),
    .B1(_06543_),
    .C1(_06546_),
    .Y(_06656_));
 sky130_fd_sc_hd__o21ai_2 _14575_ (.A1(_06457_),
    .A2(_06542_),
    .B1(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__a31oi_1 _14576_ (.A1(_06445_),
    .A2(_06543_),
    .A3(_06546_),
    .B1(_06545_),
    .Y(_06659_));
 sky130_fd_sc_hd__a2bb2oi_1 _14577_ (.A1_N(_06650_),
    .A2_N(_06652_),
    .B1(_06656_),
    .B2(_06544_),
    .Y(_06660_));
 sky130_fd_sc_hd__o211ai_1 _14578_ (.A1(_06457_),
    .A2(_06542_),
    .B1(_06653_),
    .C1(_06656_),
    .Y(_06661_));
 sky130_fd_sc_hd__o211ai_2 _14579_ (.A1(_06648_),
    .A2(_06649_),
    .B1(_06655_),
    .C1(_06543_),
    .Y(_06662_));
 sky130_fd_sc_hd__and2_1 _14580_ (.A(_06661_),
    .B(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__xor2_1 _14581_ (.A(_06552_),
    .B(_06663_),
    .X(net107));
 sky130_fd_sc_hd__a32o_1 _14582_ (.A1(_02432_),
    .A2(_02237_),
    .A3(_02236_),
    .B1(_02097_),
    .B2(_02356_),
    .X(_06664_));
 sky130_fd_sc_hd__or4_2 _14583_ (.A(_02241_),
    .B(_02355_),
    .C(_02433_),
    .D(_02096_),
    .X(_06665_));
 sky130_fd_sc_hd__o221a_1 _14584_ (.A1(_06598_),
    .A2(_06633_),
    .B1(_06488_),
    .B2(_06491_),
    .C1(_06489_),
    .X(_06666_));
 sky130_fd_sc_hd__a21o_1 _14585_ (.A1(_06598_),
    .A2(_06633_),
    .B1(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__o21ai_1 _14586_ (.A1(_06623_),
    .A2(_06632_),
    .B1(_06624_),
    .Y(_06669_));
 sky130_fd_sc_hd__o21ba_1 _14587_ (.A1(_06627_),
    .A2(_06629_),
    .B1_N(_06628_),
    .X(_06670_));
 sky130_fd_sc_hd__o41a_1 _14588_ (.A1(_01058_),
    .A2(_03319_),
    .A3(_06357_),
    .A4(_06613_),
    .B1(_06612_),
    .X(_06671_));
 sky130_fd_sc_hd__nand2_1 _14589_ (.A(_06670_),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__inv_2 _14590_ (.A(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nor2_1 _14591_ (.A(_06670_),
    .B(_06671_),
    .Y(_06674_));
 sky130_fd_sc_hd__or4_1 _14592_ (.A(_01221_),
    .B(net136),
    .C(_03319_),
    .D(_03652_),
    .X(_06675_));
 sky130_fd_sc_hd__o311a_1 _14593_ (.A1(_01399_),
    .A2(_01404_),
    .A3(_03319_),
    .B1(_03653_),
    .C1(_01222_),
    .X(_06676_));
 sky130_fd_sc_hd__and3_1 _14594_ (.A(_06608_),
    .B(net137),
    .C(_03320_),
    .X(_06677_));
 sky130_fd_sc_hd__nor2_1 _14595_ (.A(_06676_),
    .B(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__a2111oi_1 _14596_ (.A1(_03834_),
    .A2(_06678_),
    .B1(_06608_),
    .C1(_01058_),
    .D1(_03319_),
    .Y(_06680_));
 sky130_fd_sc_hd__o211a_1 _14597_ (.A1(_01058_),
    .A2(_03834_),
    .B1(_06609_),
    .C1(_06678_),
    .X(_06681_));
 sky130_fd_sc_hd__nor2_1 _14598_ (.A(_06680_),
    .B(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__xor2_1 _14599_ (.A(_06604_),
    .B(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__o21ai_1 _14600_ (.A1(_06673_),
    .A2(_06674_),
    .B1(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__or3_1 _14601_ (.A(_06673_),
    .B(_06674_),
    .C(_06683_),
    .X(_06685_));
 sky130_fd_sc_hd__and2_1 _14602_ (.A(_06684_),
    .B(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__nor2_1 _14603_ (.A(_06600_),
    .B(_06618_),
    .Y(_06687_));
 sky130_fd_sc_hd__nor2_1 _14604_ (.A(_06601_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__xor2_1 _14605_ (.A(_06686_),
    .B(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__or4_1 _14606_ (.A(_02049_),
    .B(_02051_),
    .C(_02692_),
    .D(_02694_),
    .X(_06691_));
 sky130_fd_sc_hd__or4_1 _14607_ (.A(_01589_),
    .B(_01822_),
    .C(_02925_),
    .D(_03086_),
    .X(_06692_));
 sky130_fd_sc_hd__o32a_1 _14608_ (.A1(_01589_),
    .A2(net131),
    .A3(net130),
    .B1(_01822_),
    .B2(_02925_),
    .X(_06693_));
 sky130_fd_sc_hd__a31oi_1 _14609_ (.A1(_01823_),
    .A2(_03087_),
    .A3(_06602_),
    .B1(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__xnor2_1 _14610_ (.A(_06691_),
    .B(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__xnor2_1 _14611_ (.A(_06689_),
    .B(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__or2_1 _14612_ (.A(_06669_),
    .B(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__and2_1 _14613_ (.A(_06696_),
    .B(_06669_),
    .X(_06698_));
 sky130_fd_sc_hd__and3_1 _14614_ (.A(_06667_),
    .B(_06669_),
    .C(_06696_),
    .X(_06699_));
 sky130_fd_sc_hd__o21ai_2 _14615_ (.A1(_06698_),
    .A2(_06667_),
    .B1(_06697_),
    .Y(_06700_));
 sky130_fd_sc_hd__o22ai_1 _14616_ (.A1(_06667_),
    .A2(_06697_),
    .B1(_06699_),
    .B2(_06700_),
    .Y(_06702_));
 sky130_fd_sc_hd__a21o_1 _14617_ (.A1(_06664_),
    .A2(_06665_),
    .B1(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__inv_2 _14618_ (.A(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__and3_1 _14619_ (.A(_06702_),
    .B(_06665_),
    .C(_06664_),
    .X(_06705_));
 sky130_fd_sc_hd__or2_1 _14620_ (.A(_06582_),
    .B(_06585_),
    .X(_06706_));
 sky130_fd_sc_hd__and4_1 _14621_ (.A(_01189_),
    .B(_01273_),
    .C(_03450_),
    .D(_03584_),
    .X(_06707_));
 sky130_fd_sc_hd__o32a_1 _14622_ (.A1(_01188_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(_01272_),
    .B2(_03449_),
    .X(_06708_));
 sky130_fd_sc_hd__nor2_1 _14623_ (.A(_06707_),
    .B(_06708_),
    .Y(_06709_));
 sky130_fd_sc_hd__a31o_1 _14624_ (.A1(_01034_),
    .A2(_01036_),
    .A3(net129),
    .B1(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__a21boi_2 _14625_ (.A1(_06569_),
    .A2(_06572_),
    .B1_N(_06571_),
    .Y(_06711_));
 sky130_fd_sc_hd__or4_1 _14626_ (.A(_01037_),
    .B(_03583_),
    .C(_06510_),
    .D(_06711_),
    .X(_06713_));
 sky130_fd_sc_hd__xor2_1 _14627_ (.A(_06583_),
    .B(_06711_),
    .X(_06714_));
 sky130_fd_sc_hd__o32a_1 _14628_ (.A1(_01882_),
    .A2(_02628_),
    .A3(_02630_),
    .B1(_02857_),
    .B2(_01662_),
    .X(_06715_));
 sky130_fd_sc_hd__and4_1 _14629_ (.A(_01664_),
    .B(_01883_),
    .C(_02633_),
    .D(_02858_),
    .X(_06716_));
 sky130_fd_sc_hd__o22ai_1 _14630_ (.A1(_01542_),
    .A2(_03179_),
    .B1(_06715_),
    .B2(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__or4_1 _14631_ (.A(_01542_),
    .B(_03179_),
    .C(_06715_),
    .D(_06716_),
    .X(_06718_));
 sky130_fd_sc_hd__a31o_1 _14632_ (.A1(_01544_),
    .A2(_02858_),
    .A3(_06566_),
    .B1(_06564_),
    .X(_06719_));
 sky130_fd_sc_hd__a21oi_1 _14633_ (.A1(_06717_),
    .A2(_06718_),
    .B1(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__nand3_1 _14634_ (.A(_06717_),
    .B(_06718_),
    .C(_06719_),
    .Y(_06721_));
 sky130_fd_sc_hd__nand2b_1 _14635_ (.A_N(_06720_),
    .B(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__xnor2_1 _14636_ (.A(_06562_),
    .B(_06722_),
    .Y(_06724_));
 sky130_fd_sc_hd__a21o_1 _14637_ (.A1(_06583_),
    .A2(_06711_),
    .B1(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__xor2_1 _14638_ (.A(_06714_),
    .B(_06724_),
    .X(_06726_));
 sky130_fd_sc_hd__o21a_1 _14639_ (.A1(_06558_),
    .A2(_06575_),
    .B1(_06557_),
    .X(_06727_));
 sky130_fd_sc_hd__xnor2_1 _14640_ (.A(_06726_),
    .B(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__xor2_1 _14641_ (.A(_06710_),
    .B(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__and3_1 _14642_ (.A(_06729_),
    .B(_06706_),
    .C(_06580_),
    .X(_06730_));
 sky130_fd_sc_hd__a211o_1 _14643_ (.A1(_06585_),
    .A2(_06580_),
    .B1(_06582_),
    .C1(_06729_),
    .X(_06731_));
 sky130_fd_sc_hd__nand2b_1 _14644_ (.A_N(_06730_),
    .B(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__a21oi_2 _14645_ (.A1(_06595_),
    .A2(_06589_),
    .B1(_06590_),
    .Y(_06733_));
 sky130_fd_sc_hd__xor2_2 _14646_ (.A(_06732_),
    .B(_06733_),
    .X(_06735_));
 sky130_fd_sc_hd__o21ai_1 _14647_ (.A1(_06704_),
    .A2(_06705_),
    .B1(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__or3_1 _14648_ (.A(_06704_),
    .B(_06705_),
    .C(_06735_),
    .X(_06737_));
 sky130_fd_sc_hd__and2_1 _14649_ (.A(_06736_),
    .B(_06737_),
    .X(_06738_));
 sky130_fd_sc_hd__or2_1 _14650_ (.A(_06641_),
    .B(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__o211a_1 _14651_ (.A1(_06596_),
    .A2(_06639_),
    .B1(_06638_),
    .C1(_06738_),
    .X(_06740_));
 sky130_fd_sc_hd__nand2_1 _14652_ (.A(_06738_),
    .B(_06641_),
    .Y(_06741_));
 sky130_fd_sc_hd__nand2_1 _14653_ (.A(_06739_),
    .B(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__and2b_1 _14654_ (.A_N(_06651_),
    .B(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__a211oi_2 _14655_ (.A1(_06553_),
    .A2(_06645_),
    .B1(_06644_),
    .C1(_06742_),
    .Y(_06744_));
 sky130_fd_sc_hd__or2_2 _14656_ (.A(_06743_),
    .B(_06744_),
    .X(_06746_));
 sky130_fd_sc_hd__inv_2 _14657_ (.A(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__o21ai_1 _14658_ (.A1(_06654_),
    .A2(_06659_),
    .B1(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__o2111ai_4 _14659_ (.A1(_06743_),
    .A2(_06744_),
    .B1(_06543_),
    .C1(_06653_),
    .D1(_06655_),
    .Y(_06749_));
 sky130_fd_sc_hd__nand2_1 _14660_ (.A(_06748_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__nand4_2 _14661_ (.A(_06550_),
    .B(_06661_),
    .C(_06662_),
    .D(_06455_),
    .Y(_06751_));
 sky130_fd_sc_hd__a311o_1 _14662_ (.A1(_06663_),
    .A2(_06455_),
    .A3(_06550_),
    .B1(_00834_),
    .C1(_06750_),
    .X(_06752_));
 sky130_fd_sc_hd__a22o_1 _14663_ (.A1(_06748_),
    .A2(_06749_),
    .B1(_06751_),
    .B2(_00845_),
    .X(_06753_));
 sky130_fd_sc_hd__and2_1 _14664_ (.A(_06752_),
    .B(_06753_),
    .X(net108));
 sky130_fd_sc_hd__a21oi_1 _14665_ (.A1(_06703_),
    .A2(_06735_),
    .B1(_06705_),
    .Y(_06754_));
 sky130_fd_sc_hd__or3_1 _14666_ (.A(_02692_),
    .B(_02694_),
    .C(_02241_),
    .X(_06756_));
 sky130_fd_sc_hd__a32o_1 _14667_ (.A1(_02356_),
    .A2(_02427_),
    .A3(_02428_),
    .B1(_02240_),
    .B2(_02697_),
    .X(_06757_));
 sky130_fd_sc_hd__or4_2 _14668_ (.A(_02241_),
    .B(_02355_),
    .C(_02433_),
    .D(_02696_),
    .X(_06758_));
 sky130_fd_sc_hd__a32o_1 _14669_ (.A1(_02093_),
    .A2(_02095_),
    .A3(_02633_),
    .B1(_06757_),
    .B2(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__inv_2 _14670_ (.A(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand4_1 _14671_ (.A(_02097_),
    .B(_02633_),
    .C(_06757_),
    .D(_06758_),
    .Y(_06761_));
 sky130_fd_sc_hd__and3_1 _14672_ (.A(_06665_),
    .B(_06759_),
    .C(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__a21oi_1 _14673_ (.A1(_06759_),
    .A2(_06761_),
    .B1(_06665_),
    .Y(_06763_));
 sky130_fd_sc_hd__or4_1 _14674_ (.A(_02049_),
    .B(_02051_),
    .C(_02920_),
    .D(_02923_),
    .X(_06764_));
 sky130_fd_sc_hd__a211o_1 _14675_ (.A1(_03315_),
    .A2(_03312_),
    .B1(_01822_),
    .C1(_03317_),
    .X(_06765_));
 sky130_fd_sc_hd__a32o_1 _14676_ (.A1(_01590_),
    .A2(_03316_),
    .A3(_03318_),
    .B1(_01823_),
    .B2(_03087_),
    .X(_06767_));
 sky130_fd_sc_hd__o31a_1 _14677_ (.A1(_01589_),
    .A2(_03086_),
    .A3(_06765_),
    .B1(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__xnor2_1 _14678_ (.A(_06764_),
    .B(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__or2_1 _14679_ (.A(_06674_),
    .B(_06683_),
    .X(_06770_));
 sky130_fd_sc_hd__o32a_1 _14680_ (.A1(net136),
    .A2(_03652_),
    .A3(_06606_),
    .B1(_03832_),
    .B2(_01221_),
    .X(_06771_));
 sky130_fd_sc_hd__a21oi_1 _14681_ (.A1(_06604_),
    .A2(_06682_),
    .B1(_06680_),
    .Y(_06772_));
 sky130_fd_sc_hd__o311a_1 _14682_ (.A1(_02053_),
    .A2(_02696_),
    .A3(_06693_),
    .B1(_06772_),
    .C1(_06692_),
    .X(_06773_));
 sky130_fd_sc_hd__inv_2 _14683_ (.A(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__a211o_1 _14684_ (.A1(_06691_),
    .A2(_06692_),
    .B1(_06693_),
    .C1(_06772_),
    .X(_06775_));
 sky130_fd_sc_hd__and3_1 _14685_ (.A(_06774_),
    .B(_06775_),
    .C(_06771_),
    .X(_06776_));
 sky130_fd_sc_hd__a21oi_1 _14686_ (.A1(_06774_),
    .A2(_06775_),
    .B1(_06771_),
    .Y(_06778_));
 sky130_fd_sc_hd__o211a_1 _14687_ (.A1(_06776_),
    .A2(_06778_),
    .B1(_06672_),
    .C1(_06770_),
    .X(_06779_));
 sky130_fd_sc_hd__a2111oi_1 _14688_ (.A1(_06672_),
    .A2(_06683_),
    .B1(_06776_),
    .C1(_06778_),
    .D1(_06674_),
    .Y(_06780_));
 sky130_fd_sc_hd__o21bai_1 _14689_ (.A1(_06769_),
    .A2(_06779_),
    .B1_N(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__o21ai_1 _14690_ (.A1(_06779_),
    .A2(_06780_),
    .B1(_06769_),
    .Y(_06782_));
 sky130_fd_sc_hd__or3_1 _14691_ (.A(_06769_),
    .B(_06779_),
    .C(_06780_),
    .X(_06783_));
 sky130_fd_sc_hd__and2_1 _14692_ (.A(_06782_),
    .B(_06783_),
    .X(_06784_));
 sky130_fd_sc_hd__a21bo_1 _14693_ (.A1(_06686_),
    .A2(_06688_),
    .B1_N(_06695_),
    .X(_06785_));
 sky130_fd_sc_hd__o21a_1 _14694_ (.A1(_06686_),
    .A2(_06688_),
    .B1(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__nand2_1 _14695_ (.A(_06784_),
    .B(_06786_),
    .Y(_06787_));
 sky130_fd_sc_hd__nor2_1 _14696_ (.A(_06784_),
    .B(_06786_),
    .Y(_06789_));
 sky130_fd_sc_hd__a21oi_1 _14697_ (.A1(_06700_),
    .A2(_06787_),
    .B1(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__and2_1 _14698_ (.A(_06790_),
    .B(_06787_),
    .X(_06791_));
 sky130_fd_sc_hd__nand3b_1 _14699_ (.A_N(_06789_),
    .B(_06700_),
    .C(_06787_),
    .Y(_06792_));
 sky130_fd_sc_hd__o21a_1 _14700_ (.A1(_06700_),
    .A2(_06791_),
    .B1(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__nor3_1 _14701_ (.A(_06762_),
    .B(_06763_),
    .C(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__or3_1 _14702_ (.A(_06762_),
    .B(_06763_),
    .C(_06793_),
    .X(_06795_));
 sky130_fd_sc_hd__o21a_1 _14703_ (.A1(_06762_),
    .A2(_06763_),
    .B1(_06793_),
    .X(_06796_));
 sky130_fd_sc_hd__nor2_1 _14704_ (.A(_06794_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__and3_1 _14705_ (.A(_01539_),
    .B(_01541_),
    .C(_03584_),
    .X(_06798_));
 sky130_fd_sc_hd__o32a_1 _14706_ (.A1(_01272_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(_01542_),
    .B2(_03449_),
    .X(_06800_));
 sky130_fd_sc_hd__a31o_1 _14707_ (.A1(_06798_),
    .A2(_03450_),
    .A3(_01273_),
    .B1(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__o21ai_1 _14708_ (.A1(_01188_),
    .A2(_03912_),
    .B1(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__o41a_1 _14709_ (.A1(_01188_),
    .A2(_01272_),
    .A3(_03179_),
    .A4(_03449_),
    .B1(_06721_),
    .X(_06803_));
 sky130_fd_sc_hd__or3b_1 _14710_ (.A(_06720_),
    .B(_06803_),
    .C_N(_06707_),
    .X(_06804_));
 sky130_fd_sc_hd__o21bai_1 _14711_ (.A1(_06720_),
    .A2(_06803_),
    .B1_N(_06707_),
    .Y(_06805_));
 sky130_fd_sc_hd__or4_2 _14712_ (.A(_01658_),
    .B(_01660_),
    .C(_03175_),
    .D(_03177_),
    .X(_06806_));
 sky130_fd_sc_hd__o32ai_1 _14713_ (.A1(_01542_),
    .A2(_03179_),
    .A3(_06715_),
    .B1(_01662_),
    .B2(_02632_),
    .Y(_06807_));
 sky130_fd_sc_hd__or3b_1 _14714_ (.A(_01882_),
    .B(_02857_),
    .C_N(_06807_),
    .X(_06808_));
 sky130_fd_sc_hd__o32a_1 _14715_ (.A1(_01542_),
    .A2(_03179_),
    .A3(_06715_),
    .B1(_01882_),
    .B2(_02857_),
    .X(_06809_));
 sky130_fd_sc_hd__a31o_1 _14716_ (.A1(_01883_),
    .A2(_02858_),
    .A3(_06807_),
    .B1(_06809_),
    .X(_06811_));
 sky130_fd_sc_hd__xnor2_1 _14717_ (.A(_06806_),
    .B(_06811_),
    .Y(_06812_));
 sky130_fd_sc_hd__a21oi_1 _14718_ (.A1(_06804_),
    .A2(_06805_),
    .B1(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__and3_1 _14719_ (.A(_06804_),
    .B(_06805_),
    .C(_06812_),
    .X(_06814_));
 sky130_fd_sc_hd__nor2_1 _14720_ (.A(_06813_),
    .B(_06814_),
    .Y(_06815_));
 sky130_fd_sc_hd__and3_1 _14721_ (.A(_06815_),
    .B(_06725_),
    .C(_06713_),
    .X(_06816_));
 sky130_fd_sc_hd__a21oi_1 _14722_ (.A1(_06713_),
    .A2(_06725_),
    .B1(_06815_),
    .Y(_06817_));
 sky130_fd_sc_hd__or2_1 _14723_ (.A(_06802_),
    .B(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__o21ai_1 _14724_ (.A1(_06816_),
    .A2(_06817_),
    .B1(_06802_),
    .Y(_06819_));
 sky130_fd_sc_hd__o21a_1 _14725_ (.A1(_06816_),
    .A2(_06818_),
    .B1(_06819_),
    .X(_06820_));
 sky130_fd_sc_hd__o21bai_1 _14726_ (.A1(_06726_),
    .A2(_06727_),
    .B1_N(_06710_),
    .Y(_06822_));
 sky130_fd_sc_hd__a21bo_1 _14727_ (.A1(_06726_),
    .A2(_06727_),
    .B1_N(_06822_),
    .X(_06823_));
 sky130_fd_sc_hd__xor2_1 _14728_ (.A(_06820_),
    .B(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__o21ai_1 _14729_ (.A1(_06730_),
    .A2(_06733_),
    .B1(_06731_),
    .Y(_06825_));
 sky130_fd_sc_hd__xor2_2 _14730_ (.A(_06824_),
    .B(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__xnor2_1 _14731_ (.A(_06797_),
    .B(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__xnor2_1 _14732_ (.A(_06754_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__o21a_1 _14733_ (.A1(_06740_),
    .A2(_06651_),
    .B1(_06739_),
    .X(_06829_));
 sky130_fd_sc_hd__and2b_1 _14734_ (.A_N(_06828_),
    .B(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__and2b_1 _14735_ (.A_N(_06829_),
    .B(_06828_),
    .X(_06831_));
 sky130_fd_sc_hd__or2_2 _14736_ (.A(_06830_),
    .B(_06831_),
    .X(_06833_));
 sky130_fd_sc_hd__inv_2 _14737_ (.A(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__nand2_1 _14738_ (.A(_06749_),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__o2111a_1 _14739_ (.A1(_06830_),
    .A2(_06831_),
    .B1(_06543_),
    .C1(_06653_),
    .D1(_06655_),
    .X(_06836_));
 sky130_fd_sc_hd__o2111ai_4 _14740_ (.A1(_06830_),
    .A2(_06831_),
    .B1(_06543_),
    .C1(_06653_),
    .D1(_06655_),
    .Y(_06837_));
 sky130_fd_sc_hd__o2111ai_4 _14741_ (.A1(_06650_),
    .A2(_06652_),
    .B1(_06746_),
    .C1(_06833_),
    .D1(_06657_),
    .Y(_06838_));
 sky130_fd_sc_hd__o21ai_1 _14742_ (.A1(_06747_),
    .A2(_06837_),
    .B1(_06835_),
    .Y(_06839_));
 sky130_fd_sc_hd__a31o_1 _14743_ (.A1(_06551_),
    .A2(_06663_),
    .A3(_06750_),
    .B1(_00834_),
    .X(_06840_));
 sky130_fd_sc_hd__xor2_1 _14744_ (.A(_06839_),
    .B(_06840_),
    .X(net110));
 sky130_fd_sc_hd__o31ai_1 _14745_ (.A1(_01589_),
    .A2(_03086_),
    .A3(_06765_),
    .B1(_06764_),
    .Y(_06841_));
 sky130_fd_sc_hd__and3b_1 _14746_ (.A_N(_06675_),
    .B(_06767_),
    .C(_06841_),
    .X(_06843_));
 sky130_fd_sc_hd__a21boi_1 _14747_ (.A1(_06767_),
    .A2(_06841_),
    .B1_N(_06675_),
    .Y(_06844_));
 sky130_fd_sc_hd__a32o_1 _14748_ (.A1(_01590_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_01823_),
    .B2(_03320_),
    .X(_06845_));
 sky130_fd_sc_hd__or4_1 _14749_ (.A(_01589_),
    .B(_01822_),
    .C(_03319_),
    .D(_03652_),
    .X(_06846_));
 sky130_fd_sc_hd__a22o_1 _14750_ (.A1(net137),
    .A2(_03831_),
    .B1(_06845_),
    .B2(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__o21ai_1 _14751_ (.A1(_06843_),
    .A2(_06844_),
    .B1(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__or3_1 _14752_ (.A(_06847_),
    .B(_06844_),
    .C(_06843_),
    .X(_06849_));
 sky130_fd_sc_hd__and2_1 _14753_ (.A(_06848_),
    .B(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__a21o_1 _14754_ (.A1(_06775_),
    .A2(_06771_),
    .B1(_06773_),
    .X(_06851_));
 sky130_fd_sc_hd__xnor2_1 _14755_ (.A(_06850_),
    .B(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__o21ai_1 _14756_ (.A1(_02053_),
    .A2(_03086_),
    .B1(_06852_),
    .Y(_06854_));
 sky130_fd_sc_hd__or4_1 _14757_ (.A(_02053_),
    .B(net131),
    .C(net130),
    .D(_06852_),
    .X(_06855_));
 sky130_fd_sc_hd__nand2_1 _14758_ (.A(_06854_),
    .B(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__and2_1 _14759_ (.A(_06856_),
    .B(_06781_),
    .X(_06857_));
 sky130_fd_sc_hd__nor2_1 _14760_ (.A(_06781_),
    .B(_06856_),
    .Y(_06858_));
 sky130_fd_sc_hd__o21ai_1 _14761_ (.A1(_06857_),
    .A2(_06858_),
    .B1(_06790_),
    .Y(_06859_));
 sky130_fd_sc_hd__or3_1 _14762_ (.A(_06790_),
    .B(_06857_),
    .C(_06858_),
    .X(_06860_));
 sky130_fd_sc_hd__nand2_1 _14763_ (.A(_06859_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__a32o_1 _14764_ (.A1(_02356_),
    .A2(_02693_),
    .A3(_02695_),
    .B1(_02926_),
    .B2(_02240_),
    .X(_06862_));
 sky130_fd_sc_hd__o31a_1 _14765_ (.A1(_02355_),
    .A2(_02925_),
    .A3(_06756_),
    .B1(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__a21oi_2 _14766_ (.A1(_02432_),
    .A2(_02633_),
    .B1(_06863_),
    .Y(_06865_));
 sky130_fd_sc_hd__and3_1 _14767_ (.A(_02432_),
    .B(_06863_),
    .C(_02633_),
    .X(_06866_));
 sky130_fd_sc_hd__or4b_1 _14768_ (.A(_02433_),
    .B(_02628_),
    .C(_02630_),
    .D_N(_06863_),
    .X(_06867_));
 sky130_fd_sc_hd__o32a_1 _14769_ (.A1(net133),
    .A2(_02094_),
    .A3(_02857_),
    .B1(_06865_),
    .B2(_06866_),
    .X(_06868_));
 sky130_fd_sc_hd__a2111oi_2 _14770_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_06865_),
    .C1(_06866_),
    .D1(_02096_),
    .Y(_06869_));
 sky130_fd_sc_hd__nor3_1 _14771_ (.A(_06758_),
    .B(_06868_),
    .C(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__o21a_1 _14772_ (.A1(_06868_),
    .A2(_06869_),
    .B1(_06758_),
    .X(_06871_));
 sky130_fd_sc_hd__o21ai_1 _14773_ (.A1(_06868_),
    .A2(_06869_),
    .B1(_06758_),
    .Y(_06872_));
 sky130_fd_sc_hd__o21ai_1 _14774_ (.A1(_06665_),
    .A2(_06760_),
    .B1(_06761_),
    .Y(_06873_));
 sky130_fd_sc_hd__o21ai_1 _14775_ (.A1(_06870_),
    .A2(_06871_),
    .B1(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__or3_1 _14776_ (.A(_06870_),
    .B(_06871_),
    .C(_06873_),
    .X(_06876_));
 sky130_fd_sc_hd__and2_1 _14777_ (.A(_06874_),
    .B(_06876_),
    .X(_06877_));
 sky130_fd_sc_hd__nor2_1 _14778_ (.A(_06877_),
    .B(_06861_),
    .Y(_06878_));
 sky130_fd_sc_hd__nand2_1 _14779_ (.A(_06861_),
    .B(_06877_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2b_1 _14780_ (.A_N(_06878_),
    .B(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__o21ba_1 _14781_ (.A1(_06802_),
    .A2(_06817_),
    .B1_N(_06816_),
    .X(_06881_));
 sky130_fd_sc_hd__a21boi_1 _14782_ (.A1(_06804_),
    .A2(_06812_),
    .B1_N(_06805_),
    .Y(_06882_));
 sky130_fd_sc_hd__and3_1 _14783_ (.A(_01664_),
    .B(_03445_),
    .C(_03448_),
    .X(_06883_));
 sky130_fd_sc_hd__a31o_1 _14784_ (.A1(_01883_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_06883_),
    .X(_06884_));
 sky130_fd_sc_hd__and3_1 _14785_ (.A(_06883_),
    .B(_03180_),
    .C(_01883_),
    .X(_06885_));
 sky130_fd_sc_hd__o31a_1 _14786_ (.A1(_01882_),
    .A2(_03449_),
    .A3(_06806_),
    .B1(_06884_),
    .X(_06887_));
 sky130_fd_sc_hd__xor2_1 _14787_ (.A(_06798_),
    .B(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__o21ai_1 _14788_ (.A1(_06806_),
    .A2(_06809_),
    .B1(_06808_),
    .Y(_06889_));
 sky130_fd_sc_hd__a31oi_2 _14789_ (.A1(_01273_),
    .A2(_03450_),
    .A3(_06798_),
    .B1(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__and4_1 _14790_ (.A(_06798_),
    .B(_06889_),
    .C(_01273_),
    .D(_03450_),
    .X(_06891_));
 sky130_fd_sc_hd__o21bai_1 _14791_ (.A1(_06890_),
    .A2(_06891_),
    .B1_N(_06888_),
    .Y(_06892_));
 sky130_fd_sc_hd__or3b_1 _14792_ (.A(_06890_),
    .B(_06891_),
    .C_N(_06888_),
    .X(_06893_));
 sky130_fd_sc_hd__nor2_1 _14793_ (.A(_06888_),
    .B(_06891_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand2_1 _14794_ (.A(_06892_),
    .B(_06893_),
    .Y(_06895_));
 sky130_fd_sc_hd__and2b_1 _14795_ (.A_N(_06882_),
    .B(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__and2b_1 _14796_ (.A_N(_06895_),
    .B(_06882_),
    .X(_06898_));
 sky130_fd_sc_hd__nor2_1 _14797_ (.A(_06896_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__a31o_1 _14798_ (.A1(_01269_),
    .A2(_01271_),
    .A3(net129),
    .B1(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__nor2_1 _14799_ (.A(_06881_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__and2_1 _14800_ (.A(_06881_),
    .B(_06900_),
    .X(_06902_));
 sky130_fd_sc_hd__o221ai_1 _14801_ (.A1(_06820_),
    .A2(_06823_),
    .B1(_06730_),
    .B2(_06733_),
    .C1(_06731_),
    .Y(_06903_));
 sky130_fd_sc_hd__a21bo_1 _14802_ (.A1(_06820_),
    .A2(_06823_),
    .B1_N(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__o21ai_1 _14803_ (.A1(_06901_),
    .A2(_06902_),
    .B1(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__or3_1 _14804_ (.A(_06901_),
    .B(_06902_),
    .C(_06904_),
    .X(_06906_));
 sky130_fd_sc_hd__and2_2 _14805_ (.A(_06905_),
    .B(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__xnor2_1 _14806_ (.A(_06880_),
    .B(_06907_),
    .Y(_06909_));
 sky130_fd_sc_hd__o21a_1 _14807_ (.A1(_06796_),
    .A2(_06826_),
    .B1(_06795_),
    .X(_06910_));
 sky130_fd_sc_hd__nand2_1 _14808_ (.A(_06909_),
    .B(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__nor2_1 _14809_ (.A(_06909_),
    .B(_06910_),
    .Y(_06912_));
 sky130_fd_sc_hd__or2_1 _14810_ (.A(_06909_),
    .B(_06910_),
    .X(_06913_));
 sky130_fd_sc_hd__nand2_2 _14811_ (.A(_06911_),
    .B(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__o221a_1 _14812_ (.A1(_06754_),
    .A2(_06827_),
    .B1(_06740_),
    .B2(_06651_),
    .C1(_06739_),
    .X(_06915_));
 sky130_fd_sc_hd__a21o_2 _14813_ (.A1(_06754_),
    .A2(_06827_),
    .B1(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__xnor2_4 _14814_ (.A(_06914_),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__inv_2 _14815_ (.A(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__a31o_1 _14816_ (.A1(_06660_),
    .A2(_06746_),
    .A3(_06833_),
    .B1(_06918_),
    .X(_06920_));
 sky130_fd_sc_hd__o2111ai_1 _14817_ (.A1(_06650_),
    .A2(_06652_),
    .B1(_06918_),
    .C1(_06833_),
    .D1(_06657_),
    .Y(_06921_));
 sky130_fd_sc_hd__nor3_1 _14818_ (.A(_06747_),
    .B(_06917_),
    .C(_06837_),
    .Y(_06922_));
 sky130_fd_sc_hd__o21ai_2 _14819_ (.A1(_06747_),
    .A2(_06921_),
    .B1(_06920_),
    .Y(_06923_));
 sky130_fd_sc_hd__a221oi_2 _14820_ (.A1(_06748_),
    .A2(_06749_),
    .B1(_06835_),
    .B2(_06838_),
    .C1(_06751_),
    .Y(_06924_));
 sky130_fd_sc_hd__nor2_1 _14821_ (.A(_00834_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__xnor2_1 _14822_ (.A(_06923_),
    .B(_06925_),
    .Y(net111));
 sky130_fd_sc_hd__o21ai_2 _14823_ (.A1(_06912_),
    .A2(_06916_),
    .B1(_06911_),
    .Y(_06926_));
 sky130_fd_sc_hd__or4_1 _14824_ (.A(net133),
    .B(_02094_),
    .C(_03175_),
    .D(_03177_),
    .X(_06927_));
 sky130_fd_sc_hd__or3_1 _14825_ (.A(net131),
    .B(net130),
    .C(_02241_),
    .X(_06928_));
 sky130_fd_sc_hd__and3_1 _14826_ (.A(_03087_),
    .B(_02240_),
    .C(_02356_),
    .X(_06930_));
 sky130_fd_sc_hd__o311a_1 _14827_ (.A1(_02355_),
    .A2(_02920_),
    .A3(_02923_),
    .B1(_03087_),
    .C1(_02240_),
    .X(_06931_));
 sky130_fd_sc_hd__o311a_1 _14828_ (.A1(net131),
    .A2(net130),
    .A3(_02241_),
    .B1(_02356_),
    .C1(_02926_),
    .X(_06932_));
 sky130_fd_sc_hd__a311oi_1 _14829_ (.A1(_02633_),
    .A2(_02693_),
    .A3(_02695_),
    .B1(_06931_),
    .C1(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__a311o_1 _14830_ (.A1(_02633_),
    .A2(_02693_),
    .A3(_02695_),
    .B1(_06931_),
    .C1(_06932_),
    .X(_06934_));
 sky130_fd_sc_hd__o211a_1 _14831_ (.A1(_06931_),
    .A2(_06932_),
    .B1(_02633_),
    .C1(_02697_),
    .X(_06935_));
 sky130_fd_sc_hd__o22a_1 _14832_ (.A1(_02857_),
    .A2(_02433_),
    .B1(_06935_),
    .B2(_06933_),
    .X(_06936_));
 sky130_fd_sc_hd__a2111oi_1 _14833_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_06935_),
    .C1(_02433_),
    .D1(_06933_),
    .Y(_06937_));
 sky130_fd_sc_hd__or2_1 _14834_ (.A(_06936_),
    .B(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__o31a_1 _14835_ (.A1(_02355_),
    .A2(_02925_),
    .A3(_06756_),
    .B1(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__or4_1 _14836_ (.A(_02355_),
    .B(_02925_),
    .C(_06756_),
    .D(_06938_),
    .X(_06941_));
 sky130_fd_sc_hd__and2b_1 _14837_ (.A_N(_06939_),
    .B(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__xor2_1 _14838_ (.A(_06927_),
    .B(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__a31o_1 _14839_ (.A1(_02093_),
    .A2(_02095_),
    .A3(_02858_),
    .B1(_06866_),
    .X(_06944_));
 sky130_fd_sc_hd__or3b_1 _14840_ (.A(_06865_),
    .B(_06943_),
    .C_N(_06944_),
    .X(_06945_));
 sky130_fd_sc_hd__o311a_1 _14841_ (.A1(_02096_),
    .A2(_02857_),
    .A3(_06865_),
    .B1(_06867_),
    .C1(_06943_),
    .X(_06946_));
 sky130_fd_sc_hd__o311ai_1 _14842_ (.A1(_02096_),
    .A2(_02857_),
    .A3(_06865_),
    .B1(_06867_),
    .C1(_06943_),
    .Y(_06947_));
 sky130_fd_sc_hd__nand2_1 _14843_ (.A(_06945_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__a21oi_1 _14844_ (.A1(_06872_),
    .A2(_06873_),
    .B1(_06870_),
    .Y(_06949_));
 sky130_fd_sc_hd__xnor2_1 _14845_ (.A(_06948_),
    .B(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__o21ba_1 _14846_ (.A1(_06790_),
    .A2(_06857_),
    .B1_N(_06858_),
    .X(_06952_));
 sky130_fd_sc_hd__o22a_1 _14847_ (.A1(_02053_),
    .A2(_03319_),
    .B1(_03652_),
    .B2(_01822_),
    .X(_06953_));
 sky130_fd_sc_hd__and4_1 _14848_ (.A(_01823_),
    .B(_02054_),
    .C(_03320_),
    .D(_03653_),
    .X(_06954_));
 sky130_fd_sc_hd__a2bb2o_1 _14849_ (.A1_N(_06953_),
    .A2_N(_06954_),
    .B1(_01590_),
    .B2(_03831_),
    .X(_06955_));
 sky130_fd_sc_hd__o21ba_1 _14850_ (.A1(_06847_),
    .A2(_06843_),
    .B1_N(_06844_),
    .X(_06956_));
 sky130_fd_sc_hd__or2_1 _14851_ (.A(_06955_),
    .B(_06956_),
    .X(_06957_));
 sky130_fd_sc_hd__nand2_1 _14852_ (.A(_06955_),
    .B(_06956_),
    .Y(_06958_));
 sky130_fd_sc_hd__and2_1 _14853_ (.A(_06957_),
    .B(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__xor2_1 _14854_ (.A(_06846_),
    .B(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__o32a_1 _14855_ (.A1(_02053_),
    .A2(net131),
    .A3(net130),
    .B1(_06850_),
    .B2(_06851_),
    .X(_06961_));
 sky130_fd_sc_hd__a211o_1 _14856_ (.A1(_06850_),
    .A2(_06851_),
    .B1(_02053_),
    .C1(_03086_),
    .X(_06963_));
 sky130_fd_sc_hd__a211o_1 _14857_ (.A1(_06850_),
    .A2(_06851_),
    .B1(_06960_),
    .C1(_06961_),
    .X(_06964_));
 sky130_fd_sc_hd__o211a_1 _14858_ (.A1(_06850_),
    .A2(_06851_),
    .B1(_06960_),
    .C1(_06963_),
    .X(_06965_));
 sky130_fd_sc_hd__nand2_1 _14859_ (.A(_06952_),
    .B(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__o21a_1 _14860_ (.A1(_06965_),
    .A2(_06952_),
    .B1(_06964_),
    .X(_06967_));
 sky130_fd_sc_hd__o2bb2a_1 _14861_ (.A1_N(_06966_),
    .A2_N(_06967_),
    .B1(_06952_),
    .B2(_06964_),
    .X(_06968_));
 sky130_fd_sc_hd__xnor2_1 _14862_ (.A(_06950_),
    .B(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__or4_1 _14863_ (.A(_01662_),
    .B(_01882_),
    .C(_03449_),
    .D(_03583_),
    .X(_06970_));
 sky130_fd_sc_hd__o32a_1 _14864_ (.A1(_01662_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(_01882_),
    .B2(_03449_),
    .X(_06971_));
 sky130_fd_sc_hd__a31o_1 _14865_ (.A1(_01883_),
    .A2(_03584_),
    .A3(_06883_),
    .B1(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__o31a_1 _14866_ (.A1(_01538_),
    .A2(_01540_),
    .A3(_03912_),
    .B1(_06972_),
    .X(_06974_));
 sky130_fd_sc_hd__o221a_1 _14867_ (.A1(_01542_),
    .A2(_03912_),
    .B1(_06890_),
    .B2(_06894_),
    .C1(_06972_),
    .X(_06975_));
 sky130_fd_sc_hd__inv_2 _14868_ (.A(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__or3_1 _14869_ (.A(_06890_),
    .B(_06894_),
    .C(_06974_),
    .X(_06977_));
 sky130_fd_sc_hd__a31o_1 _14870_ (.A1(_01544_),
    .A2(_03584_),
    .A3(_06884_),
    .B1(_06885_),
    .X(_06978_));
 sky130_fd_sc_hd__a21oi_1 _14871_ (.A1(_06976_),
    .A2(_06977_),
    .B1(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__and3_1 _14872_ (.A(_06976_),
    .B(_06977_),
    .C(_06978_),
    .X(_06980_));
 sky130_fd_sc_hd__o21bai_1 _14873_ (.A1(_06979_),
    .A2(_06980_),
    .B1_N(_06898_),
    .Y(_06981_));
 sky130_fd_sc_hd__or4b_1 _14874_ (.A(_06895_),
    .B(_06979_),
    .C(_06980_),
    .D_N(_06882_),
    .X(_06982_));
 sky130_fd_sc_hd__o21bai_1 _14875_ (.A1(_06901_),
    .A2(_06904_),
    .B1_N(_06902_),
    .Y(_06983_));
 sky130_fd_sc_hd__a21oi_1 _14876_ (.A1(_06981_),
    .A2(_06982_),
    .B1(_06983_),
    .Y(_06985_));
 sky130_fd_sc_hd__a21o_1 _14877_ (.A1(_06981_),
    .A2(_06983_),
    .B1(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__and2b_1 _14878_ (.A_N(_06969_),
    .B(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__and2b_1 _14879_ (.A_N(_06986_),
    .B(_06969_),
    .X(_06988_));
 sky130_fd_sc_hd__o21a_1 _14880_ (.A1(_06878_),
    .A2(_06907_),
    .B1(_06879_),
    .X(_06989_));
 sky130_fd_sc_hd__nor3_1 _14881_ (.A(_06989_),
    .B(_06988_),
    .C(_06987_),
    .Y(_06990_));
 sky130_fd_sc_hd__o221a_1 _14882_ (.A1(_06878_),
    .A2(_06907_),
    .B1(_06987_),
    .B2(_06988_),
    .C1(_06879_),
    .X(_06991_));
 sky130_fd_sc_hd__o21ba_1 _14883_ (.A1(_06926_),
    .A2(_06991_),
    .B1_N(_06990_),
    .X(_06992_));
 sky130_fd_sc_hd__a21bo_1 _14884_ (.A1(_06926_),
    .A2(_06991_),
    .B1_N(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__o41a_4 _14885_ (.A1(_06926_),
    .A2(_06987_),
    .A3(_06988_),
    .A4(_06989_),
    .B1(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__inv_2 _14886_ (.A(_06994_),
    .Y(_06996_));
 sky130_fd_sc_hd__a41o_1 _14887_ (.A1(_06660_),
    .A2(_06746_),
    .A3(_06833_),
    .A4(_06918_),
    .B1(_06994_),
    .X(_06997_));
 sky130_fd_sc_hd__nand4_1 _14888_ (.A(_06660_),
    .B(_06746_),
    .C(_06833_),
    .D(_06994_),
    .Y(_06998_));
 sky130_fd_sc_hd__nor4_1 _14889_ (.A(_06747_),
    .B(_06917_),
    .C(_06996_),
    .D(_06837_),
    .Y(_06999_));
 sky130_fd_sc_hd__o21ai_2 _14890_ (.A1(_06917_),
    .A2(_06998_),
    .B1(_06997_),
    .Y(_07000_));
 sky130_fd_sc_hd__and4b_1 _14891_ (.A_N(_06751_),
    .B(_06839_),
    .C(_06923_),
    .D(_06750_),
    .X(_07001_));
 sky130_fd_sc_hd__o2bb2a_1 _14892_ (.A1_N(_06923_),
    .A2_N(_06924_),
    .B1(_00812_),
    .B2(_00823_),
    .X(_07002_));
 sky130_fd_sc_hd__xnor2_1 _14893_ (.A(_07000_),
    .B(_07002_),
    .Y(net112));
 sky130_fd_sc_hd__a21o_1 _14894_ (.A1(_06950_),
    .A2(_06968_),
    .B1(_06986_),
    .X(_07003_));
 sky130_fd_sc_hd__o21a_1 _14895_ (.A1(_06950_),
    .A2(_06968_),
    .B1(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__or4_1 _14896_ (.A(_01882_),
    .B(_03581_),
    .C(_03582_),
    .D(_06883_),
    .X(_07006_));
 sky130_fd_sc_hd__or4_1 _14897_ (.A(_00321_),
    .B(net24),
    .C(_03580_),
    .D(_01662_),
    .X(_07007_));
 sky130_fd_sc_hd__a21boi_1 _14898_ (.A1(_06976_),
    .A2(_06978_),
    .B1_N(_06977_),
    .Y(_07008_));
 sky130_fd_sc_hd__o211ai_1 _14899_ (.A1(_01662_),
    .A2(_03912_),
    .B1(_07006_),
    .C1(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__a21o_1 _14900_ (.A1(_07006_),
    .A2(_07007_),
    .B1(_07008_),
    .X(_07010_));
 sky130_fd_sc_hd__nand2_1 _14901_ (.A(_07009_),
    .B(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__a21bo_1 _14902_ (.A1(_06983_),
    .A2(_06981_),
    .B1_N(_06982_),
    .X(_07012_));
 sky130_fd_sc_hd__nand2_1 _14903_ (.A(_07012_),
    .B(_07009_),
    .Y(_07013_));
 sky130_fd_sc_hd__xor2_2 _14904_ (.A(_07011_),
    .B(_07012_),
    .X(_07014_));
 sky130_fd_sc_hd__and3_1 _14905_ (.A(_02054_),
    .B(_03653_),
    .C(_06765_),
    .X(_07015_));
 sky130_fd_sc_hd__a31o_1 _14906_ (.A1(_01820_),
    .A2(_01821_),
    .A3(_03831_),
    .B1(_07015_),
    .X(_07017_));
 sky130_fd_sc_hd__a21bo_1 _14907_ (.A1(_06955_),
    .A2(_06956_),
    .B1_N(_06846_),
    .X(_07018_));
 sky130_fd_sc_hd__a21oi_1 _14908_ (.A1(_06957_),
    .A2(_07018_),
    .B1(_07017_),
    .Y(_07019_));
 sky130_fd_sc_hd__and3_1 _14909_ (.A(_06957_),
    .B(_07017_),
    .C(_07018_),
    .X(_07020_));
 sky130_fd_sc_hd__o221a_1 _14910_ (.A1(_07019_),
    .A2(_07020_),
    .B1(_06965_),
    .B2(_06952_),
    .C1(_06964_),
    .X(_07021_));
 sky130_fd_sc_hd__nor2_1 _14911_ (.A(_07019_),
    .B(_06967_),
    .Y(_07022_));
 sky130_fd_sc_hd__or2_1 _14912_ (.A(_07021_),
    .B(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__o32a_1 _14913_ (.A1(_03175_),
    .A2(_03177_),
    .A3(_02433_),
    .B1(_02696_),
    .B2(_02857_),
    .X(_07024_));
 sky130_fd_sc_hd__and4_1 _14914_ (.A(_02697_),
    .B(_02858_),
    .C(_03180_),
    .D(_02432_),
    .X(_07025_));
 sky130_fd_sc_hd__nor2_1 _14915_ (.A(_07024_),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__and3_1 _14916_ (.A(_06930_),
    .B(_03318_),
    .C(_03316_),
    .X(_07028_));
 sky130_fd_sc_hd__or4_1 _14917_ (.A(_02241_),
    .B(_02355_),
    .C(_03086_),
    .D(_03319_),
    .X(_07029_));
 sky130_fd_sc_hd__a32o_1 _14918_ (.A1(_02356_),
    .A2(_03082_),
    .A3(_03084_),
    .B1(_03320_),
    .B2(_02240_),
    .X(_07030_));
 sky130_fd_sc_hd__a2111oi_1 _14919_ (.A1(_07029_),
    .A2(_07030_),
    .B1(_02632_),
    .C1(_02920_),
    .D1(_02923_),
    .Y(_07031_));
 sky130_fd_sc_hd__o311a_1 _14920_ (.A1(_02632_),
    .A2(_02920_),
    .A3(_02923_),
    .B1(_07029_),
    .C1(_07030_),
    .X(_07032_));
 sky130_fd_sc_hd__or2_1 _14921_ (.A(_07031_),
    .B(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__xnor2_1 _14922_ (.A(_07026_),
    .B(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__or4_1 _14923_ (.A(_02355_),
    .B(_02925_),
    .C(_06928_),
    .D(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__o31ai_1 _14924_ (.A1(_02355_),
    .A2(_02925_),
    .A3(_06928_),
    .B1(_07034_),
    .Y(_07036_));
 sky130_fd_sc_hd__a31o_1 _14925_ (.A1(_02432_),
    .A2(_02854_),
    .A3(_02856_),
    .B1(_06935_),
    .X(_07037_));
 sky130_fd_sc_hd__a22o_1 _14926_ (.A1(_07035_),
    .A2(_07036_),
    .B1(_07037_),
    .B2(_06934_),
    .X(_07039_));
 sky130_fd_sc_hd__nand4_1 _14927_ (.A(_06934_),
    .B(_07035_),
    .C(_07036_),
    .D(_07037_),
    .Y(_07040_));
 sky130_fd_sc_hd__and4_1 _14928_ (.A(_02097_),
    .B(_03450_),
    .C(_07039_),
    .D(_07040_),
    .X(_07041_));
 sky130_fd_sc_hd__a22oi_1 _14929_ (.A1(_02097_),
    .A2(_03450_),
    .B1(_07039_),
    .B2(_07040_),
    .Y(_07042_));
 sky130_fd_sc_hd__nor2_1 _14930_ (.A(_07041_),
    .B(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__o21ai_1 _14931_ (.A1(_06927_),
    .A2(_06939_),
    .B1(_06941_),
    .Y(_07044_));
 sky130_fd_sc_hd__or2_1 _14932_ (.A(_07043_),
    .B(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__nand2_1 _14933_ (.A(_07043_),
    .B(_07044_),
    .Y(_07046_));
 sky130_fd_sc_hd__a21oi_1 _14934_ (.A1(_06945_),
    .A2(_06949_),
    .B1(_06946_),
    .Y(_07047_));
 sky130_fd_sc_hd__a21oi_1 _14935_ (.A1(_07045_),
    .A2(_07046_),
    .B1(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__and3_1 _14936_ (.A(_07045_),
    .B(_07046_),
    .C(_07047_),
    .X(_07050_));
 sky130_fd_sc_hd__or4_1 _14937_ (.A(_07021_),
    .B(_07022_),
    .C(_07048_),
    .D(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__nor2_1 _14938_ (.A(_07014_),
    .B(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__o22a_1 _14939_ (.A1(_07021_),
    .A2(_07022_),
    .B1(_07048_),
    .B2(_07050_),
    .X(_07053_));
 sky130_fd_sc_hd__o32a_1 _14940_ (.A1(_07023_),
    .A2(_07048_),
    .A3(_07050_),
    .B1(_07014_),
    .B2(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__a2bb2o_1 _14941_ (.A1_N(_07052_),
    .A2_N(_07054_),
    .B1(_07053_),
    .B2(_07014_),
    .X(_07055_));
 sky130_fd_sc_hd__nor2_1 _14942_ (.A(_07004_),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand2_1 _14943_ (.A(_07004_),
    .B(_07055_),
    .Y(_07057_));
 sky130_fd_sc_hd__and2b_1 _14944_ (.A_N(_07056_),
    .B(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__xnor2_1 _14945_ (.A(_06992_),
    .B(_07058_),
    .Y(_07059_));
 sky130_fd_sc_hd__inv_2 _14946_ (.A(_07059_),
    .Y(_07061_));
 sky130_fd_sc_hd__a41oi_1 _14947_ (.A1(_06836_),
    .A2(_06918_),
    .A3(_06994_),
    .A4(_06746_),
    .B1(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__nor4_1 _14948_ (.A(_06917_),
    .B(_06996_),
    .C(_07059_),
    .D(_06838_),
    .Y(_07063_));
 sky130_fd_sc_hd__or2_1 _14949_ (.A(_07062_),
    .B(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__a31o_1 _14950_ (.A1(_06924_),
    .A2(_07000_),
    .A3(_06923_),
    .B1(_00834_),
    .X(_07065_));
 sky130_fd_sc_hd__xor2_1 _14951_ (.A(_07064_),
    .B(_07065_),
    .X(net113));
 sky130_fd_sc_hd__a21oi_2 _14952_ (.A1(_06992_),
    .A2(_07057_),
    .B1(_07056_),
    .Y(_07066_));
 sky130_fd_sc_hd__o2111a_2 _14953_ (.A1(_01882_),
    .A2(_03912_),
    .B1(_06970_),
    .C1(_07010_),
    .D1(_07013_),
    .X(_07067_));
 sky130_fd_sc_hd__a2111o_1 _14954_ (.A1(_02054_),
    .A2(_03831_),
    .B1(_06954_),
    .C1(_07020_),
    .D1(_07022_),
    .X(_07068_));
 sky130_fd_sc_hd__and3_1 _14955_ (.A(_02633_),
    .B(_02926_),
    .C(_07030_),
    .X(_07069_));
 sky130_fd_sc_hd__or3_1 _14956_ (.A(_07025_),
    .B(_07028_),
    .C(_07069_),
    .X(_07071_));
 sky130_fd_sc_hd__o21ai_1 _14957_ (.A1(_07028_),
    .A2(_07069_),
    .B1(_07025_),
    .Y(_07072_));
 sky130_fd_sc_hd__and3_1 _14958_ (.A(_02858_),
    .B(_02922_),
    .C(_02924_),
    .X(_07073_));
 sky130_fd_sc_hd__or3_1 _14959_ (.A(_02353_),
    .B(_02354_),
    .C(_03319_),
    .X(_07074_));
 sky130_fd_sc_hd__a22o_1 _14960_ (.A1(_02238_),
    .A2(_02239_),
    .B1(_03647_),
    .B2(_03648_),
    .X(_07075_));
 sky130_fd_sc_hd__xnor2_1 _14961_ (.A(_07074_),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__and4b_1 _14962_ (.A_N(_07076_),
    .B(_03084_),
    .C(_03082_),
    .D(_02633_),
    .X(_07077_));
 sky130_fd_sc_hd__or4_1 _14963_ (.A(_02632_),
    .B(net131),
    .C(net130),
    .D(_07076_),
    .X(_07078_));
 sky130_fd_sc_hd__o21ai_2 _14964_ (.A1(_02632_),
    .A2(_03086_),
    .B1(_07076_),
    .Y(_07079_));
 sky130_fd_sc_hd__a32o_1 _14965_ (.A1(_02858_),
    .A2(_02922_),
    .A3(_02924_),
    .B1(_07078_),
    .B2(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__or4b_1 _14966_ (.A(_02857_),
    .B(_02925_),
    .C(_07077_),
    .D_N(_07079_),
    .X(_07082_));
 sky130_fd_sc_hd__nand2_1 _14967_ (.A(_07080_),
    .B(_07082_),
    .Y(_07083_));
 sky130_fd_sc_hd__a21o_1 _14968_ (.A1(_07071_),
    .A2(_07072_),
    .B1(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__inv_2 _14969_ (.A(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__and3_1 _14970_ (.A(_07083_),
    .B(_07072_),
    .C(_07071_),
    .X(_07086_));
 sky130_fd_sc_hd__a22o_1 _14971_ (.A1(_06930_),
    .A2(_02926_),
    .B1(_07033_),
    .B2(_07026_),
    .X(_07087_));
 sky130_fd_sc_hd__o21a_1 _14972_ (.A1(_07026_),
    .A2(_07033_),
    .B1(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__nor3_1 _14973_ (.A(_07088_),
    .B(_07086_),
    .C(_07085_),
    .Y(_07089_));
 sky130_fd_sc_hd__o221a_1 _14974_ (.A1(_07026_),
    .A2(_07033_),
    .B1(_07085_),
    .B2(_07086_),
    .C1(_07087_),
    .X(_07090_));
 sky130_fd_sc_hd__and3_1 _14975_ (.A(_02432_),
    .B(_03445_),
    .C(_03448_),
    .X(_07091_));
 sky130_fd_sc_hd__o32a_1 _14976_ (.A1(_03444_),
    .A2(_03447_),
    .A3(_02433_),
    .B1(_02696_),
    .B2(_03179_),
    .X(_07093_));
 sky130_fd_sc_hd__a31o_1 _14977_ (.A1(_02697_),
    .A2(_03176_),
    .A3(_03178_),
    .B1(_07091_),
    .X(_07094_));
 sky130_fd_sc_hd__and3_1 _14978_ (.A(_07091_),
    .B(_03180_),
    .C(_02697_),
    .X(_07095_));
 sky130_fd_sc_hd__o32a_1 _14979_ (.A1(_02096_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(_07093_),
    .B2(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__or4_1 _14980_ (.A(_02096_),
    .B(_03583_),
    .C(_07093_),
    .D(_07095_),
    .X(_07097_));
 sky130_fd_sc_hd__and2b_1 _14981_ (.A_N(_07096_),
    .B(_07097_),
    .X(_07098_));
 sky130_fd_sc_hd__o21ai_1 _14982_ (.A1(_07089_),
    .A2(_07090_),
    .B1(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__or3_1 _14983_ (.A(_07089_),
    .B(_07090_),
    .C(_07098_),
    .X(_07100_));
 sky130_fd_sc_hd__nand2_1 _14984_ (.A(_07099_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__o21ai_1 _14985_ (.A1(_02096_),
    .A2(_03449_),
    .B1(_07040_),
    .Y(_07102_));
 sky130_fd_sc_hd__and3_1 _14986_ (.A(_07101_),
    .B(_07102_),
    .C(_07039_),
    .X(_07104_));
 sky130_fd_sc_hd__a21o_1 _14987_ (.A1(_07039_),
    .A2(_07102_),
    .B1(_07101_),
    .X(_07105_));
 sky130_fd_sc_hd__nand2b_1 _14988_ (.A_N(_07104_),
    .B(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__a21bo_1 _14989_ (.A1(_07045_),
    .A2(_07047_),
    .B1_N(_07046_),
    .X(_07107_));
 sky130_fd_sc_hd__xnor2_1 _14990_ (.A(_07106_),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__or2_1 _14991_ (.A(_07068_),
    .B(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__nand2_1 _14992_ (.A(_07068_),
    .B(_07108_),
    .Y(_07110_));
 sky130_fd_sc_hd__nand2_1 _14993_ (.A(_07110_),
    .B(_07067_),
    .Y(_07111_));
 sky130_fd_sc_hd__nand3_2 _14994_ (.A(_07109_),
    .B(_07110_),
    .C(_07067_),
    .Y(_07112_));
 sky130_fd_sc_hd__a21o_1 _14995_ (.A1(_07109_),
    .A2(_07110_),
    .B1(_07067_),
    .X(_07113_));
 sky130_fd_sc_hd__a221o_1 _14996_ (.A1(_07014_),
    .A2(_07051_),
    .B1(_07112_),
    .B2(_07113_),
    .C1(_07053_),
    .X(_07115_));
 sky130_fd_sc_hd__and4_1 _14997_ (.A(_07066_),
    .B(_07112_),
    .C(_07113_),
    .D(_07054_),
    .X(_07116_));
 sky130_fd_sc_hd__a32oi_4 _14998_ (.A1(_07054_),
    .A2(_07112_),
    .A3(_07113_),
    .B1(_07115_),
    .B2(_07066_),
    .Y(_07117_));
 sky130_fd_sc_hd__o22ai_1 _14999_ (.A1(_07066_),
    .A2(_07115_),
    .B1(_07116_),
    .B2(_07117_),
    .Y(_07118_));
 sky130_fd_sc_hd__a31o_1 _15000_ (.A1(_06922_),
    .A2(_06994_),
    .A3(_07061_),
    .B1(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__and2_2 _15001_ (.A(_07118_),
    .B(_07061_),
    .X(_07120_));
 sky130_fd_sc_hd__inv_2 _15002_ (.A(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__nor4_1 _15003_ (.A(_06917_),
    .B(_06996_),
    .C(_07121_),
    .D(_06838_),
    .Y(_07122_));
 sky130_fd_sc_hd__nand4b_4 _15004_ (.A_N(_06838_),
    .B(_06918_),
    .C(_06994_),
    .D(_07120_),
    .Y(_07123_));
 sky130_fd_sc_hd__nand2_2 _15005_ (.A(_07119_),
    .B(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__o2111a_1 _15006_ (.A1(_07062_),
    .A2(_07063_),
    .B1(_06923_),
    .C1(_07000_),
    .D1(_06924_),
    .X(_07126_));
 sky130_fd_sc_hd__o2bb2a_1 _15007_ (.A1_N(_07119_),
    .A2_N(_07123_),
    .B1(_07126_),
    .B2(_00834_),
    .X(_07127_));
 sky130_fd_sc_hd__a311oi_1 _15008_ (.A1(_07001_),
    .A2(_07064_),
    .A3(_07000_),
    .B1(_07124_),
    .C1(_00834_),
    .Y(_07128_));
 sky130_fd_sc_hd__nor2_1 _15009_ (.A(_07127_),
    .B(_07128_),
    .Y(net114));
 sky130_fd_sc_hd__a21oi_1 _15010_ (.A1(_07105_),
    .A2(_07107_),
    .B1(_07104_),
    .Y(_07129_));
 sky130_fd_sc_hd__o21ba_1 _15011_ (.A1(_07090_),
    .A2(_07098_),
    .B1_N(_07089_),
    .X(_07130_));
 sky130_fd_sc_hd__o32a_1 _15012_ (.A1(_03582_),
    .A2(_02433_),
    .A3(_03581_),
    .B1(_02696_),
    .B2(_03449_),
    .X(_07131_));
 sky130_fd_sc_hd__a31o_1 _15013_ (.A1(_02697_),
    .A2(_03584_),
    .A3(_07091_),
    .B1(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__o21ai_2 _15014_ (.A1(_02096_),
    .A2(_03912_),
    .B1(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__a31o_1 _15015_ (.A1(_02097_),
    .A2(_03584_),
    .A3(_07094_),
    .B1(_07095_),
    .X(_07134_));
 sky130_fd_sc_hd__a31o_1 _15016_ (.A1(_02858_),
    .A2(_02926_),
    .A3(_07079_),
    .B1(_07077_),
    .X(_07136_));
 sky130_fd_sc_hd__nand2_1 _15017_ (.A(_07136_),
    .B(_07134_),
    .Y(_07137_));
 sky130_fd_sc_hd__a311o_1 _15018_ (.A1(_02858_),
    .A2(_02926_),
    .A3(_07079_),
    .B1(_07134_),
    .C1(_07077_),
    .X(_07138_));
 sky130_fd_sc_hd__or4_1 _15019_ (.A(_02857_),
    .B(_02925_),
    .C(_03086_),
    .D(_03179_),
    .X(_07139_));
 sky130_fd_sc_hd__o32a_1 _15020_ (.A1(_02857_),
    .A2(net131),
    .A3(net130),
    .B1(_03179_),
    .B2(_02925_),
    .X(_07140_));
 sky130_fd_sc_hd__a31o_1 _15021_ (.A1(_03087_),
    .A2(_03180_),
    .A3(_07073_),
    .B1(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__o32a_1 _15022_ (.A1(_02353_),
    .A2(_02354_),
    .A3(_03652_),
    .B1(_03319_),
    .B2(_02632_),
    .X(_07142_));
 sky130_fd_sc_hd__or3_1 _15023_ (.A(_02628_),
    .B(_02630_),
    .C(_03652_),
    .X(_07143_));
 sky130_fd_sc_hd__and4_1 _15024_ (.A(_02356_),
    .B(_02633_),
    .C(_03320_),
    .D(_03653_),
    .X(_07144_));
 sky130_fd_sc_hd__o22a_1 _15025_ (.A1(_02241_),
    .A2(_03832_),
    .B1(_07142_),
    .B2(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__xor2_1 _15026_ (.A(_07141_),
    .B(_07145_),
    .X(_07147_));
 sky130_fd_sc_hd__o31a_1 _15027_ (.A1(_02241_),
    .A2(_03652_),
    .A3(_07074_),
    .B1(_07147_),
    .X(_07148_));
 sky130_fd_sc_hd__or4_1 _15028_ (.A(_02241_),
    .B(_03652_),
    .C(_07074_),
    .D(_07147_),
    .X(_07149_));
 sky130_fd_sc_hd__and2b_1 _15029_ (.A_N(_07148_),
    .B(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__a21oi_1 _15030_ (.A1(_07137_),
    .A2(_07138_),
    .B1(_07150_),
    .Y(_07151_));
 sky130_fd_sc_hd__and3_1 _15031_ (.A(_07137_),
    .B(_07138_),
    .C(_07150_),
    .X(_07152_));
 sky130_fd_sc_hd__or2_1 _15032_ (.A(_07151_),
    .B(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__a21bo_1 _15033_ (.A1(_07083_),
    .A2(_07072_),
    .B1_N(_07071_),
    .X(_07154_));
 sky130_fd_sc_hd__nand2b_1 _15034_ (.A_N(_07153_),
    .B(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__and2b_1 _15035_ (.A_N(_07154_),
    .B(_07153_),
    .X(_07156_));
 sky130_fd_sc_hd__inv_2 _15036_ (.A(_07156_),
    .Y(_07158_));
 sky130_fd_sc_hd__nand3_1 _15037_ (.A(_07133_),
    .B(_07155_),
    .C(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__a21o_1 _15038_ (.A1(_07155_),
    .A2(_07158_),
    .B1(_07133_),
    .X(_07160_));
 sky130_fd_sc_hd__a21oi_1 _15039_ (.A1(_07159_),
    .A2(_07160_),
    .B1(_07130_),
    .Y(_07161_));
 sky130_fd_sc_hd__nand3_1 _15040_ (.A(_07130_),
    .B(_07159_),
    .C(_07160_),
    .Y(_07162_));
 sky130_fd_sc_hd__inv_2 _15041_ (.A(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__o21a_1 _15042_ (.A1(_07161_),
    .A2(_07129_),
    .B1(_07162_),
    .X(_07164_));
 sky130_fd_sc_hd__or3_1 _15043_ (.A(_07161_),
    .B(_07163_),
    .C(_07129_),
    .X(_07165_));
 sky130_fd_sc_hd__o21ai_1 _15044_ (.A1(_07161_),
    .A2(_07163_),
    .B1(_07129_),
    .Y(_07166_));
 sky130_fd_sc_hd__a22o_1 _15045_ (.A1(_07109_),
    .A2(_07111_),
    .B1(_07165_),
    .B2(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__nand4_1 _15046_ (.A(_07109_),
    .B(_07111_),
    .C(_07165_),
    .D(_07166_),
    .Y(_07169_));
 sky130_fd_sc_hd__a21oi_2 _15047_ (.A1(_07167_),
    .A2(_07169_),
    .B1(_07117_),
    .Y(_07170_));
 sky130_fd_sc_hd__and3_1 _15048_ (.A(_07117_),
    .B(_07167_),
    .C(_07169_),
    .X(_07171_));
 sky130_fd_sc_hd__nor2_2 _15049_ (.A(_07170_),
    .B(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__a31o_1 _15050_ (.A1(_06922_),
    .A2(_06994_),
    .A3(_07120_),
    .B1(_07172_),
    .X(_07173_));
 sky130_fd_sc_hd__and3_1 _15051_ (.A(_06999_),
    .B(_07120_),
    .C(_07172_),
    .X(_07174_));
 sky130_fd_sc_hd__nand2_1 _15052_ (.A(_07122_),
    .B(_07172_),
    .Y(_07175_));
 sky130_fd_sc_hd__nand2_1 _15053_ (.A(_07173_),
    .B(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__a41o_1 _15054_ (.A1(_07001_),
    .A2(_07064_),
    .A3(_07124_),
    .A4(_07000_),
    .B1(_00834_),
    .X(_07177_));
 sky130_fd_sc_hd__xor2_1 _15055_ (.A(_07176_),
    .B(_07177_),
    .X(net115));
 sky130_fd_sc_hd__o21a_1 _15056_ (.A1(_07133_),
    .A2(_07156_),
    .B1(_07155_),
    .X(_07179_));
 sky130_fd_sc_hd__or4_1 _15057_ (.A(_02696_),
    .B(_03581_),
    .C(_03582_),
    .D(_07139_),
    .X(_07180_));
 sky130_fd_sc_hd__a32o_1 _15058_ (.A1(_07073_),
    .A2(_03180_),
    .A3(_03087_),
    .B1(_02697_),
    .B2(_03584_),
    .X(_07181_));
 sky130_fd_sc_hd__a22o_2 _15059_ (.A1(_02432_),
    .A2(net129),
    .B1(_07180_),
    .B2(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__nand2_1 _15060_ (.A(_07137_),
    .B(_07150_),
    .Y(_07183_));
 sky130_fd_sc_hd__a211o_1 _15061_ (.A1(_07145_),
    .A2(_07141_),
    .B1(_07075_),
    .C1(_07074_),
    .X(_07184_));
 sky130_fd_sc_hd__o21ai_1 _15062_ (.A1(_07141_),
    .A2(_07145_),
    .B1(_07184_),
    .Y(_07185_));
 sky130_fd_sc_hd__a31o_1 _15063_ (.A1(_02697_),
    .A2(_03584_),
    .A3(_07091_),
    .B1(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__inv_2 _15064_ (.A(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__and4_1 _15065_ (.A(_07091_),
    .B(_07185_),
    .C(_02697_),
    .D(_03584_),
    .X(_07188_));
 sky130_fd_sc_hd__and4_1 _15066_ (.A(_02926_),
    .B(_03087_),
    .C(_03180_),
    .D(_03450_),
    .X(_07190_));
 sky130_fd_sc_hd__or4_1 _15067_ (.A(_02925_),
    .B(_03086_),
    .C(_03179_),
    .D(_03449_),
    .X(_07191_));
 sky130_fd_sc_hd__o32a_1 _15068_ (.A1(net131),
    .A2(net130),
    .A3(_03179_),
    .B1(_03449_),
    .B2(_02925_),
    .X(_07192_));
 sky130_fd_sc_hd__a221o_4 _15069_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_03312_),
    .B2(_03315_),
    .C1(_03317_),
    .X(_07193_));
 sky130_fd_sc_hd__xnor2_1 _15070_ (.A(_07143_),
    .B(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__or4_1 _15071_ (.A(_03830_),
    .B(_02353_),
    .C(_03645_),
    .D(_02354_),
    .X(_07195_));
 sky130_fd_sc_hd__a211oi_1 _15072_ (.A1(_07194_),
    .A2(_07195_),
    .B1(_07190_),
    .C1(_07192_),
    .Y(_07196_));
 sky130_fd_sc_hd__o221a_1 _15073_ (.A1(_02355_),
    .A2(_03834_),
    .B1(_07190_),
    .B2(_07192_),
    .C1(_07194_),
    .X(_07197_));
 sky130_fd_sc_hd__nor3_1 _15074_ (.A(_07144_),
    .B(_07196_),
    .C(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__o21a_1 _15075_ (.A1(_07196_),
    .A2(_07197_),
    .B1(_07144_),
    .X(_07199_));
 sky130_fd_sc_hd__or2_1 _15076_ (.A(_07198_),
    .B(_07199_),
    .X(_07201_));
 sky130_fd_sc_hd__o22a_1 _15077_ (.A1(_07187_),
    .A2(_07188_),
    .B1(_07198_),
    .B2(_07199_),
    .X(_07202_));
 sky130_fd_sc_hd__nor2_1 _15078_ (.A(_07188_),
    .B(_07201_),
    .Y(_07203_));
 sky130_fd_sc_hd__a21o_1 _15079_ (.A1(_07203_),
    .A2(_07186_),
    .B1(_07202_),
    .X(_07204_));
 sky130_fd_sc_hd__a221o_2 _15080_ (.A1(_07138_),
    .A2(_07183_),
    .B1(_07203_),
    .B2(_07186_),
    .C1(_07202_),
    .X(_07205_));
 sky130_fd_sc_hd__o211ai_2 _15081_ (.A1(_07134_),
    .A2(_07136_),
    .B1(_07183_),
    .C1(_07204_),
    .Y(_07206_));
 sky130_fd_sc_hd__a21oi_1 _15082_ (.A1(_07205_),
    .A2(_07206_),
    .B1(_07182_),
    .Y(_07207_));
 sky130_fd_sc_hd__a21boi_4 _15083_ (.A1(_07182_),
    .A2(_07205_),
    .B1_N(_07206_),
    .Y(_07208_));
 sky130_fd_sc_hd__a31oi_2 _15084_ (.A1(_07182_),
    .A2(_07205_),
    .A3(_07206_),
    .B1(_07207_),
    .Y(_07209_));
 sky130_fd_sc_hd__o211a_1 _15085_ (.A1(_07133_),
    .A2(_07156_),
    .B1(_07155_),
    .C1(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__nand2_1 _15086_ (.A(_07209_),
    .B(_07179_),
    .Y(_07212_));
 sky130_fd_sc_hd__nor2_1 _15087_ (.A(_07179_),
    .B(_07209_),
    .Y(_07213_));
 sky130_fd_sc_hd__nor2_1 _15088_ (.A(_07210_),
    .B(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__xnor2_1 _15089_ (.A(_07164_),
    .B(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__a21boi_1 _15090_ (.A1(_07117_),
    .A2(_07167_),
    .B1_N(_07169_),
    .Y(_07216_));
 sky130_fd_sc_hd__nand2b_1 _15091_ (.A_N(_07215_),
    .B(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__and2b_2 _15092_ (.A_N(_07216_),
    .B(_07215_),
    .X(_07218_));
 sky130_fd_sc_hd__inv_2 _15093_ (.A(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__and2_2 _15094_ (.A(_07217_),
    .B(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__inv_2 _15095_ (.A(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__and4_1 _15096_ (.A(_06999_),
    .B(_07120_),
    .C(_07172_),
    .D(_07220_),
    .X(_07223_));
 sky130_fd_sc_hd__a41o_1 _15097_ (.A1(_06922_),
    .A2(_06994_),
    .A3(_07120_),
    .A4(_07172_),
    .B1(_07220_),
    .X(_07224_));
 sky130_fd_sc_hd__o41ai_4 _15098_ (.A1(_07170_),
    .A2(_07171_),
    .A3(_07221_),
    .A4(_07123_),
    .B1(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__a31oi_1 _15099_ (.A1(_07126_),
    .A2(_07176_),
    .A3(_07124_),
    .B1(_00834_),
    .Y(_07226_));
 sky130_fd_sc_hd__xnor2_1 _15100_ (.A(_07225_),
    .B(_07226_),
    .Y(net116));
 sky130_fd_sc_hd__o21bai_1 _15101_ (.A1(_07144_),
    .A2(_07196_),
    .B1_N(_07197_),
    .Y(_07227_));
 sky130_fd_sc_hd__nand2_1 _15102_ (.A(_07227_),
    .B(_07180_),
    .Y(_07228_));
 sky130_fd_sc_hd__or4_1 _15103_ (.A(_02696_),
    .B(_03583_),
    .C(_07139_),
    .D(_07227_),
    .X(_07229_));
 sky130_fd_sc_hd__a32o_1 _15104_ (.A1(_02858_),
    .A2(_03650_),
    .A3(_03651_),
    .B1(_03180_),
    .B2(_03320_),
    .X(_07230_));
 sky130_fd_sc_hd__o31ai_1 _15105_ (.A1(_03179_),
    .A2(_03652_),
    .A3(_07193_),
    .B1(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__o221a_1 _15106_ (.A1(_03834_),
    .A2(_02632_),
    .B1(_07193_),
    .B2(_07143_),
    .C1(_07231_),
    .X(_07233_));
 sky130_fd_sc_hd__a2111oi_2 _15107_ (.A1(_03834_),
    .A2(_07231_),
    .B1(_07193_),
    .C1(_02632_),
    .D1(_03652_),
    .Y(_07234_));
 sky130_fd_sc_hd__o21ai_1 _15108_ (.A1(_07233_),
    .A2(_07234_),
    .B1(_07190_),
    .Y(_07235_));
 sky130_fd_sc_hd__o31ai_1 _15109_ (.A1(_07190_),
    .A2(_07233_),
    .A3(_07234_),
    .B1(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__and3_1 _15110_ (.A(_07228_),
    .B(_07229_),
    .C(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__a21oi_1 _15111_ (.A1(_07228_),
    .A2(_07229_),
    .B1(_07236_),
    .Y(_07238_));
 sky130_fd_sc_hd__o311ai_2 _15112_ (.A1(_07190_),
    .A2(_07233_),
    .A3(_07234_),
    .B1(_07235_),
    .C1(_07229_),
    .Y(_07239_));
 sky130_fd_sc_hd__or2_1 _15113_ (.A(_07237_),
    .B(_07238_),
    .X(_07240_));
 sky130_fd_sc_hd__o21a_1 _15114_ (.A1(_07187_),
    .A2(_07203_),
    .B1(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__or3_1 _15115_ (.A(_07187_),
    .B(_07203_),
    .C(_07240_),
    .X(_07242_));
 sky130_fd_sc_hd__nand2b_2 _15116_ (.A_N(_07241_),
    .B(_07242_),
    .Y(_07244_));
 sky130_fd_sc_hd__or4_1 _15117_ (.A(_02925_),
    .B(_03086_),
    .C(_03449_),
    .D(_03583_),
    .X(_07245_));
 sky130_fd_sc_hd__a32o_1 _15118_ (.A1(_03087_),
    .A2(_03445_),
    .A3(_03448_),
    .B1(_03584_),
    .B2(_02926_),
    .X(_07246_));
 sky130_fd_sc_hd__o2bb2a_2 _15119_ (.A1_N(_07245_),
    .A2_N(_07246_),
    .B1(_02696_),
    .B2(_03912_),
    .X(_07247_));
 sky130_fd_sc_hd__xnor2_4 _15120_ (.A(_07244_),
    .B(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__xor2_2 _15121_ (.A(_07208_),
    .B(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__a21oi_2 _15122_ (.A1(_07164_),
    .A2(_07212_),
    .B1(_07213_),
    .Y(_07250_));
 sky130_fd_sc_hd__xnor2_4 _15123_ (.A(_07249_),
    .B(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__inv_2 _15124_ (.A(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__nor2_1 _15125_ (.A(_07251_),
    .B(_07219_),
    .Y(_07253_));
 sky130_fd_sc_hd__xnor2_4 _15126_ (.A(_07218_),
    .B(_07251_),
    .Y(_07255_));
 sky130_fd_sc_hd__a41oi_2 _15127_ (.A1(_06999_),
    .A2(_07120_),
    .A3(_07172_),
    .A4(_07220_),
    .B1(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand4_1 _15128_ (.A(_07122_),
    .B(_07172_),
    .C(_07220_),
    .D(_07255_),
    .Y(_07257_));
 sky130_fd_sc_hd__a41oi_4 _15129_ (.A1(_07174_),
    .A2(_07217_),
    .A3(_07219_),
    .A4(_07252_),
    .B1(_07256_),
    .Y(_07258_));
 sky130_fd_sc_hd__nand4_2 _15130_ (.A(_07126_),
    .B(_07176_),
    .C(_07225_),
    .D(_07124_),
    .Y(_07259_));
 sky130_fd_sc_hd__a41o_1 _15131_ (.A1(_07126_),
    .A2(_07176_),
    .A3(_07225_),
    .A4(_07124_),
    .B1(_00834_),
    .X(_07260_));
 sky130_fd_sc_hd__xnor2_1 _15132_ (.A(_07258_),
    .B(_07260_),
    .Y(net117));
 sky130_fd_sc_hd__a21oi_1 _15133_ (.A1(_07242_),
    .A2(_07247_),
    .B1(_07241_),
    .Y(_07261_));
 sky130_fd_sc_hd__o21ba_1 _15134_ (.A1(_07191_),
    .A2(_07233_),
    .B1_N(_07234_),
    .X(_07262_));
 sky130_fd_sc_hd__o41a_1 _15135_ (.A1(_02925_),
    .A2(_03086_),
    .A3(_03449_),
    .A4(_03583_),
    .B1(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__and4b_1 _15136_ (.A_N(_07262_),
    .B(_03584_),
    .C(_02924_),
    .D(_02922_),
    .X(_07265_));
 sky130_fd_sc_hd__a31o_1 _15137_ (.A1(_07265_),
    .A2(_03450_),
    .A3(_03087_),
    .B1(_07263_),
    .X(_07266_));
 sky130_fd_sc_hd__a32o_1 _15138_ (.A1(_03180_),
    .A2(_03653_),
    .A3(_07193_),
    .B1(_03831_),
    .B2(_02858_),
    .X(_07267_));
 sky130_fd_sc_hd__o21bai_1 _15139_ (.A1(_07245_),
    .A2(_07262_),
    .B1_N(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__a2bb2o_1 _15140_ (.A1_N(_07263_),
    .A2_N(_07268_),
    .B1(_07267_),
    .B2(_07266_),
    .X(_07269_));
 sky130_fd_sc_hd__and3_1 _15141_ (.A(_07228_),
    .B(_07239_),
    .C(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__a21oi_1 _15142_ (.A1(_07228_),
    .A2(_07239_),
    .B1(_07269_),
    .Y(_07271_));
 sky130_fd_sc_hd__a32o_1 _15143_ (.A1(_03320_),
    .A2(_03445_),
    .A3(_03448_),
    .B1(_03584_),
    .B2(_03087_),
    .X(_07272_));
 sky130_fd_sc_hd__or4_2 _15144_ (.A(_03086_),
    .B(_03319_),
    .C(_03449_),
    .D(_03583_),
    .X(_07273_));
 sky130_fd_sc_hd__a22o_1 _15145_ (.A1(net129),
    .A2(_02926_),
    .B1(_07273_),
    .B2(_07272_),
    .X(_07274_));
 sky130_fd_sc_hd__o21bai_1 _15146_ (.A1(_07270_),
    .A2(_07271_),
    .B1_N(_07274_),
    .Y(_07276_));
 sky130_fd_sc_hd__or3b_1 _15147_ (.A(_07270_),
    .B(_07271_),
    .C_N(_07274_),
    .X(_07277_));
 sky130_fd_sc_hd__a21oi_1 _15148_ (.A1(_07276_),
    .A2(_07277_),
    .B1(_07261_),
    .Y(_07278_));
 sky130_fd_sc_hd__nand3_1 _15149_ (.A(_07261_),
    .B(_07276_),
    .C(_07277_),
    .Y(_07279_));
 sky130_fd_sc_hd__and2b_1 _15150_ (.A_N(_07278_),
    .B(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__o21ba_1 _15151_ (.A1(_07208_),
    .A2(_07248_),
    .B1_N(_07250_),
    .X(_07281_));
 sky130_fd_sc_hd__a21oi_4 _15152_ (.A1(_07208_),
    .A2(_07248_),
    .B1(_07281_),
    .Y(_07282_));
 sky130_fd_sc_hd__inv_2 _15153_ (.A(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__xor2_4 _15154_ (.A(_07280_),
    .B(_07282_),
    .X(_07284_));
 sky130_fd_sc_hd__inv_2 _15155_ (.A(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__xnor2_1 _15156_ (.A(_07253_),
    .B(_07285_),
    .Y(_07287_));
 sky130_fd_sc_hd__a41oi_2 _15157_ (.A1(_07122_),
    .A2(_07172_),
    .A3(_07220_),
    .A4(_07255_),
    .B1(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__a31oi_2 _15158_ (.A1(_07223_),
    .A2(_07255_),
    .A3(_07284_),
    .B1(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__o22ai_4 _15159_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_07258_),
    .B2(_07259_),
    .Y(_07290_));
 sky130_fd_sc_hd__xnor2_1 _15160_ (.A(_07289_),
    .B(_07290_),
    .Y(net118));
 sky130_fd_sc_hd__o21ai_2 _15161_ (.A1(_07278_),
    .A2(_07283_),
    .B1(_07279_),
    .Y(_07291_));
 sky130_fd_sc_hd__a21bo_1 _15162_ (.A1(_07245_),
    .A2(_07262_),
    .B1_N(_07268_),
    .X(_07292_));
 sky130_fd_sc_hd__o31a_1 _15163_ (.A1(_03179_),
    .A2(_03652_),
    .A3(_07193_),
    .B1(_07273_),
    .X(_07293_));
 sky130_fd_sc_hd__nor4_1 _15164_ (.A(_03179_),
    .B(_03652_),
    .C(_07193_),
    .D(_07273_),
    .Y(_07294_));
 sky130_fd_sc_hd__nor2_1 _15165_ (.A(_07293_),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__o32a_1 _15166_ (.A1(_03319_),
    .A2(_03581_),
    .A3(_03582_),
    .B1(_03652_),
    .B2(_03449_),
    .X(_07297_));
 sky130_fd_sc_hd__or3_1 _15167_ (.A(_03581_),
    .B(_03582_),
    .C(_03652_),
    .X(_07298_));
 sky130_fd_sc_hd__and4_1 _15168_ (.A(_03320_),
    .B(_03450_),
    .C(_03584_),
    .D(_03653_),
    .X(_07299_));
 sky130_fd_sc_hd__a2bb2o_1 _15169_ (.A1_N(_07297_),
    .A2_N(_07299_),
    .B1(_03180_),
    .B2(_03831_),
    .X(_07300_));
 sky130_fd_sc_hd__or2_1 _15170_ (.A(_07300_),
    .B(_07295_),
    .X(_07301_));
 sky130_fd_sc_hd__nand2_1 _15171_ (.A(_07295_),
    .B(_07300_),
    .Y(_07302_));
 sky130_fd_sc_hd__and2_1 _15172_ (.A(_07301_),
    .B(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__and4b_1 _15173_ (.A_N(_07263_),
    .B(_07268_),
    .C(_07301_),
    .D(_07302_),
    .X(_07304_));
 sky130_fd_sc_hd__xnor2_1 _15174_ (.A(_07292_),
    .B(_07303_),
    .Y(_07305_));
 sky130_fd_sc_hd__and3_1 _15175_ (.A(net129),
    .B(_03084_),
    .C(_03082_),
    .X(_07306_));
 sky130_fd_sc_hd__o21bai_1 _15176_ (.A1(_07274_),
    .A2(_07270_),
    .B1_N(_07271_),
    .Y(_07308_));
 sky130_fd_sc_hd__o21ba_1 _15177_ (.A1(_07305_),
    .A2(_07306_),
    .B1_N(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__or3b_1 _15178_ (.A(_07305_),
    .B(_07306_),
    .C_N(_07308_),
    .X(_07310_));
 sky130_fd_sc_hd__and2b_1 _15179_ (.A_N(_07309_),
    .B(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__xor2_2 _15180_ (.A(_07291_),
    .B(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__xnor2_1 _15181_ (.A(_07291_),
    .B(_07311_),
    .Y(_07313_));
 sky130_fd_sc_hd__or4_1 _15182_ (.A(_07251_),
    .B(_07285_),
    .C(_07313_),
    .D(_07219_),
    .X(_07314_));
 sky130_fd_sc_hd__a31o_1 _15183_ (.A1(_07218_),
    .A2(_07252_),
    .A3(_07284_),
    .B1(_07312_),
    .X(_07315_));
 sky130_fd_sc_hd__o2bb2ai_1 _15184_ (.A1_N(_07314_),
    .A2_N(_07315_),
    .B1(_07257_),
    .B2(_07285_),
    .Y(_07316_));
 sky130_fd_sc_hd__nor3_1 _15185_ (.A(_07257_),
    .B(_07285_),
    .C(_07313_),
    .Y(_07317_));
 sky130_fd_sc_hd__nand4_4 _15186_ (.A(_07223_),
    .B(_07255_),
    .C(_07284_),
    .D(_07312_),
    .Y(_07319_));
 sky130_fd_sc_hd__nand2_2 _15187_ (.A(_07316_),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__a311o_1 _15188_ (.A1(_07223_),
    .A2(_07255_),
    .A3(_07284_),
    .B1(_07288_),
    .C1(_00834_),
    .X(_07321_));
 sky130_fd_sc_hd__o31ai_2 _15189_ (.A1(_07258_),
    .A2(_07289_),
    .A3(_07259_),
    .B1(_00845_),
    .Y(_07322_));
 sky130_fd_sc_hd__xor2_1 _15190_ (.A(_07320_),
    .B(_07322_),
    .X(net119));
 sky130_fd_sc_hd__o221a_1 _15191_ (.A1(_03449_),
    .A2(_03832_),
    .B1(_03912_),
    .B2(_03319_),
    .C1(_07298_),
    .X(_07323_));
 sky130_fd_sc_hd__o41a_1 _15192_ (.A1(_03179_),
    .A2(_03652_),
    .A3(_07193_),
    .A4(_07273_),
    .B1(_07302_),
    .X(_07324_));
 sky130_fd_sc_hd__nor2_1 _15193_ (.A(_07323_),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__nand2_1 _15194_ (.A(_07324_),
    .B(_07323_),
    .Y(_07326_));
 sky130_fd_sc_hd__or3b_1 _15195_ (.A(_07299_),
    .B(_07325_),
    .C_N(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__o41a_1 _15196_ (.A1(_03179_),
    .A2(_03652_),
    .A3(_07193_),
    .A4(_07273_),
    .B1(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__nor3b_1 _15197_ (.A(_07294_),
    .B(_07304_),
    .C_N(_07327_),
    .Y(_07329_));
 sky130_fd_sc_hd__a21oi_1 _15198_ (.A1(_07291_),
    .A2(_07310_),
    .B1(_07309_),
    .Y(_07330_));
 sky130_fd_sc_hd__and4bb_1 _15199_ (.A_N(_07294_),
    .B_N(_07304_),
    .C(_07327_),
    .D(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__or3b_1 _15200_ (.A(_07292_),
    .B(_07328_),
    .C_N(_07303_),
    .X(_07332_));
 sky130_fd_sc_hd__o21ai_1 _15201_ (.A1(_07329_),
    .A2(_07330_),
    .B1(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__or2_2 _15202_ (.A(_07331_),
    .B(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__inv_2 _15203_ (.A(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__o41a_1 _15204_ (.A1(_07251_),
    .A2(_07285_),
    .A3(_07313_),
    .A4(_07219_),
    .B1(_07334_),
    .X(_07336_));
 sky130_fd_sc_hd__and4_1 _15205_ (.A(_07253_),
    .B(_07284_),
    .C(_07312_),
    .D(_07335_),
    .X(_07337_));
 sky130_fd_sc_hd__o21ai_2 _15206_ (.A1(_07336_),
    .A2(_07337_),
    .B1(_07319_),
    .Y(_07339_));
 sky130_fd_sc_hd__or4_1 _15207_ (.A(_07257_),
    .B(_07285_),
    .C(_07313_),
    .D(_07334_),
    .X(_07340_));
 sky130_fd_sc_hd__o211ai_1 _15208_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_07316_),
    .C1(_07319_),
    .Y(_07341_));
 sky130_fd_sc_hd__o2111ai_1 _15209_ (.A1(_00834_),
    .A2(_07320_),
    .B1(_07339_),
    .C1(_07340_),
    .D1(_07322_),
    .Y(_07342_));
 sky130_fd_sc_hd__a32o_1 _15210_ (.A1(_07290_),
    .A2(_07321_),
    .A3(_07341_),
    .B1(_07340_),
    .B2(_07339_),
    .X(_07343_));
 sky130_fd_sc_hd__nand2_1 _15211_ (.A(_07342_),
    .B(_07343_),
    .Y(net121));
 sky130_fd_sc_hd__or4_1 _15212_ (.A(_03645_),
    .B(_03830_),
    .C(_03581_),
    .D(_03582_),
    .X(_07344_));
 sky130_fd_sc_hd__o221a_1 _15213_ (.A1(_03652_),
    .A2(_03912_),
    .B1(_07323_),
    .B2(_07324_),
    .C1(_07344_),
    .X(_07345_));
 sky130_fd_sc_hd__or4b_2 _15214_ (.A(_07299_),
    .B(_07333_),
    .C(_07337_),
    .D_N(_07345_),
    .X(_07346_));
 sky130_fd_sc_hd__o21bai_1 _15215_ (.A1(_07319_),
    .A2(_07334_),
    .B1_N(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__nand3_1 _15216_ (.A(_07317_),
    .B(_07335_),
    .C(_07346_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand2_1 _15217_ (.A(_07347_),
    .B(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__o221ai_4 _15218_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_07319_),
    .B2(_07334_),
    .C1(_07339_),
    .Y(_07351_));
 sky130_fd_sc_hd__o2111a_1 _15219_ (.A1(_00834_),
    .A2(_07320_),
    .B1(_07321_),
    .C1(_07351_),
    .D1(_07290_),
    .X(_07352_));
 sky130_fd_sc_hd__o2111ai_2 _15220_ (.A1(_00834_),
    .A2(_07320_),
    .B1(_07321_),
    .C1(_07351_),
    .D1(_07290_),
    .Y(_07353_));
 sky130_fd_sc_hd__xnor2_1 _15221_ (.A(_07350_),
    .B(_07353_),
    .Y(net122));
 sky130_fd_sc_hd__nor2_1 _15222_ (.A(_03832_),
    .B(_03912_),
    .Y(_07354_));
 sky130_fd_sc_hd__nand4_2 _15223_ (.A(_07317_),
    .B(_07335_),
    .C(_07346_),
    .D(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__a31o_1 _15224_ (.A1(_07317_),
    .A2(_07335_),
    .A3(_07346_),
    .B1(_07354_),
    .X(_07356_));
 sky130_fd_sc_hd__and3_1 _15225_ (.A(_00845_),
    .B(_07347_),
    .C(_07349_),
    .X(_07357_));
 sky130_fd_sc_hd__o211ai_1 _15226_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_07347_),
    .C1(_07349_),
    .Y(_07359_));
 sky130_fd_sc_hd__o2111a_1 _15227_ (.A1(_00834_),
    .A2(_07320_),
    .B1(_07351_),
    .C1(_07359_),
    .D1(_07322_),
    .X(_07360_));
 sky130_fd_sc_hd__o2111ai_1 _15228_ (.A1(_00834_),
    .A2(_07350_),
    .B1(_07355_),
    .C1(_07356_),
    .D1(_07352_),
    .Y(_07361_));
 sky130_fd_sc_hd__o2bb2ai_1 _15229_ (.A1_N(_07355_),
    .A2_N(_07356_),
    .B1(_07353_),
    .B2(_07357_),
    .Y(_07362_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_07361_),
    .B(_07362_),
    .Y(net123));
 sky130_fd_sc_hd__o211ai_1 _15231_ (.A1(_00812_),
    .A2(_00823_),
    .B1(_07355_),
    .C1(_07356_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand4_1 _15232_ (.A(_07352_),
    .B(_07355_),
    .C(_07359_),
    .D(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__o21a_1 _15233_ (.A1(_07355_),
    .A2(_07360_),
    .B1(_07364_),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_16 input1 (.A(signed_A[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_8 input2 (.A(signed_A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_8 input3 (.A(signed_A[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(signed_A[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(signed_A[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(signed_A[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input7 (.A(signed_A[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(signed_A[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_8 input9 (.A(signed_A[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(signed_A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(signed_A[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(signed_A[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_8 input13 (.A(signed_A[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(signed_A[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(signed_A[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(signed_A[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(signed_A[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(signed_A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_8 input19 (.A(signed_A[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(signed_A[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(signed_A[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(signed_A[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(signed_A[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(signed_A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_12 input25 (.A(signed_A[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(signed_A[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(signed_A[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(signed_A[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(signed_A[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(signed_A[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(signed_A[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(signed_A[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_16 input33 (.A(signed_B[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(signed_B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_8 input35 (.A(signed_B[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(signed_B[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_8 input37 (.A(signed_B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_8 input38 (.A(signed_B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(signed_B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 input40 (.A(signed_B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_4 input41 (.A(signed_B[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 input42 (.A(signed_B[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_8 input43 (.A(signed_B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(signed_B[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_6 input45 (.A(signed_B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_8 input46 (.A(signed_B[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_8 input47 (.A(signed_B[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(signed_B[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(signed_B[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input50 (.A(signed_B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 input51 (.A(signed_B[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(signed_B[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(signed_B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_4 input54 (.A(signed_B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(signed_B[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_4 input56 (.A(signed_B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_12 input57 (.A(signed_B[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 input58 (.A(signed_B[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 input59 (.A(signed_B[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_6 input60 (.A(signed_B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_8 input61 (.A(signed_B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_8 input62 (.A(signed_B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_4 input63 (.A(signed_B[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(signed_B[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(product[0]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(product[10]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(product[11]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(product[12]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(product[13]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(product[14]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(product[15]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(product[16]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(product[17]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(product[18]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(product[19]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(product[1]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(product[20]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(product[21]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(product[22]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(product[23]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(product[24]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(product[25]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(product[26]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(product[27]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(product[28]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(product[29]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(product[2]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(product[30]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(product[31]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(product[32]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(product[33]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(product[34]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(product[35]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(product[36]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(product[37]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(product[38]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(product[39]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(product[3]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(product[40]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(product[41]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(product[42]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(product[43]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(product[44]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(product[45]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(product[46]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(product[47]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(product[48]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(product[49]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(product[4]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(product[50]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(product[51]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(product[52]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(product[53]));
 sky130_fd_sc_hd__buf_1 output114 (.A(net114),
    .X(product[54]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(product[55]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(product[56]));
 sky130_fd_sc_hd__buf_1 output117 (.A(net117),
    .X(product[57]));
 sky130_fd_sc_hd__buf_1 output118 (.A(net118),
    .X(product[58]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(product[59]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(product[5]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(product[60]));
 sky130_fd_sc_hd__buf_1 output122 (.A(net122),
    .X(product[61]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(product[62]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(product[63]));
 sky130_fd_sc_hd__buf_1 output125 (.A(net125),
    .X(product[6]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(product[7]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(product[8]));
 sky130_fd_sc_hd__buf_1 output128 (.A(net128),
    .X(product[9]));
 sky130_fd_sc_hd__buf_4 max_cap129 (.A(_03911_),
    .X(net129));
 sky130_fd_sc_hd__buf_8 max_cap130 (.A(_03083_),
    .X(net130));
 sky130_fd_sc_hd__buf_4 wire131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_4 max_cap132 (.A(_03081_),
    .X(net132));
 sky130_fd_sc_hd__buf_6 max_cap133 (.A(_02092_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 max_cap134 (.A(_01880_),
    .X(net134));
 sky130_fd_sc_hd__buf_6 max_cap135 (.A(_01879_),
    .X(net135));
 sky130_fd_sc_hd__buf_12 max_cap136 (.A(_01406_),
    .X(net136));
 sky130_fd_sc_hd__buf_8 wire137 (.A(_01405_),
    .X(net137));
 sky130_fd_sc_hd__buf_4 wire138 (.A(_02426_),
    .X(net138));
 sky130_fd_sc_hd__buf_8 max_cap139 (.A(_02236_),
    .X(net139));
 sky130_fd_sc_hd__buf_8 max_cap140 (.A(_01661_),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_16 max_cap141 (.A(_01059_),
    .X(net141));
 sky130_fd_sc_hd__buf_8 max_cap142 (.A(_00428_),
    .X(net142));
 sky130_fd_sc_hd__buf_12 max_cap143 (.A(_00149_),
    .X(net143));
 sky130_fd_sc_hd__buf_12 max_cap144 (.A(_00149_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_8 max_cap145 (.A(_01218_),
    .X(net145));
 sky130_fd_sc_hd__buf_8 max_cap146 (.A(_00566_),
    .X(net146));
 sky130_fd_sc_hd__buf_8 max_cap147 (.A(_00565_),
    .X(net147));
 sky130_fd_sc_hd__buf_8 max_cap148 (.A(_00071_),
    .X(net148));
 sky130_fd_sc_hd__buf_6 max_cap149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__buf_6 max_cap150 (.A(_07539_),
    .X(net150));
 sky130_fd_sc_hd__buf_12 max_cap151 (.A(_07370_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_8 max_cap152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_8 max_cap153 (.A(_07369_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_8 max_cap154 (.A(_07437_),
    .X(net154));
 sky130_fd_sc_hd__buf_6 max_cap155 (.A(_04715_),
    .X(net155));
 sky130_fd_sc_hd__buf_8 max_cap156 (.A(_03555_),
    .X(net156));
 sky130_fd_sc_hd__buf_6 max_cap157 (.A(_03555_),
    .X(net157));
 sky130_fd_sc_hd__buf_8 max_cap158 (.A(_03544_),
    .X(net158));
 sky130_fd_sc_hd__buf_12 max_cap159 (.A(_02855_),
    .X(net159));
 sky130_fd_sc_hd__buf_4 max_cap160 (.A(_00063_),
    .X(net160));
 sky130_fd_sc_hd__buf_4 max_cap161 (.A(_07504_),
    .X(net161));
 sky130_fd_sc_hd__buf_6 max_cap162 (.A(_07436_),
    .X(net162));
 sky130_fd_sc_hd__buf_8 max_cap163 (.A(_02800_),
    .X(net163));
 sky130_fd_sc_hd__buf_12 max_cap164 (.A(_01194_),
    .X(net164));
 sky130_fd_sc_hd__buf_8 max_cap165 (.A(_01183_),
    .X(net165));
 sky130_fd_sc_hd__buf_6 max_cap166 (.A(_01183_),
    .X(net166));
 sky130_fd_sc_hd__buf_4 max_cap167 (.A(_02811_),
    .X(net167));
 sky130_fd_sc_hd__buf_4 max_cap168 (.A(_02790_),
    .X(net168));
 sky130_fd_sc_hd__buf_6 max_cap169 (.A(_02790_),
    .X(net169));
 sky130_fd_sc_hd__buf_4 max_cap170 (.A(_02035_),
    .X(net170));
 sky130_fd_sc_hd__buf_4 max_cap171 (.A(_01870_),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 max_cap172 (.A(_00921_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_16 max_cap173 (.A(net57),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_16 max_cap174 (.A(net25),
    .X(net174));
endmodule
